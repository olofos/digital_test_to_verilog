//  A testbench for adder_tb
`timescale 1us/1ns

module adder_tb;
    reg [7:0] A;
    reg [7:0] B;
    wire [7:0] S;
    wire C;

  adder adder0 (
    .A(A),
    .B(B),
    .S(S),
    .C(C)
  );

    reg [24:0] patterns[0:65537];
    integer i;

    initial begin
      patterns[0] = 25'b00000001_00000001_00000010_0;
      patterns[1] = 25'b11111111_00000001_00000000_1;
      patterns[2] = 25'b00000000_00000000_00000000_0;
      patterns[3] = 25'b00000000_00000001_00000001_0;
      patterns[4] = 25'b00000000_00000010_00000010_0;
      patterns[5] = 25'b00000000_00000011_00000011_0;
      patterns[6] = 25'b00000000_00000100_00000100_0;
      patterns[7] = 25'b00000000_00000101_00000101_0;
      patterns[8] = 25'b00000000_00000110_00000110_0;
      patterns[9] = 25'b00000000_00000111_00000111_0;
      patterns[10] = 25'b00000000_00001000_00001000_0;
      patterns[11] = 25'b00000000_00001001_00001001_0;
      patterns[12] = 25'b00000000_00001010_00001010_0;
      patterns[13] = 25'b00000000_00001011_00001011_0;
      patterns[14] = 25'b00000000_00001100_00001100_0;
      patterns[15] = 25'b00000000_00001101_00001101_0;
      patterns[16] = 25'b00000000_00001110_00001110_0;
      patterns[17] = 25'b00000000_00001111_00001111_0;
      patterns[18] = 25'b00000000_00010000_00010000_0;
      patterns[19] = 25'b00000000_00010001_00010001_0;
      patterns[20] = 25'b00000000_00010010_00010010_0;
      patterns[21] = 25'b00000000_00010011_00010011_0;
      patterns[22] = 25'b00000000_00010100_00010100_0;
      patterns[23] = 25'b00000000_00010101_00010101_0;
      patterns[24] = 25'b00000000_00010110_00010110_0;
      patterns[25] = 25'b00000000_00010111_00010111_0;
      patterns[26] = 25'b00000000_00011000_00011000_0;
      patterns[27] = 25'b00000000_00011001_00011001_0;
      patterns[28] = 25'b00000000_00011010_00011010_0;
      patterns[29] = 25'b00000000_00011011_00011011_0;
      patterns[30] = 25'b00000000_00011100_00011100_0;
      patterns[31] = 25'b00000000_00011101_00011101_0;
      patterns[32] = 25'b00000000_00011110_00011110_0;
      patterns[33] = 25'b00000000_00011111_00011111_0;
      patterns[34] = 25'b00000000_00100000_00100000_0;
      patterns[35] = 25'b00000000_00100001_00100001_0;
      patterns[36] = 25'b00000000_00100010_00100010_0;
      patterns[37] = 25'b00000000_00100011_00100011_0;
      patterns[38] = 25'b00000000_00100100_00100100_0;
      patterns[39] = 25'b00000000_00100101_00100101_0;
      patterns[40] = 25'b00000000_00100110_00100110_0;
      patterns[41] = 25'b00000000_00100111_00100111_0;
      patterns[42] = 25'b00000000_00101000_00101000_0;
      patterns[43] = 25'b00000000_00101001_00101001_0;
      patterns[44] = 25'b00000000_00101010_00101010_0;
      patterns[45] = 25'b00000000_00101011_00101011_0;
      patterns[46] = 25'b00000000_00101100_00101100_0;
      patterns[47] = 25'b00000000_00101101_00101101_0;
      patterns[48] = 25'b00000000_00101110_00101110_0;
      patterns[49] = 25'b00000000_00101111_00101111_0;
      patterns[50] = 25'b00000000_00110000_00110000_0;
      patterns[51] = 25'b00000000_00110001_00110001_0;
      patterns[52] = 25'b00000000_00110010_00110010_0;
      patterns[53] = 25'b00000000_00110011_00110011_0;
      patterns[54] = 25'b00000000_00110100_00110100_0;
      patterns[55] = 25'b00000000_00110101_00110101_0;
      patterns[56] = 25'b00000000_00110110_00110110_0;
      patterns[57] = 25'b00000000_00110111_00110111_0;
      patterns[58] = 25'b00000000_00111000_00111000_0;
      patterns[59] = 25'b00000000_00111001_00111001_0;
      patterns[60] = 25'b00000000_00111010_00111010_0;
      patterns[61] = 25'b00000000_00111011_00111011_0;
      patterns[62] = 25'b00000000_00111100_00111100_0;
      patterns[63] = 25'b00000000_00111101_00111101_0;
      patterns[64] = 25'b00000000_00111110_00111110_0;
      patterns[65] = 25'b00000000_00111111_00111111_0;
      patterns[66] = 25'b00000000_01000000_01000000_0;
      patterns[67] = 25'b00000000_01000001_01000001_0;
      patterns[68] = 25'b00000000_01000010_01000010_0;
      patterns[69] = 25'b00000000_01000011_01000011_0;
      patterns[70] = 25'b00000000_01000100_01000100_0;
      patterns[71] = 25'b00000000_01000101_01000101_0;
      patterns[72] = 25'b00000000_01000110_01000110_0;
      patterns[73] = 25'b00000000_01000111_01000111_0;
      patterns[74] = 25'b00000000_01001000_01001000_0;
      patterns[75] = 25'b00000000_01001001_01001001_0;
      patterns[76] = 25'b00000000_01001010_01001010_0;
      patterns[77] = 25'b00000000_01001011_01001011_0;
      patterns[78] = 25'b00000000_01001100_01001100_0;
      patterns[79] = 25'b00000000_01001101_01001101_0;
      patterns[80] = 25'b00000000_01001110_01001110_0;
      patterns[81] = 25'b00000000_01001111_01001111_0;
      patterns[82] = 25'b00000000_01010000_01010000_0;
      patterns[83] = 25'b00000000_01010001_01010001_0;
      patterns[84] = 25'b00000000_01010010_01010010_0;
      patterns[85] = 25'b00000000_01010011_01010011_0;
      patterns[86] = 25'b00000000_01010100_01010100_0;
      patterns[87] = 25'b00000000_01010101_01010101_0;
      patterns[88] = 25'b00000000_01010110_01010110_0;
      patterns[89] = 25'b00000000_01010111_01010111_0;
      patterns[90] = 25'b00000000_01011000_01011000_0;
      patterns[91] = 25'b00000000_01011001_01011001_0;
      patterns[92] = 25'b00000000_01011010_01011010_0;
      patterns[93] = 25'b00000000_01011011_01011011_0;
      patterns[94] = 25'b00000000_01011100_01011100_0;
      patterns[95] = 25'b00000000_01011101_01011101_0;
      patterns[96] = 25'b00000000_01011110_01011110_0;
      patterns[97] = 25'b00000000_01011111_01011111_0;
      patterns[98] = 25'b00000000_01100000_01100000_0;
      patterns[99] = 25'b00000000_01100001_01100001_0;
      patterns[100] = 25'b00000000_01100010_01100010_0;
      patterns[101] = 25'b00000000_01100011_01100011_0;
      patterns[102] = 25'b00000000_01100100_01100100_0;
      patterns[103] = 25'b00000000_01100101_01100101_0;
      patterns[104] = 25'b00000000_01100110_01100110_0;
      patterns[105] = 25'b00000000_01100111_01100111_0;
      patterns[106] = 25'b00000000_01101000_01101000_0;
      patterns[107] = 25'b00000000_01101001_01101001_0;
      patterns[108] = 25'b00000000_01101010_01101010_0;
      patterns[109] = 25'b00000000_01101011_01101011_0;
      patterns[110] = 25'b00000000_01101100_01101100_0;
      patterns[111] = 25'b00000000_01101101_01101101_0;
      patterns[112] = 25'b00000000_01101110_01101110_0;
      patterns[113] = 25'b00000000_01101111_01101111_0;
      patterns[114] = 25'b00000000_01110000_01110000_0;
      patterns[115] = 25'b00000000_01110001_01110001_0;
      patterns[116] = 25'b00000000_01110010_01110010_0;
      patterns[117] = 25'b00000000_01110011_01110011_0;
      patterns[118] = 25'b00000000_01110100_01110100_0;
      patterns[119] = 25'b00000000_01110101_01110101_0;
      patterns[120] = 25'b00000000_01110110_01110110_0;
      patterns[121] = 25'b00000000_01110111_01110111_0;
      patterns[122] = 25'b00000000_01111000_01111000_0;
      patterns[123] = 25'b00000000_01111001_01111001_0;
      patterns[124] = 25'b00000000_01111010_01111010_0;
      patterns[125] = 25'b00000000_01111011_01111011_0;
      patterns[126] = 25'b00000000_01111100_01111100_0;
      patterns[127] = 25'b00000000_01111101_01111101_0;
      patterns[128] = 25'b00000000_01111110_01111110_0;
      patterns[129] = 25'b00000000_01111111_01111111_0;
      patterns[130] = 25'b00000000_10000000_10000000_0;
      patterns[131] = 25'b00000000_10000001_10000001_0;
      patterns[132] = 25'b00000000_10000010_10000010_0;
      patterns[133] = 25'b00000000_10000011_10000011_0;
      patterns[134] = 25'b00000000_10000100_10000100_0;
      patterns[135] = 25'b00000000_10000101_10000101_0;
      patterns[136] = 25'b00000000_10000110_10000110_0;
      patterns[137] = 25'b00000000_10000111_10000111_0;
      patterns[138] = 25'b00000000_10001000_10001000_0;
      patterns[139] = 25'b00000000_10001001_10001001_0;
      patterns[140] = 25'b00000000_10001010_10001010_0;
      patterns[141] = 25'b00000000_10001011_10001011_0;
      patterns[142] = 25'b00000000_10001100_10001100_0;
      patterns[143] = 25'b00000000_10001101_10001101_0;
      patterns[144] = 25'b00000000_10001110_10001110_0;
      patterns[145] = 25'b00000000_10001111_10001111_0;
      patterns[146] = 25'b00000000_10010000_10010000_0;
      patterns[147] = 25'b00000000_10010001_10010001_0;
      patterns[148] = 25'b00000000_10010010_10010010_0;
      patterns[149] = 25'b00000000_10010011_10010011_0;
      patterns[150] = 25'b00000000_10010100_10010100_0;
      patterns[151] = 25'b00000000_10010101_10010101_0;
      patterns[152] = 25'b00000000_10010110_10010110_0;
      patterns[153] = 25'b00000000_10010111_10010111_0;
      patterns[154] = 25'b00000000_10011000_10011000_0;
      patterns[155] = 25'b00000000_10011001_10011001_0;
      patterns[156] = 25'b00000000_10011010_10011010_0;
      patterns[157] = 25'b00000000_10011011_10011011_0;
      patterns[158] = 25'b00000000_10011100_10011100_0;
      patterns[159] = 25'b00000000_10011101_10011101_0;
      patterns[160] = 25'b00000000_10011110_10011110_0;
      patterns[161] = 25'b00000000_10011111_10011111_0;
      patterns[162] = 25'b00000000_10100000_10100000_0;
      patterns[163] = 25'b00000000_10100001_10100001_0;
      patterns[164] = 25'b00000000_10100010_10100010_0;
      patterns[165] = 25'b00000000_10100011_10100011_0;
      patterns[166] = 25'b00000000_10100100_10100100_0;
      patterns[167] = 25'b00000000_10100101_10100101_0;
      patterns[168] = 25'b00000000_10100110_10100110_0;
      patterns[169] = 25'b00000000_10100111_10100111_0;
      patterns[170] = 25'b00000000_10101000_10101000_0;
      patterns[171] = 25'b00000000_10101001_10101001_0;
      patterns[172] = 25'b00000000_10101010_10101010_0;
      patterns[173] = 25'b00000000_10101011_10101011_0;
      patterns[174] = 25'b00000000_10101100_10101100_0;
      patterns[175] = 25'b00000000_10101101_10101101_0;
      patterns[176] = 25'b00000000_10101110_10101110_0;
      patterns[177] = 25'b00000000_10101111_10101111_0;
      patterns[178] = 25'b00000000_10110000_10110000_0;
      patterns[179] = 25'b00000000_10110001_10110001_0;
      patterns[180] = 25'b00000000_10110010_10110010_0;
      patterns[181] = 25'b00000000_10110011_10110011_0;
      patterns[182] = 25'b00000000_10110100_10110100_0;
      patterns[183] = 25'b00000000_10110101_10110101_0;
      patterns[184] = 25'b00000000_10110110_10110110_0;
      patterns[185] = 25'b00000000_10110111_10110111_0;
      patterns[186] = 25'b00000000_10111000_10111000_0;
      patterns[187] = 25'b00000000_10111001_10111001_0;
      patterns[188] = 25'b00000000_10111010_10111010_0;
      patterns[189] = 25'b00000000_10111011_10111011_0;
      patterns[190] = 25'b00000000_10111100_10111100_0;
      patterns[191] = 25'b00000000_10111101_10111101_0;
      patterns[192] = 25'b00000000_10111110_10111110_0;
      patterns[193] = 25'b00000000_10111111_10111111_0;
      patterns[194] = 25'b00000000_11000000_11000000_0;
      patterns[195] = 25'b00000000_11000001_11000001_0;
      patterns[196] = 25'b00000000_11000010_11000010_0;
      patterns[197] = 25'b00000000_11000011_11000011_0;
      patterns[198] = 25'b00000000_11000100_11000100_0;
      patterns[199] = 25'b00000000_11000101_11000101_0;
      patterns[200] = 25'b00000000_11000110_11000110_0;
      patterns[201] = 25'b00000000_11000111_11000111_0;
      patterns[202] = 25'b00000000_11001000_11001000_0;
      patterns[203] = 25'b00000000_11001001_11001001_0;
      patterns[204] = 25'b00000000_11001010_11001010_0;
      patterns[205] = 25'b00000000_11001011_11001011_0;
      patterns[206] = 25'b00000000_11001100_11001100_0;
      patterns[207] = 25'b00000000_11001101_11001101_0;
      patterns[208] = 25'b00000000_11001110_11001110_0;
      patterns[209] = 25'b00000000_11001111_11001111_0;
      patterns[210] = 25'b00000000_11010000_11010000_0;
      patterns[211] = 25'b00000000_11010001_11010001_0;
      patterns[212] = 25'b00000000_11010010_11010010_0;
      patterns[213] = 25'b00000000_11010011_11010011_0;
      patterns[214] = 25'b00000000_11010100_11010100_0;
      patterns[215] = 25'b00000000_11010101_11010101_0;
      patterns[216] = 25'b00000000_11010110_11010110_0;
      patterns[217] = 25'b00000000_11010111_11010111_0;
      patterns[218] = 25'b00000000_11011000_11011000_0;
      patterns[219] = 25'b00000000_11011001_11011001_0;
      patterns[220] = 25'b00000000_11011010_11011010_0;
      patterns[221] = 25'b00000000_11011011_11011011_0;
      patterns[222] = 25'b00000000_11011100_11011100_0;
      patterns[223] = 25'b00000000_11011101_11011101_0;
      patterns[224] = 25'b00000000_11011110_11011110_0;
      patterns[225] = 25'b00000000_11011111_11011111_0;
      patterns[226] = 25'b00000000_11100000_11100000_0;
      patterns[227] = 25'b00000000_11100001_11100001_0;
      patterns[228] = 25'b00000000_11100010_11100010_0;
      patterns[229] = 25'b00000000_11100011_11100011_0;
      patterns[230] = 25'b00000000_11100100_11100100_0;
      patterns[231] = 25'b00000000_11100101_11100101_0;
      patterns[232] = 25'b00000000_11100110_11100110_0;
      patterns[233] = 25'b00000000_11100111_11100111_0;
      patterns[234] = 25'b00000000_11101000_11101000_0;
      patterns[235] = 25'b00000000_11101001_11101001_0;
      patterns[236] = 25'b00000000_11101010_11101010_0;
      patterns[237] = 25'b00000000_11101011_11101011_0;
      patterns[238] = 25'b00000000_11101100_11101100_0;
      patterns[239] = 25'b00000000_11101101_11101101_0;
      patterns[240] = 25'b00000000_11101110_11101110_0;
      patterns[241] = 25'b00000000_11101111_11101111_0;
      patterns[242] = 25'b00000000_11110000_11110000_0;
      patterns[243] = 25'b00000000_11110001_11110001_0;
      patterns[244] = 25'b00000000_11110010_11110010_0;
      patterns[245] = 25'b00000000_11110011_11110011_0;
      patterns[246] = 25'b00000000_11110100_11110100_0;
      patterns[247] = 25'b00000000_11110101_11110101_0;
      patterns[248] = 25'b00000000_11110110_11110110_0;
      patterns[249] = 25'b00000000_11110111_11110111_0;
      patterns[250] = 25'b00000000_11111000_11111000_0;
      patterns[251] = 25'b00000000_11111001_11111001_0;
      patterns[252] = 25'b00000000_11111010_11111010_0;
      patterns[253] = 25'b00000000_11111011_11111011_0;
      patterns[254] = 25'b00000000_11111100_11111100_0;
      patterns[255] = 25'b00000000_11111101_11111101_0;
      patterns[256] = 25'b00000000_11111110_11111110_0;
      patterns[257] = 25'b00000000_11111111_11111111_0;
      patterns[258] = 25'b00000001_00000000_00000001_0;
      patterns[259] = 25'b00000001_00000001_00000010_0;
      patterns[260] = 25'b00000001_00000010_00000011_0;
      patterns[261] = 25'b00000001_00000011_00000100_0;
      patterns[262] = 25'b00000001_00000100_00000101_0;
      patterns[263] = 25'b00000001_00000101_00000110_0;
      patterns[264] = 25'b00000001_00000110_00000111_0;
      patterns[265] = 25'b00000001_00000111_00001000_0;
      patterns[266] = 25'b00000001_00001000_00001001_0;
      patterns[267] = 25'b00000001_00001001_00001010_0;
      patterns[268] = 25'b00000001_00001010_00001011_0;
      patterns[269] = 25'b00000001_00001011_00001100_0;
      patterns[270] = 25'b00000001_00001100_00001101_0;
      patterns[271] = 25'b00000001_00001101_00001110_0;
      patterns[272] = 25'b00000001_00001110_00001111_0;
      patterns[273] = 25'b00000001_00001111_00010000_0;
      patterns[274] = 25'b00000001_00010000_00010001_0;
      patterns[275] = 25'b00000001_00010001_00010010_0;
      patterns[276] = 25'b00000001_00010010_00010011_0;
      patterns[277] = 25'b00000001_00010011_00010100_0;
      patterns[278] = 25'b00000001_00010100_00010101_0;
      patterns[279] = 25'b00000001_00010101_00010110_0;
      patterns[280] = 25'b00000001_00010110_00010111_0;
      patterns[281] = 25'b00000001_00010111_00011000_0;
      patterns[282] = 25'b00000001_00011000_00011001_0;
      patterns[283] = 25'b00000001_00011001_00011010_0;
      patterns[284] = 25'b00000001_00011010_00011011_0;
      patterns[285] = 25'b00000001_00011011_00011100_0;
      patterns[286] = 25'b00000001_00011100_00011101_0;
      patterns[287] = 25'b00000001_00011101_00011110_0;
      patterns[288] = 25'b00000001_00011110_00011111_0;
      patterns[289] = 25'b00000001_00011111_00100000_0;
      patterns[290] = 25'b00000001_00100000_00100001_0;
      patterns[291] = 25'b00000001_00100001_00100010_0;
      patterns[292] = 25'b00000001_00100010_00100011_0;
      patterns[293] = 25'b00000001_00100011_00100100_0;
      patterns[294] = 25'b00000001_00100100_00100101_0;
      patterns[295] = 25'b00000001_00100101_00100110_0;
      patterns[296] = 25'b00000001_00100110_00100111_0;
      patterns[297] = 25'b00000001_00100111_00101000_0;
      patterns[298] = 25'b00000001_00101000_00101001_0;
      patterns[299] = 25'b00000001_00101001_00101010_0;
      patterns[300] = 25'b00000001_00101010_00101011_0;
      patterns[301] = 25'b00000001_00101011_00101100_0;
      patterns[302] = 25'b00000001_00101100_00101101_0;
      patterns[303] = 25'b00000001_00101101_00101110_0;
      patterns[304] = 25'b00000001_00101110_00101111_0;
      patterns[305] = 25'b00000001_00101111_00110000_0;
      patterns[306] = 25'b00000001_00110000_00110001_0;
      patterns[307] = 25'b00000001_00110001_00110010_0;
      patterns[308] = 25'b00000001_00110010_00110011_0;
      patterns[309] = 25'b00000001_00110011_00110100_0;
      patterns[310] = 25'b00000001_00110100_00110101_0;
      patterns[311] = 25'b00000001_00110101_00110110_0;
      patterns[312] = 25'b00000001_00110110_00110111_0;
      patterns[313] = 25'b00000001_00110111_00111000_0;
      patterns[314] = 25'b00000001_00111000_00111001_0;
      patterns[315] = 25'b00000001_00111001_00111010_0;
      patterns[316] = 25'b00000001_00111010_00111011_0;
      patterns[317] = 25'b00000001_00111011_00111100_0;
      patterns[318] = 25'b00000001_00111100_00111101_0;
      patterns[319] = 25'b00000001_00111101_00111110_0;
      patterns[320] = 25'b00000001_00111110_00111111_0;
      patterns[321] = 25'b00000001_00111111_01000000_0;
      patterns[322] = 25'b00000001_01000000_01000001_0;
      patterns[323] = 25'b00000001_01000001_01000010_0;
      patterns[324] = 25'b00000001_01000010_01000011_0;
      patterns[325] = 25'b00000001_01000011_01000100_0;
      patterns[326] = 25'b00000001_01000100_01000101_0;
      patterns[327] = 25'b00000001_01000101_01000110_0;
      patterns[328] = 25'b00000001_01000110_01000111_0;
      patterns[329] = 25'b00000001_01000111_01001000_0;
      patterns[330] = 25'b00000001_01001000_01001001_0;
      patterns[331] = 25'b00000001_01001001_01001010_0;
      patterns[332] = 25'b00000001_01001010_01001011_0;
      patterns[333] = 25'b00000001_01001011_01001100_0;
      patterns[334] = 25'b00000001_01001100_01001101_0;
      patterns[335] = 25'b00000001_01001101_01001110_0;
      patterns[336] = 25'b00000001_01001110_01001111_0;
      patterns[337] = 25'b00000001_01001111_01010000_0;
      patterns[338] = 25'b00000001_01010000_01010001_0;
      patterns[339] = 25'b00000001_01010001_01010010_0;
      patterns[340] = 25'b00000001_01010010_01010011_0;
      patterns[341] = 25'b00000001_01010011_01010100_0;
      patterns[342] = 25'b00000001_01010100_01010101_0;
      patterns[343] = 25'b00000001_01010101_01010110_0;
      patterns[344] = 25'b00000001_01010110_01010111_0;
      patterns[345] = 25'b00000001_01010111_01011000_0;
      patterns[346] = 25'b00000001_01011000_01011001_0;
      patterns[347] = 25'b00000001_01011001_01011010_0;
      patterns[348] = 25'b00000001_01011010_01011011_0;
      patterns[349] = 25'b00000001_01011011_01011100_0;
      patterns[350] = 25'b00000001_01011100_01011101_0;
      patterns[351] = 25'b00000001_01011101_01011110_0;
      patterns[352] = 25'b00000001_01011110_01011111_0;
      patterns[353] = 25'b00000001_01011111_01100000_0;
      patterns[354] = 25'b00000001_01100000_01100001_0;
      patterns[355] = 25'b00000001_01100001_01100010_0;
      patterns[356] = 25'b00000001_01100010_01100011_0;
      patterns[357] = 25'b00000001_01100011_01100100_0;
      patterns[358] = 25'b00000001_01100100_01100101_0;
      patterns[359] = 25'b00000001_01100101_01100110_0;
      patterns[360] = 25'b00000001_01100110_01100111_0;
      patterns[361] = 25'b00000001_01100111_01101000_0;
      patterns[362] = 25'b00000001_01101000_01101001_0;
      patterns[363] = 25'b00000001_01101001_01101010_0;
      patterns[364] = 25'b00000001_01101010_01101011_0;
      patterns[365] = 25'b00000001_01101011_01101100_0;
      patterns[366] = 25'b00000001_01101100_01101101_0;
      patterns[367] = 25'b00000001_01101101_01101110_0;
      patterns[368] = 25'b00000001_01101110_01101111_0;
      patterns[369] = 25'b00000001_01101111_01110000_0;
      patterns[370] = 25'b00000001_01110000_01110001_0;
      patterns[371] = 25'b00000001_01110001_01110010_0;
      patterns[372] = 25'b00000001_01110010_01110011_0;
      patterns[373] = 25'b00000001_01110011_01110100_0;
      patterns[374] = 25'b00000001_01110100_01110101_0;
      patterns[375] = 25'b00000001_01110101_01110110_0;
      patterns[376] = 25'b00000001_01110110_01110111_0;
      patterns[377] = 25'b00000001_01110111_01111000_0;
      patterns[378] = 25'b00000001_01111000_01111001_0;
      patterns[379] = 25'b00000001_01111001_01111010_0;
      patterns[380] = 25'b00000001_01111010_01111011_0;
      patterns[381] = 25'b00000001_01111011_01111100_0;
      patterns[382] = 25'b00000001_01111100_01111101_0;
      patterns[383] = 25'b00000001_01111101_01111110_0;
      patterns[384] = 25'b00000001_01111110_01111111_0;
      patterns[385] = 25'b00000001_01111111_10000000_0;
      patterns[386] = 25'b00000001_10000000_10000001_0;
      patterns[387] = 25'b00000001_10000001_10000010_0;
      patterns[388] = 25'b00000001_10000010_10000011_0;
      patterns[389] = 25'b00000001_10000011_10000100_0;
      patterns[390] = 25'b00000001_10000100_10000101_0;
      patterns[391] = 25'b00000001_10000101_10000110_0;
      patterns[392] = 25'b00000001_10000110_10000111_0;
      patterns[393] = 25'b00000001_10000111_10001000_0;
      patterns[394] = 25'b00000001_10001000_10001001_0;
      patterns[395] = 25'b00000001_10001001_10001010_0;
      patterns[396] = 25'b00000001_10001010_10001011_0;
      patterns[397] = 25'b00000001_10001011_10001100_0;
      patterns[398] = 25'b00000001_10001100_10001101_0;
      patterns[399] = 25'b00000001_10001101_10001110_0;
      patterns[400] = 25'b00000001_10001110_10001111_0;
      patterns[401] = 25'b00000001_10001111_10010000_0;
      patterns[402] = 25'b00000001_10010000_10010001_0;
      patterns[403] = 25'b00000001_10010001_10010010_0;
      patterns[404] = 25'b00000001_10010010_10010011_0;
      patterns[405] = 25'b00000001_10010011_10010100_0;
      patterns[406] = 25'b00000001_10010100_10010101_0;
      patterns[407] = 25'b00000001_10010101_10010110_0;
      patterns[408] = 25'b00000001_10010110_10010111_0;
      patterns[409] = 25'b00000001_10010111_10011000_0;
      patterns[410] = 25'b00000001_10011000_10011001_0;
      patterns[411] = 25'b00000001_10011001_10011010_0;
      patterns[412] = 25'b00000001_10011010_10011011_0;
      patterns[413] = 25'b00000001_10011011_10011100_0;
      patterns[414] = 25'b00000001_10011100_10011101_0;
      patterns[415] = 25'b00000001_10011101_10011110_0;
      patterns[416] = 25'b00000001_10011110_10011111_0;
      patterns[417] = 25'b00000001_10011111_10100000_0;
      patterns[418] = 25'b00000001_10100000_10100001_0;
      patterns[419] = 25'b00000001_10100001_10100010_0;
      patterns[420] = 25'b00000001_10100010_10100011_0;
      patterns[421] = 25'b00000001_10100011_10100100_0;
      patterns[422] = 25'b00000001_10100100_10100101_0;
      patterns[423] = 25'b00000001_10100101_10100110_0;
      patterns[424] = 25'b00000001_10100110_10100111_0;
      patterns[425] = 25'b00000001_10100111_10101000_0;
      patterns[426] = 25'b00000001_10101000_10101001_0;
      patterns[427] = 25'b00000001_10101001_10101010_0;
      patterns[428] = 25'b00000001_10101010_10101011_0;
      patterns[429] = 25'b00000001_10101011_10101100_0;
      patterns[430] = 25'b00000001_10101100_10101101_0;
      patterns[431] = 25'b00000001_10101101_10101110_0;
      patterns[432] = 25'b00000001_10101110_10101111_0;
      patterns[433] = 25'b00000001_10101111_10110000_0;
      patterns[434] = 25'b00000001_10110000_10110001_0;
      patterns[435] = 25'b00000001_10110001_10110010_0;
      patterns[436] = 25'b00000001_10110010_10110011_0;
      patterns[437] = 25'b00000001_10110011_10110100_0;
      patterns[438] = 25'b00000001_10110100_10110101_0;
      patterns[439] = 25'b00000001_10110101_10110110_0;
      patterns[440] = 25'b00000001_10110110_10110111_0;
      patterns[441] = 25'b00000001_10110111_10111000_0;
      patterns[442] = 25'b00000001_10111000_10111001_0;
      patterns[443] = 25'b00000001_10111001_10111010_0;
      patterns[444] = 25'b00000001_10111010_10111011_0;
      patterns[445] = 25'b00000001_10111011_10111100_0;
      patterns[446] = 25'b00000001_10111100_10111101_0;
      patterns[447] = 25'b00000001_10111101_10111110_0;
      patterns[448] = 25'b00000001_10111110_10111111_0;
      patterns[449] = 25'b00000001_10111111_11000000_0;
      patterns[450] = 25'b00000001_11000000_11000001_0;
      patterns[451] = 25'b00000001_11000001_11000010_0;
      patterns[452] = 25'b00000001_11000010_11000011_0;
      patterns[453] = 25'b00000001_11000011_11000100_0;
      patterns[454] = 25'b00000001_11000100_11000101_0;
      patterns[455] = 25'b00000001_11000101_11000110_0;
      patterns[456] = 25'b00000001_11000110_11000111_0;
      patterns[457] = 25'b00000001_11000111_11001000_0;
      patterns[458] = 25'b00000001_11001000_11001001_0;
      patterns[459] = 25'b00000001_11001001_11001010_0;
      patterns[460] = 25'b00000001_11001010_11001011_0;
      patterns[461] = 25'b00000001_11001011_11001100_0;
      patterns[462] = 25'b00000001_11001100_11001101_0;
      patterns[463] = 25'b00000001_11001101_11001110_0;
      patterns[464] = 25'b00000001_11001110_11001111_0;
      patterns[465] = 25'b00000001_11001111_11010000_0;
      patterns[466] = 25'b00000001_11010000_11010001_0;
      patterns[467] = 25'b00000001_11010001_11010010_0;
      patterns[468] = 25'b00000001_11010010_11010011_0;
      patterns[469] = 25'b00000001_11010011_11010100_0;
      patterns[470] = 25'b00000001_11010100_11010101_0;
      patterns[471] = 25'b00000001_11010101_11010110_0;
      patterns[472] = 25'b00000001_11010110_11010111_0;
      patterns[473] = 25'b00000001_11010111_11011000_0;
      patterns[474] = 25'b00000001_11011000_11011001_0;
      patterns[475] = 25'b00000001_11011001_11011010_0;
      patterns[476] = 25'b00000001_11011010_11011011_0;
      patterns[477] = 25'b00000001_11011011_11011100_0;
      patterns[478] = 25'b00000001_11011100_11011101_0;
      patterns[479] = 25'b00000001_11011101_11011110_0;
      patterns[480] = 25'b00000001_11011110_11011111_0;
      patterns[481] = 25'b00000001_11011111_11100000_0;
      patterns[482] = 25'b00000001_11100000_11100001_0;
      patterns[483] = 25'b00000001_11100001_11100010_0;
      patterns[484] = 25'b00000001_11100010_11100011_0;
      patterns[485] = 25'b00000001_11100011_11100100_0;
      patterns[486] = 25'b00000001_11100100_11100101_0;
      patterns[487] = 25'b00000001_11100101_11100110_0;
      patterns[488] = 25'b00000001_11100110_11100111_0;
      patterns[489] = 25'b00000001_11100111_11101000_0;
      patterns[490] = 25'b00000001_11101000_11101001_0;
      patterns[491] = 25'b00000001_11101001_11101010_0;
      patterns[492] = 25'b00000001_11101010_11101011_0;
      patterns[493] = 25'b00000001_11101011_11101100_0;
      patterns[494] = 25'b00000001_11101100_11101101_0;
      patterns[495] = 25'b00000001_11101101_11101110_0;
      patterns[496] = 25'b00000001_11101110_11101111_0;
      patterns[497] = 25'b00000001_11101111_11110000_0;
      patterns[498] = 25'b00000001_11110000_11110001_0;
      patterns[499] = 25'b00000001_11110001_11110010_0;
      patterns[500] = 25'b00000001_11110010_11110011_0;
      patterns[501] = 25'b00000001_11110011_11110100_0;
      patterns[502] = 25'b00000001_11110100_11110101_0;
      patterns[503] = 25'b00000001_11110101_11110110_0;
      patterns[504] = 25'b00000001_11110110_11110111_0;
      patterns[505] = 25'b00000001_11110111_11111000_0;
      patterns[506] = 25'b00000001_11111000_11111001_0;
      patterns[507] = 25'b00000001_11111001_11111010_0;
      patterns[508] = 25'b00000001_11111010_11111011_0;
      patterns[509] = 25'b00000001_11111011_11111100_0;
      patterns[510] = 25'b00000001_11111100_11111101_0;
      patterns[511] = 25'b00000001_11111101_11111110_0;
      patterns[512] = 25'b00000001_11111110_11111111_0;
      patterns[513] = 25'b00000001_11111111_00000000_1;
      patterns[514] = 25'b00000010_00000000_00000010_0;
      patterns[515] = 25'b00000010_00000001_00000011_0;
      patterns[516] = 25'b00000010_00000010_00000100_0;
      patterns[517] = 25'b00000010_00000011_00000101_0;
      patterns[518] = 25'b00000010_00000100_00000110_0;
      patterns[519] = 25'b00000010_00000101_00000111_0;
      patterns[520] = 25'b00000010_00000110_00001000_0;
      patterns[521] = 25'b00000010_00000111_00001001_0;
      patterns[522] = 25'b00000010_00001000_00001010_0;
      patterns[523] = 25'b00000010_00001001_00001011_0;
      patterns[524] = 25'b00000010_00001010_00001100_0;
      patterns[525] = 25'b00000010_00001011_00001101_0;
      patterns[526] = 25'b00000010_00001100_00001110_0;
      patterns[527] = 25'b00000010_00001101_00001111_0;
      patterns[528] = 25'b00000010_00001110_00010000_0;
      patterns[529] = 25'b00000010_00001111_00010001_0;
      patterns[530] = 25'b00000010_00010000_00010010_0;
      patterns[531] = 25'b00000010_00010001_00010011_0;
      patterns[532] = 25'b00000010_00010010_00010100_0;
      patterns[533] = 25'b00000010_00010011_00010101_0;
      patterns[534] = 25'b00000010_00010100_00010110_0;
      patterns[535] = 25'b00000010_00010101_00010111_0;
      patterns[536] = 25'b00000010_00010110_00011000_0;
      patterns[537] = 25'b00000010_00010111_00011001_0;
      patterns[538] = 25'b00000010_00011000_00011010_0;
      patterns[539] = 25'b00000010_00011001_00011011_0;
      patterns[540] = 25'b00000010_00011010_00011100_0;
      patterns[541] = 25'b00000010_00011011_00011101_0;
      patterns[542] = 25'b00000010_00011100_00011110_0;
      patterns[543] = 25'b00000010_00011101_00011111_0;
      patterns[544] = 25'b00000010_00011110_00100000_0;
      patterns[545] = 25'b00000010_00011111_00100001_0;
      patterns[546] = 25'b00000010_00100000_00100010_0;
      patterns[547] = 25'b00000010_00100001_00100011_0;
      patterns[548] = 25'b00000010_00100010_00100100_0;
      patterns[549] = 25'b00000010_00100011_00100101_0;
      patterns[550] = 25'b00000010_00100100_00100110_0;
      patterns[551] = 25'b00000010_00100101_00100111_0;
      patterns[552] = 25'b00000010_00100110_00101000_0;
      patterns[553] = 25'b00000010_00100111_00101001_0;
      patterns[554] = 25'b00000010_00101000_00101010_0;
      patterns[555] = 25'b00000010_00101001_00101011_0;
      patterns[556] = 25'b00000010_00101010_00101100_0;
      patterns[557] = 25'b00000010_00101011_00101101_0;
      patterns[558] = 25'b00000010_00101100_00101110_0;
      patterns[559] = 25'b00000010_00101101_00101111_0;
      patterns[560] = 25'b00000010_00101110_00110000_0;
      patterns[561] = 25'b00000010_00101111_00110001_0;
      patterns[562] = 25'b00000010_00110000_00110010_0;
      patterns[563] = 25'b00000010_00110001_00110011_0;
      patterns[564] = 25'b00000010_00110010_00110100_0;
      patterns[565] = 25'b00000010_00110011_00110101_0;
      patterns[566] = 25'b00000010_00110100_00110110_0;
      patterns[567] = 25'b00000010_00110101_00110111_0;
      patterns[568] = 25'b00000010_00110110_00111000_0;
      patterns[569] = 25'b00000010_00110111_00111001_0;
      patterns[570] = 25'b00000010_00111000_00111010_0;
      patterns[571] = 25'b00000010_00111001_00111011_0;
      patterns[572] = 25'b00000010_00111010_00111100_0;
      patterns[573] = 25'b00000010_00111011_00111101_0;
      patterns[574] = 25'b00000010_00111100_00111110_0;
      patterns[575] = 25'b00000010_00111101_00111111_0;
      patterns[576] = 25'b00000010_00111110_01000000_0;
      patterns[577] = 25'b00000010_00111111_01000001_0;
      patterns[578] = 25'b00000010_01000000_01000010_0;
      patterns[579] = 25'b00000010_01000001_01000011_0;
      patterns[580] = 25'b00000010_01000010_01000100_0;
      patterns[581] = 25'b00000010_01000011_01000101_0;
      patterns[582] = 25'b00000010_01000100_01000110_0;
      patterns[583] = 25'b00000010_01000101_01000111_0;
      patterns[584] = 25'b00000010_01000110_01001000_0;
      patterns[585] = 25'b00000010_01000111_01001001_0;
      patterns[586] = 25'b00000010_01001000_01001010_0;
      patterns[587] = 25'b00000010_01001001_01001011_0;
      patterns[588] = 25'b00000010_01001010_01001100_0;
      patterns[589] = 25'b00000010_01001011_01001101_0;
      patterns[590] = 25'b00000010_01001100_01001110_0;
      patterns[591] = 25'b00000010_01001101_01001111_0;
      patterns[592] = 25'b00000010_01001110_01010000_0;
      patterns[593] = 25'b00000010_01001111_01010001_0;
      patterns[594] = 25'b00000010_01010000_01010010_0;
      patterns[595] = 25'b00000010_01010001_01010011_0;
      patterns[596] = 25'b00000010_01010010_01010100_0;
      patterns[597] = 25'b00000010_01010011_01010101_0;
      patterns[598] = 25'b00000010_01010100_01010110_0;
      patterns[599] = 25'b00000010_01010101_01010111_0;
      patterns[600] = 25'b00000010_01010110_01011000_0;
      patterns[601] = 25'b00000010_01010111_01011001_0;
      patterns[602] = 25'b00000010_01011000_01011010_0;
      patterns[603] = 25'b00000010_01011001_01011011_0;
      patterns[604] = 25'b00000010_01011010_01011100_0;
      patterns[605] = 25'b00000010_01011011_01011101_0;
      patterns[606] = 25'b00000010_01011100_01011110_0;
      patterns[607] = 25'b00000010_01011101_01011111_0;
      patterns[608] = 25'b00000010_01011110_01100000_0;
      patterns[609] = 25'b00000010_01011111_01100001_0;
      patterns[610] = 25'b00000010_01100000_01100010_0;
      patterns[611] = 25'b00000010_01100001_01100011_0;
      patterns[612] = 25'b00000010_01100010_01100100_0;
      patterns[613] = 25'b00000010_01100011_01100101_0;
      patterns[614] = 25'b00000010_01100100_01100110_0;
      patterns[615] = 25'b00000010_01100101_01100111_0;
      patterns[616] = 25'b00000010_01100110_01101000_0;
      patterns[617] = 25'b00000010_01100111_01101001_0;
      patterns[618] = 25'b00000010_01101000_01101010_0;
      patterns[619] = 25'b00000010_01101001_01101011_0;
      patterns[620] = 25'b00000010_01101010_01101100_0;
      patterns[621] = 25'b00000010_01101011_01101101_0;
      patterns[622] = 25'b00000010_01101100_01101110_0;
      patterns[623] = 25'b00000010_01101101_01101111_0;
      patterns[624] = 25'b00000010_01101110_01110000_0;
      patterns[625] = 25'b00000010_01101111_01110001_0;
      patterns[626] = 25'b00000010_01110000_01110010_0;
      patterns[627] = 25'b00000010_01110001_01110011_0;
      patterns[628] = 25'b00000010_01110010_01110100_0;
      patterns[629] = 25'b00000010_01110011_01110101_0;
      patterns[630] = 25'b00000010_01110100_01110110_0;
      patterns[631] = 25'b00000010_01110101_01110111_0;
      patterns[632] = 25'b00000010_01110110_01111000_0;
      patterns[633] = 25'b00000010_01110111_01111001_0;
      patterns[634] = 25'b00000010_01111000_01111010_0;
      patterns[635] = 25'b00000010_01111001_01111011_0;
      patterns[636] = 25'b00000010_01111010_01111100_0;
      patterns[637] = 25'b00000010_01111011_01111101_0;
      patterns[638] = 25'b00000010_01111100_01111110_0;
      patterns[639] = 25'b00000010_01111101_01111111_0;
      patterns[640] = 25'b00000010_01111110_10000000_0;
      patterns[641] = 25'b00000010_01111111_10000001_0;
      patterns[642] = 25'b00000010_10000000_10000010_0;
      patterns[643] = 25'b00000010_10000001_10000011_0;
      patterns[644] = 25'b00000010_10000010_10000100_0;
      patterns[645] = 25'b00000010_10000011_10000101_0;
      patterns[646] = 25'b00000010_10000100_10000110_0;
      patterns[647] = 25'b00000010_10000101_10000111_0;
      patterns[648] = 25'b00000010_10000110_10001000_0;
      patterns[649] = 25'b00000010_10000111_10001001_0;
      patterns[650] = 25'b00000010_10001000_10001010_0;
      patterns[651] = 25'b00000010_10001001_10001011_0;
      patterns[652] = 25'b00000010_10001010_10001100_0;
      patterns[653] = 25'b00000010_10001011_10001101_0;
      patterns[654] = 25'b00000010_10001100_10001110_0;
      patterns[655] = 25'b00000010_10001101_10001111_0;
      patterns[656] = 25'b00000010_10001110_10010000_0;
      patterns[657] = 25'b00000010_10001111_10010001_0;
      patterns[658] = 25'b00000010_10010000_10010010_0;
      patterns[659] = 25'b00000010_10010001_10010011_0;
      patterns[660] = 25'b00000010_10010010_10010100_0;
      patterns[661] = 25'b00000010_10010011_10010101_0;
      patterns[662] = 25'b00000010_10010100_10010110_0;
      patterns[663] = 25'b00000010_10010101_10010111_0;
      patterns[664] = 25'b00000010_10010110_10011000_0;
      patterns[665] = 25'b00000010_10010111_10011001_0;
      patterns[666] = 25'b00000010_10011000_10011010_0;
      patterns[667] = 25'b00000010_10011001_10011011_0;
      patterns[668] = 25'b00000010_10011010_10011100_0;
      patterns[669] = 25'b00000010_10011011_10011101_0;
      patterns[670] = 25'b00000010_10011100_10011110_0;
      patterns[671] = 25'b00000010_10011101_10011111_0;
      patterns[672] = 25'b00000010_10011110_10100000_0;
      patterns[673] = 25'b00000010_10011111_10100001_0;
      patterns[674] = 25'b00000010_10100000_10100010_0;
      patterns[675] = 25'b00000010_10100001_10100011_0;
      patterns[676] = 25'b00000010_10100010_10100100_0;
      patterns[677] = 25'b00000010_10100011_10100101_0;
      patterns[678] = 25'b00000010_10100100_10100110_0;
      patterns[679] = 25'b00000010_10100101_10100111_0;
      patterns[680] = 25'b00000010_10100110_10101000_0;
      patterns[681] = 25'b00000010_10100111_10101001_0;
      patterns[682] = 25'b00000010_10101000_10101010_0;
      patterns[683] = 25'b00000010_10101001_10101011_0;
      patterns[684] = 25'b00000010_10101010_10101100_0;
      patterns[685] = 25'b00000010_10101011_10101101_0;
      patterns[686] = 25'b00000010_10101100_10101110_0;
      patterns[687] = 25'b00000010_10101101_10101111_0;
      patterns[688] = 25'b00000010_10101110_10110000_0;
      patterns[689] = 25'b00000010_10101111_10110001_0;
      patterns[690] = 25'b00000010_10110000_10110010_0;
      patterns[691] = 25'b00000010_10110001_10110011_0;
      patterns[692] = 25'b00000010_10110010_10110100_0;
      patterns[693] = 25'b00000010_10110011_10110101_0;
      patterns[694] = 25'b00000010_10110100_10110110_0;
      patterns[695] = 25'b00000010_10110101_10110111_0;
      patterns[696] = 25'b00000010_10110110_10111000_0;
      patterns[697] = 25'b00000010_10110111_10111001_0;
      patterns[698] = 25'b00000010_10111000_10111010_0;
      patterns[699] = 25'b00000010_10111001_10111011_0;
      patterns[700] = 25'b00000010_10111010_10111100_0;
      patterns[701] = 25'b00000010_10111011_10111101_0;
      patterns[702] = 25'b00000010_10111100_10111110_0;
      patterns[703] = 25'b00000010_10111101_10111111_0;
      patterns[704] = 25'b00000010_10111110_11000000_0;
      patterns[705] = 25'b00000010_10111111_11000001_0;
      patterns[706] = 25'b00000010_11000000_11000010_0;
      patterns[707] = 25'b00000010_11000001_11000011_0;
      patterns[708] = 25'b00000010_11000010_11000100_0;
      patterns[709] = 25'b00000010_11000011_11000101_0;
      patterns[710] = 25'b00000010_11000100_11000110_0;
      patterns[711] = 25'b00000010_11000101_11000111_0;
      patterns[712] = 25'b00000010_11000110_11001000_0;
      patterns[713] = 25'b00000010_11000111_11001001_0;
      patterns[714] = 25'b00000010_11001000_11001010_0;
      patterns[715] = 25'b00000010_11001001_11001011_0;
      patterns[716] = 25'b00000010_11001010_11001100_0;
      patterns[717] = 25'b00000010_11001011_11001101_0;
      patterns[718] = 25'b00000010_11001100_11001110_0;
      patterns[719] = 25'b00000010_11001101_11001111_0;
      patterns[720] = 25'b00000010_11001110_11010000_0;
      patterns[721] = 25'b00000010_11001111_11010001_0;
      patterns[722] = 25'b00000010_11010000_11010010_0;
      patterns[723] = 25'b00000010_11010001_11010011_0;
      patterns[724] = 25'b00000010_11010010_11010100_0;
      patterns[725] = 25'b00000010_11010011_11010101_0;
      patterns[726] = 25'b00000010_11010100_11010110_0;
      patterns[727] = 25'b00000010_11010101_11010111_0;
      patterns[728] = 25'b00000010_11010110_11011000_0;
      patterns[729] = 25'b00000010_11010111_11011001_0;
      patterns[730] = 25'b00000010_11011000_11011010_0;
      patterns[731] = 25'b00000010_11011001_11011011_0;
      patterns[732] = 25'b00000010_11011010_11011100_0;
      patterns[733] = 25'b00000010_11011011_11011101_0;
      patterns[734] = 25'b00000010_11011100_11011110_0;
      patterns[735] = 25'b00000010_11011101_11011111_0;
      patterns[736] = 25'b00000010_11011110_11100000_0;
      patterns[737] = 25'b00000010_11011111_11100001_0;
      patterns[738] = 25'b00000010_11100000_11100010_0;
      patterns[739] = 25'b00000010_11100001_11100011_0;
      patterns[740] = 25'b00000010_11100010_11100100_0;
      patterns[741] = 25'b00000010_11100011_11100101_0;
      patterns[742] = 25'b00000010_11100100_11100110_0;
      patterns[743] = 25'b00000010_11100101_11100111_0;
      patterns[744] = 25'b00000010_11100110_11101000_0;
      patterns[745] = 25'b00000010_11100111_11101001_0;
      patterns[746] = 25'b00000010_11101000_11101010_0;
      patterns[747] = 25'b00000010_11101001_11101011_0;
      patterns[748] = 25'b00000010_11101010_11101100_0;
      patterns[749] = 25'b00000010_11101011_11101101_0;
      patterns[750] = 25'b00000010_11101100_11101110_0;
      patterns[751] = 25'b00000010_11101101_11101111_0;
      patterns[752] = 25'b00000010_11101110_11110000_0;
      patterns[753] = 25'b00000010_11101111_11110001_0;
      patterns[754] = 25'b00000010_11110000_11110010_0;
      patterns[755] = 25'b00000010_11110001_11110011_0;
      patterns[756] = 25'b00000010_11110010_11110100_0;
      patterns[757] = 25'b00000010_11110011_11110101_0;
      patterns[758] = 25'b00000010_11110100_11110110_0;
      patterns[759] = 25'b00000010_11110101_11110111_0;
      patterns[760] = 25'b00000010_11110110_11111000_0;
      patterns[761] = 25'b00000010_11110111_11111001_0;
      patterns[762] = 25'b00000010_11111000_11111010_0;
      patterns[763] = 25'b00000010_11111001_11111011_0;
      patterns[764] = 25'b00000010_11111010_11111100_0;
      patterns[765] = 25'b00000010_11111011_11111101_0;
      patterns[766] = 25'b00000010_11111100_11111110_0;
      patterns[767] = 25'b00000010_11111101_11111111_0;
      patterns[768] = 25'b00000010_11111110_00000000_1;
      patterns[769] = 25'b00000010_11111111_00000001_1;
      patterns[770] = 25'b00000011_00000000_00000011_0;
      patterns[771] = 25'b00000011_00000001_00000100_0;
      patterns[772] = 25'b00000011_00000010_00000101_0;
      patterns[773] = 25'b00000011_00000011_00000110_0;
      patterns[774] = 25'b00000011_00000100_00000111_0;
      patterns[775] = 25'b00000011_00000101_00001000_0;
      patterns[776] = 25'b00000011_00000110_00001001_0;
      patterns[777] = 25'b00000011_00000111_00001010_0;
      patterns[778] = 25'b00000011_00001000_00001011_0;
      patterns[779] = 25'b00000011_00001001_00001100_0;
      patterns[780] = 25'b00000011_00001010_00001101_0;
      patterns[781] = 25'b00000011_00001011_00001110_0;
      patterns[782] = 25'b00000011_00001100_00001111_0;
      patterns[783] = 25'b00000011_00001101_00010000_0;
      patterns[784] = 25'b00000011_00001110_00010001_0;
      patterns[785] = 25'b00000011_00001111_00010010_0;
      patterns[786] = 25'b00000011_00010000_00010011_0;
      patterns[787] = 25'b00000011_00010001_00010100_0;
      patterns[788] = 25'b00000011_00010010_00010101_0;
      patterns[789] = 25'b00000011_00010011_00010110_0;
      patterns[790] = 25'b00000011_00010100_00010111_0;
      patterns[791] = 25'b00000011_00010101_00011000_0;
      patterns[792] = 25'b00000011_00010110_00011001_0;
      patterns[793] = 25'b00000011_00010111_00011010_0;
      patterns[794] = 25'b00000011_00011000_00011011_0;
      patterns[795] = 25'b00000011_00011001_00011100_0;
      patterns[796] = 25'b00000011_00011010_00011101_0;
      patterns[797] = 25'b00000011_00011011_00011110_0;
      patterns[798] = 25'b00000011_00011100_00011111_0;
      patterns[799] = 25'b00000011_00011101_00100000_0;
      patterns[800] = 25'b00000011_00011110_00100001_0;
      patterns[801] = 25'b00000011_00011111_00100010_0;
      patterns[802] = 25'b00000011_00100000_00100011_0;
      patterns[803] = 25'b00000011_00100001_00100100_0;
      patterns[804] = 25'b00000011_00100010_00100101_0;
      patterns[805] = 25'b00000011_00100011_00100110_0;
      patterns[806] = 25'b00000011_00100100_00100111_0;
      patterns[807] = 25'b00000011_00100101_00101000_0;
      patterns[808] = 25'b00000011_00100110_00101001_0;
      patterns[809] = 25'b00000011_00100111_00101010_0;
      patterns[810] = 25'b00000011_00101000_00101011_0;
      patterns[811] = 25'b00000011_00101001_00101100_0;
      patterns[812] = 25'b00000011_00101010_00101101_0;
      patterns[813] = 25'b00000011_00101011_00101110_0;
      patterns[814] = 25'b00000011_00101100_00101111_0;
      patterns[815] = 25'b00000011_00101101_00110000_0;
      patterns[816] = 25'b00000011_00101110_00110001_0;
      patterns[817] = 25'b00000011_00101111_00110010_0;
      patterns[818] = 25'b00000011_00110000_00110011_0;
      patterns[819] = 25'b00000011_00110001_00110100_0;
      patterns[820] = 25'b00000011_00110010_00110101_0;
      patterns[821] = 25'b00000011_00110011_00110110_0;
      patterns[822] = 25'b00000011_00110100_00110111_0;
      patterns[823] = 25'b00000011_00110101_00111000_0;
      patterns[824] = 25'b00000011_00110110_00111001_0;
      patterns[825] = 25'b00000011_00110111_00111010_0;
      patterns[826] = 25'b00000011_00111000_00111011_0;
      patterns[827] = 25'b00000011_00111001_00111100_0;
      patterns[828] = 25'b00000011_00111010_00111101_0;
      patterns[829] = 25'b00000011_00111011_00111110_0;
      patterns[830] = 25'b00000011_00111100_00111111_0;
      patterns[831] = 25'b00000011_00111101_01000000_0;
      patterns[832] = 25'b00000011_00111110_01000001_0;
      patterns[833] = 25'b00000011_00111111_01000010_0;
      patterns[834] = 25'b00000011_01000000_01000011_0;
      patterns[835] = 25'b00000011_01000001_01000100_0;
      patterns[836] = 25'b00000011_01000010_01000101_0;
      patterns[837] = 25'b00000011_01000011_01000110_0;
      patterns[838] = 25'b00000011_01000100_01000111_0;
      patterns[839] = 25'b00000011_01000101_01001000_0;
      patterns[840] = 25'b00000011_01000110_01001001_0;
      patterns[841] = 25'b00000011_01000111_01001010_0;
      patterns[842] = 25'b00000011_01001000_01001011_0;
      patterns[843] = 25'b00000011_01001001_01001100_0;
      patterns[844] = 25'b00000011_01001010_01001101_0;
      patterns[845] = 25'b00000011_01001011_01001110_0;
      patterns[846] = 25'b00000011_01001100_01001111_0;
      patterns[847] = 25'b00000011_01001101_01010000_0;
      patterns[848] = 25'b00000011_01001110_01010001_0;
      patterns[849] = 25'b00000011_01001111_01010010_0;
      patterns[850] = 25'b00000011_01010000_01010011_0;
      patterns[851] = 25'b00000011_01010001_01010100_0;
      patterns[852] = 25'b00000011_01010010_01010101_0;
      patterns[853] = 25'b00000011_01010011_01010110_0;
      patterns[854] = 25'b00000011_01010100_01010111_0;
      patterns[855] = 25'b00000011_01010101_01011000_0;
      patterns[856] = 25'b00000011_01010110_01011001_0;
      patterns[857] = 25'b00000011_01010111_01011010_0;
      patterns[858] = 25'b00000011_01011000_01011011_0;
      patterns[859] = 25'b00000011_01011001_01011100_0;
      patterns[860] = 25'b00000011_01011010_01011101_0;
      patterns[861] = 25'b00000011_01011011_01011110_0;
      patterns[862] = 25'b00000011_01011100_01011111_0;
      patterns[863] = 25'b00000011_01011101_01100000_0;
      patterns[864] = 25'b00000011_01011110_01100001_0;
      patterns[865] = 25'b00000011_01011111_01100010_0;
      patterns[866] = 25'b00000011_01100000_01100011_0;
      patterns[867] = 25'b00000011_01100001_01100100_0;
      patterns[868] = 25'b00000011_01100010_01100101_0;
      patterns[869] = 25'b00000011_01100011_01100110_0;
      patterns[870] = 25'b00000011_01100100_01100111_0;
      patterns[871] = 25'b00000011_01100101_01101000_0;
      patterns[872] = 25'b00000011_01100110_01101001_0;
      patterns[873] = 25'b00000011_01100111_01101010_0;
      patterns[874] = 25'b00000011_01101000_01101011_0;
      patterns[875] = 25'b00000011_01101001_01101100_0;
      patterns[876] = 25'b00000011_01101010_01101101_0;
      patterns[877] = 25'b00000011_01101011_01101110_0;
      patterns[878] = 25'b00000011_01101100_01101111_0;
      patterns[879] = 25'b00000011_01101101_01110000_0;
      patterns[880] = 25'b00000011_01101110_01110001_0;
      patterns[881] = 25'b00000011_01101111_01110010_0;
      patterns[882] = 25'b00000011_01110000_01110011_0;
      patterns[883] = 25'b00000011_01110001_01110100_0;
      patterns[884] = 25'b00000011_01110010_01110101_0;
      patterns[885] = 25'b00000011_01110011_01110110_0;
      patterns[886] = 25'b00000011_01110100_01110111_0;
      patterns[887] = 25'b00000011_01110101_01111000_0;
      patterns[888] = 25'b00000011_01110110_01111001_0;
      patterns[889] = 25'b00000011_01110111_01111010_0;
      patterns[890] = 25'b00000011_01111000_01111011_0;
      patterns[891] = 25'b00000011_01111001_01111100_0;
      patterns[892] = 25'b00000011_01111010_01111101_0;
      patterns[893] = 25'b00000011_01111011_01111110_0;
      patterns[894] = 25'b00000011_01111100_01111111_0;
      patterns[895] = 25'b00000011_01111101_10000000_0;
      patterns[896] = 25'b00000011_01111110_10000001_0;
      patterns[897] = 25'b00000011_01111111_10000010_0;
      patterns[898] = 25'b00000011_10000000_10000011_0;
      patterns[899] = 25'b00000011_10000001_10000100_0;
      patterns[900] = 25'b00000011_10000010_10000101_0;
      patterns[901] = 25'b00000011_10000011_10000110_0;
      patterns[902] = 25'b00000011_10000100_10000111_0;
      patterns[903] = 25'b00000011_10000101_10001000_0;
      patterns[904] = 25'b00000011_10000110_10001001_0;
      patterns[905] = 25'b00000011_10000111_10001010_0;
      patterns[906] = 25'b00000011_10001000_10001011_0;
      patterns[907] = 25'b00000011_10001001_10001100_0;
      patterns[908] = 25'b00000011_10001010_10001101_0;
      patterns[909] = 25'b00000011_10001011_10001110_0;
      patterns[910] = 25'b00000011_10001100_10001111_0;
      patterns[911] = 25'b00000011_10001101_10010000_0;
      patterns[912] = 25'b00000011_10001110_10010001_0;
      patterns[913] = 25'b00000011_10001111_10010010_0;
      patterns[914] = 25'b00000011_10010000_10010011_0;
      patterns[915] = 25'b00000011_10010001_10010100_0;
      patterns[916] = 25'b00000011_10010010_10010101_0;
      patterns[917] = 25'b00000011_10010011_10010110_0;
      patterns[918] = 25'b00000011_10010100_10010111_0;
      patterns[919] = 25'b00000011_10010101_10011000_0;
      patterns[920] = 25'b00000011_10010110_10011001_0;
      patterns[921] = 25'b00000011_10010111_10011010_0;
      patterns[922] = 25'b00000011_10011000_10011011_0;
      patterns[923] = 25'b00000011_10011001_10011100_0;
      patterns[924] = 25'b00000011_10011010_10011101_0;
      patterns[925] = 25'b00000011_10011011_10011110_0;
      patterns[926] = 25'b00000011_10011100_10011111_0;
      patterns[927] = 25'b00000011_10011101_10100000_0;
      patterns[928] = 25'b00000011_10011110_10100001_0;
      patterns[929] = 25'b00000011_10011111_10100010_0;
      patterns[930] = 25'b00000011_10100000_10100011_0;
      patterns[931] = 25'b00000011_10100001_10100100_0;
      patterns[932] = 25'b00000011_10100010_10100101_0;
      patterns[933] = 25'b00000011_10100011_10100110_0;
      patterns[934] = 25'b00000011_10100100_10100111_0;
      patterns[935] = 25'b00000011_10100101_10101000_0;
      patterns[936] = 25'b00000011_10100110_10101001_0;
      patterns[937] = 25'b00000011_10100111_10101010_0;
      patterns[938] = 25'b00000011_10101000_10101011_0;
      patterns[939] = 25'b00000011_10101001_10101100_0;
      patterns[940] = 25'b00000011_10101010_10101101_0;
      patterns[941] = 25'b00000011_10101011_10101110_0;
      patterns[942] = 25'b00000011_10101100_10101111_0;
      patterns[943] = 25'b00000011_10101101_10110000_0;
      patterns[944] = 25'b00000011_10101110_10110001_0;
      patterns[945] = 25'b00000011_10101111_10110010_0;
      patterns[946] = 25'b00000011_10110000_10110011_0;
      patterns[947] = 25'b00000011_10110001_10110100_0;
      patterns[948] = 25'b00000011_10110010_10110101_0;
      patterns[949] = 25'b00000011_10110011_10110110_0;
      patterns[950] = 25'b00000011_10110100_10110111_0;
      patterns[951] = 25'b00000011_10110101_10111000_0;
      patterns[952] = 25'b00000011_10110110_10111001_0;
      patterns[953] = 25'b00000011_10110111_10111010_0;
      patterns[954] = 25'b00000011_10111000_10111011_0;
      patterns[955] = 25'b00000011_10111001_10111100_0;
      patterns[956] = 25'b00000011_10111010_10111101_0;
      patterns[957] = 25'b00000011_10111011_10111110_0;
      patterns[958] = 25'b00000011_10111100_10111111_0;
      patterns[959] = 25'b00000011_10111101_11000000_0;
      patterns[960] = 25'b00000011_10111110_11000001_0;
      patterns[961] = 25'b00000011_10111111_11000010_0;
      patterns[962] = 25'b00000011_11000000_11000011_0;
      patterns[963] = 25'b00000011_11000001_11000100_0;
      patterns[964] = 25'b00000011_11000010_11000101_0;
      patterns[965] = 25'b00000011_11000011_11000110_0;
      patterns[966] = 25'b00000011_11000100_11000111_0;
      patterns[967] = 25'b00000011_11000101_11001000_0;
      patterns[968] = 25'b00000011_11000110_11001001_0;
      patterns[969] = 25'b00000011_11000111_11001010_0;
      patterns[970] = 25'b00000011_11001000_11001011_0;
      patterns[971] = 25'b00000011_11001001_11001100_0;
      patterns[972] = 25'b00000011_11001010_11001101_0;
      patterns[973] = 25'b00000011_11001011_11001110_0;
      patterns[974] = 25'b00000011_11001100_11001111_0;
      patterns[975] = 25'b00000011_11001101_11010000_0;
      patterns[976] = 25'b00000011_11001110_11010001_0;
      patterns[977] = 25'b00000011_11001111_11010010_0;
      patterns[978] = 25'b00000011_11010000_11010011_0;
      patterns[979] = 25'b00000011_11010001_11010100_0;
      patterns[980] = 25'b00000011_11010010_11010101_0;
      patterns[981] = 25'b00000011_11010011_11010110_0;
      patterns[982] = 25'b00000011_11010100_11010111_0;
      patterns[983] = 25'b00000011_11010101_11011000_0;
      patterns[984] = 25'b00000011_11010110_11011001_0;
      patterns[985] = 25'b00000011_11010111_11011010_0;
      patterns[986] = 25'b00000011_11011000_11011011_0;
      patterns[987] = 25'b00000011_11011001_11011100_0;
      patterns[988] = 25'b00000011_11011010_11011101_0;
      patterns[989] = 25'b00000011_11011011_11011110_0;
      patterns[990] = 25'b00000011_11011100_11011111_0;
      patterns[991] = 25'b00000011_11011101_11100000_0;
      patterns[992] = 25'b00000011_11011110_11100001_0;
      patterns[993] = 25'b00000011_11011111_11100010_0;
      patterns[994] = 25'b00000011_11100000_11100011_0;
      patterns[995] = 25'b00000011_11100001_11100100_0;
      patterns[996] = 25'b00000011_11100010_11100101_0;
      patterns[997] = 25'b00000011_11100011_11100110_0;
      patterns[998] = 25'b00000011_11100100_11100111_0;
      patterns[999] = 25'b00000011_11100101_11101000_0;
      patterns[1000] = 25'b00000011_11100110_11101001_0;
      patterns[1001] = 25'b00000011_11100111_11101010_0;
      patterns[1002] = 25'b00000011_11101000_11101011_0;
      patterns[1003] = 25'b00000011_11101001_11101100_0;
      patterns[1004] = 25'b00000011_11101010_11101101_0;
      patterns[1005] = 25'b00000011_11101011_11101110_0;
      patterns[1006] = 25'b00000011_11101100_11101111_0;
      patterns[1007] = 25'b00000011_11101101_11110000_0;
      patterns[1008] = 25'b00000011_11101110_11110001_0;
      patterns[1009] = 25'b00000011_11101111_11110010_0;
      patterns[1010] = 25'b00000011_11110000_11110011_0;
      patterns[1011] = 25'b00000011_11110001_11110100_0;
      patterns[1012] = 25'b00000011_11110010_11110101_0;
      patterns[1013] = 25'b00000011_11110011_11110110_0;
      patterns[1014] = 25'b00000011_11110100_11110111_0;
      patterns[1015] = 25'b00000011_11110101_11111000_0;
      patterns[1016] = 25'b00000011_11110110_11111001_0;
      patterns[1017] = 25'b00000011_11110111_11111010_0;
      patterns[1018] = 25'b00000011_11111000_11111011_0;
      patterns[1019] = 25'b00000011_11111001_11111100_0;
      patterns[1020] = 25'b00000011_11111010_11111101_0;
      patterns[1021] = 25'b00000011_11111011_11111110_0;
      patterns[1022] = 25'b00000011_11111100_11111111_0;
      patterns[1023] = 25'b00000011_11111101_00000000_1;
      patterns[1024] = 25'b00000011_11111110_00000001_1;
      patterns[1025] = 25'b00000011_11111111_00000010_1;
      patterns[1026] = 25'b00000100_00000000_00000100_0;
      patterns[1027] = 25'b00000100_00000001_00000101_0;
      patterns[1028] = 25'b00000100_00000010_00000110_0;
      patterns[1029] = 25'b00000100_00000011_00000111_0;
      patterns[1030] = 25'b00000100_00000100_00001000_0;
      patterns[1031] = 25'b00000100_00000101_00001001_0;
      patterns[1032] = 25'b00000100_00000110_00001010_0;
      patterns[1033] = 25'b00000100_00000111_00001011_0;
      patterns[1034] = 25'b00000100_00001000_00001100_0;
      patterns[1035] = 25'b00000100_00001001_00001101_0;
      patterns[1036] = 25'b00000100_00001010_00001110_0;
      patterns[1037] = 25'b00000100_00001011_00001111_0;
      patterns[1038] = 25'b00000100_00001100_00010000_0;
      patterns[1039] = 25'b00000100_00001101_00010001_0;
      patterns[1040] = 25'b00000100_00001110_00010010_0;
      patterns[1041] = 25'b00000100_00001111_00010011_0;
      patterns[1042] = 25'b00000100_00010000_00010100_0;
      patterns[1043] = 25'b00000100_00010001_00010101_0;
      patterns[1044] = 25'b00000100_00010010_00010110_0;
      patterns[1045] = 25'b00000100_00010011_00010111_0;
      patterns[1046] = 25'b00000100_00010100_00011000_0;
      patterns[1047] = 25'b00000100_00010101_00011001_0;
      patterns[1048] = 25'b00000100_00010110_00011010_0;
      patterns[1049] = 25'b00000100_00010111_00011011_0;
      patterns[1050] = 25'b00000100_00011000_00011100_0;
      patterns[1051] = 25'b00000100_00011001_00011101_0;
      patterns[1052] = 25'b00000100_00011010_00011110_0;
      patterns[1053] = 25'b00000100_00011011_00011111_0;
      patterns[1054] = 25'b00000100_00011100_00100000_0;
      patterns[1055] = 25'b00000100_00011101_00100001_0;
      patterns[1056] = 25'b00000100_00011110_00100010_0;
      patterns[1057] = 25'b00000100_00011111_00100011_0;
      patterns[1058] = 25'b00000100_00100000_00100100_0;
      patterns[1059] = 25'b00000100_00100001_00100101_0;
      patterns[1060] = 25'b00000100_00100010_00100110_0;
      patterns[1061] = 25'b00000100_00100011_00100111_0;
      patterns[1062] = 25'b00000100_00100100_00101000_0;
      patterns[1063] = 25'b00000100_00100101_00101001_0;
      patterns[1064] = 25'b00000100_00100110_00101010_0;
      patterns[1065] = 25'b00000100_00100111_00101011_0;
      patterns[1066] = 25'b00000100_00101000_00101100_0;
      patterns[1067] = 25'b00000100_00101001_00101101_0;
      patterns[1068] = 25'b00000100_00101010_00101110_0;
      patterns[1069] = 25'b00000100_00101011_00101111_0;
      patterns[1070] = 25'b00000100_00101100_00110000_0;
      patterns[1071] = 25'b00000100_00101101_00110001_0;
      patterns[1072] = 25'b00000100_00101110_00110010_0;
      patterns[1073] = 25'b00000100_00101111_00110011_0;
      patterns[1074] = 25'b00000100_00110000_00110100_0;
      patterns[1075] = 25'b00000100_00110001_00110101_0;
      patterns[1076] = 25'b00000100_00110010_00110110_0;
      patterns[1077] = 25'b00000100_00110011_00110111_0;
      patterns[1078] = 25'b00000100_00110100_00111000_0;
      patterns[1079] = 25'b00000100_00110101_00111001_0;
      patterns[1080] = 25'b00000100_00110110_00111010_0;
      patterns[1081] = 25'b00000100_00110111_00111011_0;
      patterns[1082] = 25'b00000100_00111000_00111100_0;
      patterns[1083] = 25'b00000100_00111001_00111101_0;
      patterns[1084] = 25'b00000100_00111010_00111110_0;
      patterns[1085] = 25'b00000100_00111011_00111111_0;
      patterns[1086] = 25'b00000100_00111100_01000000_0;
      patterns[1087] = 25'b00000100_00111101_01000001_0;
      patterns[1088] = 25'b00000100_00111110_01000010_0;
      patterns[1089] = 25'b00000100_00111111_01000011_0;
      patterns[1090] = 25'b00000100_01000000_01000100_0;
      patterns[1091] = 25'b00000100_01000001_01000101_0;
      patterns[1092] = 25'b00000100_01000010_01000110_0;
      patterns[1093] = 25'b00000100_01000011_01000111_0;
      patterns[1094] = 25'b00000100_01000100_01001000_0;
      patterns[1095] = 25'b00000100_01000101_01001001_0;
      patterns[1096] = 25'b00000100_01000110_01001010_0;
      patterns[1097] = 25'b00000100_01000111_01001011_0;
      patterns[1098] = 25'b00000100_01001000_01001100_0;
      patterns[1099] = 25'b00000100_01001001_01001101_0;
      patterns[1100] = 25'b00000100_01001010_01001110_0;
      patterns[1101] = 25'b00000100_01001011_01001111_0;
      patterns[1102] = 25'b00000100_01001100_01010000_0;
      patterns[1103] = 25'b00000100_01001101_01010001_0;
      patterns[1104] = 25'b00000100_01001110_01010010_0;
      patterns[1105] = 25'b00000100_01001111_01010011_0;
      patterns[1106] = 25'b00000100_01010000_01010100_0;
      patterns[1107] = 25'b00000100_01010001_01010101_0;
      patterns[1108] = 25'b00000100_01010010_01010110_0;
      patterns[1109] = 25'b00000100_01010011_01010111_0;
      patterns[1110] = 25'b00000100_01010100_01011000_0;
      patterns[1111] = 25'b00000100_01010101_01011001_0;
      patterns[1112] = 25'b00000100_01010110_01011010_0;
      patterns[1113] = 25'b00000100_01010111_01011011_0;
      patterns[1114] = 25'b00000100_01011000_01011100_0;
      patterns[1115] = 25'b00000100_01011001_01011101_0;
      patterns[1116] = 25'b00000100_01011010_01011110_0;
      patterns[1117] = 25'b00000100_01011011_01011111_0;
      patterns[1118] = 25'b00000100_01011100_01100000_0;
      patterns[1119] = 25'b00000100_01011101_01100001_0;
      patterns[1120] = 25'b00000100_01011110_01100010_0;
      patterns[1121] = 25'b00000100_01011111_01100011_0;
      patterns[1122] = 25'b00000100_01100000_01100100_0;
      patterns[1123] = 25'b00000100_01100001_01100101_0;
      patterns[1124] = 25'b00000100_01100010_01100110_0;
      patterns[1125] = 25'b00000100_01100011_01100111_0;
      patterns[1126] = 25'b00000100_01100100_01101000_0;
      patterns[1127] = 25'b00000100_01100101_01101001_0;
      patterns[1128] = 25'b00000100_01100110_01101010_0;
      patterns[1129] = 25'b00000100_01100111_01101011_0;
      patterns[1130] = 25'b00000100_01101000_01101100_0;
      patterns[1131] = 25'b00000100_01101001_01101101_0;
      patterns[1132] = 25'b00000100_01101010_01101110_0;
      patterns[1133] = 25'b00000100_01101011_01101111_0;
      patterns[1134] = 25'b00000100_01101100_01110000_0;
      patterns[1135] = 25'b00000100_01101101_01110001_0;
      patterns[1136] = 25'b00000100_01101110_01110010_0;
      patterns[1137] = 25'b00000100_01101111_01110011_0;
      patterns[1138] = 25'b00000100_01110000_01110100_0;
      patterns[1139] = 25'b00000100_01110001_01110101_0;
      patterns[1140] = 25'b00000100_01110010_01110110_0;
      patterns[1141] = 25'b00000100_01110011_01110111_0;
      patterns[1142] = 25'b00000100_01110100_01111000_0;
      patterns[1143] = 25'b00000100_01110101_01111001_0;
      patterns[1144] = 25'b00000100_01110110_01111010_0;
      patterns[1145] = 25'b00000100_01110111_01111011_0;
      patterns[1146] = 25'b00000100_01111000_01111100_0;
      patterns[1147] = 25'b00000100_01111001_01111101_0;
      patterns[1148] = 25'b00000100_01111010_01111110_0;
      patterns[1149] = 25'b00000100_01111011_01111111_0;
      patterns[1150] = 25'b00000100_01111100_10000000_0;
      patterns[1151] = 25'b00000100_01111101_10000001_0;
      patterns[1152] = 25'b00000100_01111110_10000010_0;
      patterns[1153] = 25'b00000100_01111111_10000011_0;
      patterns[1154] = 25'b00000100_10000000_10000100_0;
      patterns[1155] = 25'b00000100_10000001_10000101_0;
      patterns[1156] = 25'b00000100_10000010_10000110_0;
      patterns[1157] = 25'b00000100_10000011_10000111_0;
      patterns[1158] = 25'b00000100_10000100_10001000_0;
      patterns[1159] = 25'b00000100_10000101_10001001_0;
      patterns[1160] = 25'b00000100_10000110_10001010_0;
      patterns[1161] = 25'b00000100_10000111_10001011_0;
      patterns[1162] = 25'b00000100_10001000_10001100_0;
      patterns[1163] = 25'b00000100_10001001_10001101_0;
      patterns[1164] = 25'b00000100_10001010_10001110_0;
      patterns[1165] = 25'b00000100_10001011_10001111_0;
      patterns[1166] = 25'b00000100_10001100_10010000_0;
      patterns[1167] = 25'b00000100_10001101_10010001_0;
      patterns[1168] = 25'b00000100_10001110_10010010_0;
      patterns[1169] = 25'b00000100_10001111_10010011_0;
      patterns[1170] = 25'b00000100_10010000_10010100_0;
      patterns[1171] = 25'b00000100_10010001_10010101_0;
      patterns[1172] = 25'b00000100_10010010_10010110_0;
      patterns[1173] = 25'b00000100_10010011_10010111_0;
      patterns[1174] = 25'b00000100_10010100_10011000_0;
      patterns[1175] = 25'b00000100_10010101_10011001_0;
      patterns[1176] = 25'b00000100_10010110_10011010_0;
      patterns[1177] = 25'b00000100_10010111_10011011_0;
      patterns[1178] = 25'b00000100_10011000_10011100_0;
      patterns[1179] = 25'b00000100_10011001_10011101_0;
      patterns[1180] = 25'b00000100_10011010_10011110_0;
      patterns[1181] = 25'b00000100_10011011_10011111_0;
      patterns[1182] = 25'b00000100_10011100_10100000_0;
      patterns[1183] = 25'b00000100_10011101_10100001_0;
      patterns[1184] = 25'b00000100_10011110_10100010_0;
      patterns[1185] = 25'b00000100_10011111_10100011_0;
      patterns[1186] = 25'b00000100_10100000_10100100_0;
      patterns[1187] = 25'b00000100_10100001_10100101_0;
      patterns[1188] = 25'b00000100_10100010_10100110_0;
      patterns[1189] = 25'b00000100_10100011_10100111_0;
      patterns[1190] = 25'b00000100_10100100_10101000_0;
      patterns[1191] = 25'b00000100_10100101_10101001_0;
      patterns[1192] = 25'b00000100_10100110_10101010_0;
      patterns[1193] = 25'b00000100_10100111_10101011_0;
      patterns[1194] = 25'b00000100_10101000_10101100_0;
      patterns[1195] = 25'b00000100_10101001_10101101_0;
      patterns[1196] = 25'b00000100_10101010_10101110_0;
      patterns[1197] = 25'b00000100_10101011_10101111_0;
      patterns[1198] = 25'b00000100_10101100_10110000_0;
      patterns[1199] = 25'b00000100_10101101_10110001_0;
      patterns[1200] = 25'b00000100_10101110_10110010_0;
      patterns[1201] = 25'b00000100_10101111_10110011_0;
      patterns[1202] = 25'b00000100_10110000_10110100_0;
      patterns[1203] = 25'b00000100_10110001_10110101_0;
      patterns[1204] = 25'b00000100_10110010_10110110_0;
      patterns[1205] = 25'b00000100_10110011_10110111_0;
      patterns[1206] = 25'b00000100_10110100_10111000_0;
      patterns[1207] = 25'b00000100_10110101_10111001_0;
      patterns[1208] = 25'b00000100_10110110_10111010_0;
      patterns[1209] = 25'b00000100_10110111_10111011_0;
      patterns[1210] = 25'b00000100_10111000_10111100_0;
      patterns[1211] = 25'b00000100_10111001_10111101_0;
      patterns[1212] = 25'b00000100_10111010_10111110_0;
      patterns[1213] = 25'b00000100_10111011_10111111_0;
      patterns[1214] = 25'b00000100_10111100_11000000_0;
      patterns[1215] = 25'b00000100_10111101_11000001_0;
      patterns[1216] = 25'b00000100_10111110_11000010_0;
      patterns[1217] = 25'b00000100_10111111_11000011_0;
      patterns[1218] = 25'b00000100_11000000_11000100_0;
      patterns[1219] = 25'b00000100_11000001_11000101_0;
      patterns[1220] = 25'b00000100_11000010_11000110_0;
      patterns[1221] = 25'b00000100_11000011_11000111_0;
      patterns[1222] = 25'b00000100_11000100_11001000_0;
      patterns[1223] = 25'b00000100_11000101_11001001_0;
      patterns[1224] = 25'b00000100_11000110_11001010_0;
      patterns[1225] = 25'b00000100_11000111_11001011_0;
      patterns[1226] = 25'b00000100_11001000_11001100_0;
      patterns[1227] = 25'b00000100_11001001_11001101_0;
      patterns[1228] = 25'b00000100_11001010_11001110_0;
      patterns[1229] = 25'b00000100_11001011_11001111_0;
      patterns[1230] = 25'b00000100_11001100_11010000_0;
      patterns[1231] = 25'b00000100_11001101_11010001_0;
      patterns[1232] = 25'b00000100_11001110_11010010_0;
      patterns[1233] = 25'b00000100_11001111_11010011_0;
      patterns[1234] = 25'b00000100_11010000_11010100_0;
      patterns[1235] = 25'b00000100_11010001_11010101_0;
      patterns[1236] = 25'b00000100_11010010_11010110_0;
      patterns[1237] = 25'b00000100_11010011_11010111_0;
      patterns[1238] = 25'b00000100_11010100_11011000_0;
      patterns[1239] = 25'b00000100_11010101_11011001_0;
      patterns[1240] = 25'b00000100_11010110_11011010_0;
      patterns[1241] = 25'b00000100_11010111_11011011_0;
      patterns[1242] = 25'b00000100_11011000_11011100_0;
      patterns[1243] = 25'b00000100_11011001_11011101_0;
      patterns[1244] = 25'b00000100_11011010_11011110_0;
      patterns[1245] = 25'b00000100_11011011_11011111_0;
      patterns[1246] = 25'b00000100_11011100_11100000_0;
      patterns[1247] = 25'b00000100_11011101_11100001_0;
      patterns[1248] = 25'b00000100_11011110_11100010_0;
      patterns[1249] = 25'b00000100_11011111_11100011_0;
      patterns[1250] = 25'b00000100_11100000_11100100_0;
      patterns[1251] = 25'b00000100_11100001_11100101_0;
      patterns[1252] = 25'b00000100_11100010_11100110_0;
      patterns[1253] = 25'b00000100_11100011_11100111_0;
      patterns[1254] = 25'b00000100_11100100_11101000_0;
      patterns[1255] = 25'b00000100_11100101_11101001_0;
      patterns[1256] = 25'b00000100_11100110_11101010_0;
      patterns[1257] = 25'b00000100_11100111_11101011_0;
      patterns[1258] = 25'b00000100_11101000_11101100_0;
      patterns[1259] = 25'b00000100_11101001_11101101_0;
      patterns[1260] = 25'b00000100_11101010_11101110_0;
      patterns[1261] = 25'b00000100_11101011_11101111_0;
      patterns[1262] = 25'b00000100_11101100_11110000_0;
      patterns[1263] = 25'b00000100_11101101_11110001_0;
      patterns[1264] = 25'b00000100_11101110_11110010_0;
      patterns[1265] = 25'b00000100_11101111_11110011_0;
      patterns[1266] = 25'b00000100_11110000_11110100_0;
      patterns[1267] = 25'b00000100_11110001_11110101_0;
      patterns[1268] = 25'b00000100_11110010_11110110_0;
      patterns[1269] = 25'b00000100_11110011_11110111_0;
      patterns[1270] = 25'b00000100_11110100_11111000_0;
      patterns[1271] = 25'b00000100_11110101_11111001_0;
      patterns[1272] = 25'b00000100_11110110_11111010_0;
      patterns[1273] = 25'b00000100_11110111_11111011_0;
      patterns[1274] = 25'b00000100_11111000_11111100_0;
      patterns[1275] = 25'b00000100_11111001_11111101_0;
      patterns[1276] = 25'b00000100_11111010_11111110_0;
      patterns[1277] = 25'b00000100_11111011_11111111_0;
      patterns[1278] = 25'b00000100_11111100_00000000_1;
      patterns[1279] = 25'b00000100_11111101_00000001_1;
      patterns[1280] = 25'b00000100_11111110_00000010_1;
      patterns[1281] = 25'b00000100_11111111_00000011_1;
      patterns[1282] = 25'b00000101_00000000_00000101_0;
      patterns[1283] = 25'b00000101_00000001_00000110_0;
      patterns[1284] = 25'b00000101_00000010_00000111_0;
      patterns[1285] = 25'b00000101_00000011_00001000_0;
      patterns[1286] = 25'b00000101_00000100_00001001_0;
      patterns[1287] = 25'b00000101_00000101_00001010_0;
      patterns[1288] = 25'b00000101_00000110_00001011_0;
      patterns[1289] = 25'b00000101_00000111_00001100_0;
      patterns[1290] = 25'b00000101_00001000_00001101_0;
      patterns[1291] = 25'b00000101_00001001_00001110_0;
      patterns[1292] = 25'b00000101_00001010_00001111_0;
      patterns[1293] = 25'b00000101_00001011_00010000_0;
      patterns[1294] = 25'b00000101_00001100_00010001_0;
      patterns[1295] = 25'b00000101_00001101_00010010_0;
      patterns[1296] = 25'b00000101_00001110_00010011_0;
      patterns[1297] = 25'b00000101_00001111_00010100_0;
      patterns[1298] = 25'b00000101_00010000_00010101_0;
      patterns[1299] = 25'b00000101_00010001_00010110_0;
      patterns[1300] = 25'b00000101_00010010_00010111_0;
      patterns[1301] = 25'b00000101_00010011_00011000_0;
      patterns[1302] = 25'b00000101_00010100_00011001_0;
      patterns[1303] = 25'b00000101_00010101_00011010_0;
      patterns[1304] = 25'b00000101_00010110_00011011_0;
      patterns[1305] = 25'b00000101_00010111_00011100_0;
      patterns[1306] = 25'b00000101_00011000_00011101_0;
      patterns[1307] = 25'b00000101_00011001_00011110_0;
      patterns[1308] = 25'b00000101_00011010_00011111_0;
      patterns[1309] = 25'b00000101_00011011_00100000_0;
      patterns[1310] = 25'b00000101_00011100_00100001_0;
      patterns[1311] = 25'b00000101_00011101_00100010_0;
      patterns[1312] = 25'b00000101_00011110_00100011_0;
      patterns[1313] = 25'b00000101_00011111_00100100_0;
      patterns[1314] = 25'b00000101_00100000_00100101_0;
      patterns[1315] = 25'b00000101_00100001_00100110_0;
      patterns[1316] = 25'b00000101_00100010_00100111_0;
      patterns[1317] = 25'b00000101_00100011_00101000_0;
      patterns[1318] = 25'b00000101_00100100_00101001_0;
      patterns[1319] = 25'b00000101_00100101_00101010_0;
      patterns[1320] = 25'b00000101_00100110_00101011_0;
      patterns[1321] = 25'b00000101_00100111_00101100_0;
      patterns[1322] = 25'b00000101_00101000_00101101_0;
      patterns[1323] = 25'b00000101_00101001_00101110_0;
      patterns[1324] = 25'b00000101_00101010_00101111_0;
      patterns[1325] = 25'b00000101_00101011_00110000_0;
      patterns[1326] = 25'b00000101_00101100_00110001_0;
      patterns[1327] = 25'b00000101_00101101_00110010_0;
      patterns[1328] = 25'b00000101_00101110_00110011_0;
      patterns[1329] = 25'b00000101_00101111_00110100_0;
      patterns[1330] = 25'b00000101_00110000_00110101_0;
      patterns[1331] = 25'b00000101_00110001_00110110_0;
      patterns[1332] = 25'b00000101_00110010_00110111_0;
      patterns[1333] = 25'b00000101_00110011_00111000_0;
      patterns[1334] = 25'b00000101_00110100_00111001_0;
      patterns[1335] = 25'b00000101_00110101_00111010_0;
      patterns[1336] = 25'b00000101_00110110_00111011_0;
      patterns[1337] = 25'b00000101_00110111_00111100_0;
      patterns[1338] = 25'b00000101_00111000_00111101_0;
      patterns[1339] = 25'b00000101_00111001_00111110_0;
      patterns[1340] = 25'b00000101_00111010_00111111_0;
      patterns[1341] = 25'b00000101_00111011_01000000_0;
      patterns[1342] = 25'b00000101_00111100_01000001_0;
      patterns[1343] = 25'b00000101_00111101_01000010_0;
      patterns[1344] = 25'b00000101_00111110_01000011_0;
      patterns[1345] = 25'b00000101_00111111_01000100_0;
      patterns[1346] = 25'b00000101_01000000_01000101_0;
      patterns[1347] = 25'b00000101_01000001_01000110_0;
      patterns[1348] = 25'b00000101_01000010_01000111_0;
      patterns[1349] = 25'b00000101_01000011_01001000_0;
      patterns[1350] = 25'b00000101_01000100_01001001_0;
      patterns[1351] = 25'b00000101_01000101_01001010_0;
      patterns[1352] = 25'b00000101_01000110_01001011_0;
      patterns[1353] = 25'b00000101_01000111_01001100_0;
      patterns[1354] = 25'b00000101_01001000_01001101_0;
      patterns[1355] = 25'b00000101_01001001_01001110_0;
      patterns[1356] = 25'b00000101_01001010_01001111_0;
      patterns[1357] = 25'b00000101_01001011_01010000_0;
      patterns[1358] = 25'b00000101_01001100_01010001_0;
      patterns[1359] = 25'b00000101_01001101_01010010_0;
      patterns[1360] = 25'b00000101_01001110_01010011_0;
      patterns[1361] = 25'b00000101_01001111_01010100_0;
      patterns[1362] = 25'b00000101_01010000_01010101_0;
      patterns[1363] = 25'b00000101_01010001_01010110_0;
      patterns[1364] = 25'b00000101_01010010_01010111_0;
      patterns[1365] = 25'b00000101_01010011_01011000_0;
      patterns[1366] = 25'b00000101_01010100_01011001_0;
      patterns[1367] = 25'b00000101_01010101_01011010_0;
      patterns[1368] = 25'b00000101_01010110_01011011_0;
      patterns[1369] = 25'b00000101_01010111_01011100_0;
      patterns[1370] = 25'b00000101_01011000_01011101_0;
      patterns[1371] = 25'b00000101_01011001_01011110_0;
      patterns[1372] = 25'b00000101_01011010_01011111_0;
      patterns[1373] = 25'b00000101_01011011_01100000_0;
      patterns[1374] = 25'b00000101_01011100_01100001_0;
      patterns[1375] = 25'b00000101_01011101_01100010_0;
      patterns[1376] = 25'b00000101_01011110_01100011_0;
      patterns[1377] = 25'b00000101_01011111_01100100_0;
      patterns[1378] = 25'b00000101_01100000_01100101_0;
      patterns[1379] = 25'b00000101_01100001_01100110_0;
      patterns[1380] = 25'b00000101_01100010_01100111_0;
      patterns[1381] = 25'b00000101_01100011_01101000_0;
      patterns[1382] = 25'b00000101_01100100_01101001_0;
      patterns[1383] = 25'b00000101_01100101_01101010_0;
      patterns[1384] = 25'b00000101_01100110_01101011_0;
      patterns[1385] = 25'b00000101_01100111_01101100_0;
      patterns[1386] = 25'b00000101_01101000_01101101_0;
      patterns[1387] = 25'b00000101_01101001_01101110_0;
      patterns[1388] = 25'b00000101_01101010_01101111_0;
      patterns[1389] = 25'b00000101_01101011_01110000_0;
      patterns[1390] = 25'b00000101_01101100_01110001_0;
      patterns[1391] = 25'b00000101_01101101_01110010_0;
      patterns[1392] = 25'b00000101_01101110_01110011_0;
      patterns[1393] = 25'b00000101_01101111_01110100_0;
      patterns[1394] = 25'b00000101_01110000_01110101_0;
      patterns[1395] = 25'b00000101_01110001_01110110_0;
      patterns[1396] = 25'b00000101_01110010_01110111_0;
      patterns[1397] = 25'b00000101_01110011_01111000_0;
      patterns[1398] = 25'b00000101_01110100_01111001_0;
      patterns[1399] = 25'b00000101_01110101_01111010_0;
      patterns[1400] = 25'b00000101_01110110_01111011_0;
      patterns[1401] = 25'b00000101_01110111_01111100_0;
      patterns[1402] = 25'b00000101_01111000_01111101_0;
      patterns[1403] = 25'b00000101_01111001_01111110_0;
      patterns[1404] = 25'b00000101_01111010_01111111_0;
      patterns[1405] = 25'b00000101_01111011_10000000_0;
      patterns[1406] = 25'b00000101_01111100_10000001_0;
      patterns[1407] = 25'b00000101_01111101_10000010_0;
      patterns[1408] = 25'b00000101_01111110_10000011_0;
      patterns[1409] = 25'b00000101_01111111_10000100_0;
      patterns[1410] = 25'b00000101_10000000_10000101_0;
      patterns[1411] = 25'b00000101_10000001_10000110_0;
      patterns[1412] = 25'b00000101_10000010_10000111_0;
      patterns[1413] = 25'b00000101_10000011_10001000_0;
      patterns[1414] = 25'b00000101_10000100_10001001_0;
      patterns[1415] = 25'b00000101_10000101_10001010_0;
      patterns[1416] = 25'b00000101_10000110_10001011_0;
      patterns[1417] = 25'b00000101_10000111_10001100_0;
      patterns[1418] = 25'b00000101_10001000_10001101_0;
      patterns[1419] = 25'b00000101_10001001_10001110_0;
      patterns[1420] = 25'b00000101_10001010_10001111_0;
      patterns[1421] = 25'b00000101_10001011_10010000_0;
      patterns[1422] = 25'b00000101_10001100_10010001_0;
      patterns[1423] = 25'b00000101_10001101_10010010_0;
      patterns[1424] = 25'b00000101_10001110_10010011_0;
      patterns[1425] = 25'b00000101_10001111_10010100_0;
      patterns[1426] = 25'b00000101_10010000_10010101_0;
      patterns[1427] = 25'b00000101_10010001_10010110_0;
      patterns[1428] = 25'b00000101_10010010_10010111_0;
      patterns[1429] = 25'b00000101_10010011_10011000_0;
      patterns[1430] = 25'b00000101_10010100_10011001_0;
      patterns[1431] = 25'b00000101_10010101_10011010_0;
      patterns[1432] = 25'b00000101_10010110_10011011_0;
      patterns[1433] = 25'b00000101_10010111_10011100_0;
      patterns[1434] = 25'b00000101_10011000_10011101_0;
      patterns[1435] = 25'b00000101_10011001_10011110_0;
      patterns[1436] = 25'b00000101_10011010_10011111_0;
      patterns[1437] = 25'b00000101_10011011_10100000_0;
      patterns[1438] = 25'b00000101_10011100_10100001_0;
      patterns[1439] = 25'b00000101_10011101_10100010_0;
      patterns[1440] = 25'b00000101_10011110_10100011_0;
      patterns[1441] = 25'b00000101_10011111_10100100_0;
      patterns[1442] = 25'b00000101_10100000_10100101_0;
      patterns[1443] = 25'b00000101_10100001_10100110_0;
      patterns[1444] = 25'b00000101_10100010_10100111_0;
      patterns[1445] = 25'b00000101_10100011_10101000_0;
      patterns[1446] = 25'b00000101_10100100_10101001_0;
      patterns[1447] = 25'b00000101_10100101_10101010_0;
      patterns[1448] = 25'b00000101_10100110_10101011_0;
      patterns[1449] = 25'b00000101_10100111_10101100_0;
      patterns[1450] = 25'b00000101_10101000_10101101_0;
      patterns[1451] = 25'b00000101_10101001_10101110_0;
      patterns[1452] = 25'b00000101_10101010_10101111_0;
      patterns[1453] = 25'b00000101_10101011_10110000_0;
      patterns[1454] = 25'b00000101_10101100_10110001_0;
      patterns[1455] = 25'b00000101_10101101_10110010_0;
      patterns[1456] = 25'b00000101_10101110_10110011_0;
      patterns[1457] = 25'b00000101_10101111_10110100_0;
      patterns[1458] = 25'b00000101_10110000_10110101_0;
      patterns[1459] = 25'b00000101_10110001_10110110_0;
      patterns[1460] = 25'b00000101_10110010_10110111_0;
      patterns[1461] = 25'b00000101_10110011_10111000_0;
      patterns[1462] = 25'b00000101_10110100_10111001_0;
      patterns[1463] = 25'b00000101_10110101_10111010_0;
      patterns[1464] = 25'b00000101_10110110_10111011_0;
      patterns[1465] = 25'b00000101_10110111_10111100_0;
      patterns[1466] = 25'b00000101_10111000_10111101_0;
      patterns[1467] = 25'b00000101_10111001_10111110_0;
      patterns[1468] = 25'b00000101_10111010_10111111_0;
      patterns[1469] = 25'b00000101_10111011_11000000_0;
      patterns[1470] = 25'b00000101_10111100_11000001_0;
      patterns[1471] = 25'b00000101_10111101_11000010_0;
      patterns[1472] = 25'b00000101_10111110_11000011_0;
      patterns[1473] = 25'b00000101_10111111_11000100_0;
      patterns[1474] = 25'b00000101_11000000_11000101_0;
      patterns[1475] = 25'b00000101_11000001_11000110_0;
      patterns[1476] = 25'b00000101_11000010_11000111_0;
      patterns[1477] = 25'b00000101_11000011_11001000_0;
      patterns[1478] = 25'b00000101_11000100_11001001_0;
      patterns[1479] = 25'b00000101_11000101_11001010_0;
      patterns[1480] = 25'b00000101_11000110_11001011_0;
      patterns[1481] = 25'b00000101_11000111_11001100_0;
      patterns[1482] = 25'b00000101_11001000_11001101_0;
      patterns[1483] = 25'b00000101_11001001_11001110_0;
      patterns[1484] = 25'b00000101_11001010_11001111_0;
      patterns[1485] = 25'b00000101_11001011_11010000_0;
      patterns[1486] = 25'b00000101_11001100_11010001_0;
      patterns[1487] = 25'b00000101_11001101_11010010_0;
      patterns[1488] = 25'b00000101_11001110_11010011_0;
      patterns[1489] = 25'b00000101_11001111_11010100_0;
      patterns[1490] = 25'b00000101_11010000_11010101_0;
      patterns[1491] = 25'b00000101_11010001_11010110_0;
      patterns[1492] = 25'b00000101_11010010_11010111_0;
      patterns[1493] = 25'b00000101_11010011_11011000_0;
      patterns[1494] = 25'b00000101_11010100_11011001_0;
      patterns[1495] = 25'b00000101_11010101_11011010_0;
      patterns[1496] = 25'b00000101_11010110_11011011_0;
      patterns[1497] = 25'b00000101_11010111_11011100_0;
      patterns[1498] = 25'b00000101_11011000_11011101_0;
      patterns[1499] = 25'b00000101_11011001_11011110_0;
      patterns[1500] = 25'b00000101_11011010_11011111_0;
      patterns[1501] = 25'b00000101_11011011_11100000_0;
      patterns[1502] = 25'b00000101_11011100_11100001_0;
      patterns[1503] = 25'b00000101_11011101_11100010_0;
      patterns[1504] = 25'b00000101_11011110_11100011_0;
      patterns[1505] = 25'b00000101_11011111_11100100_0;
      patterns[1506] = 25'b00000101_11100000_11100101_0;
      patterns[1507] = 25'b00000101_11100001_11100110_0;
      patterns[1508] = 25'b00000101_11100010_11100111_0;
      patterns[1509] = 25'b00000101_11100011_11101000_0;
      patterns[1510] = 25'b00000101_11100100_11101001_0;
      patterns[1511] = 25'b00000101_11100101_11101010_0;
      patterns[1512] = 25'b00000101_11100110_11101011_0;
      patterns[1513] = 25'b00000101_11100111_11101100_0;
      patterns[1514] = 25'b00000101_11101000_11101101_0;
      patterns[1515] = 25'b00000101_11101001_11101110_0;
      patterns[1516] = 25'b00000101_11101010_11101111_0;
      patterns[1517] = 25'b00000101_11101011_11110000_0;
      patterns[1518] = 25'b00000101_11101100_11110001_0;
      patterns[1519] = 25'b00000101_11101101_11110010_0;
      patterns[1520] = 25'b00000101_11101110_11110011_0;
      patterns[1521] = 25'b00000101_11101111_11110100_0;
      patterns[1522] = 25'b00000101_11110000_11110101_0;
      patterns[1523] = 25'b00000101_11110001_11110110_0;
      patterns[1524] = 25'b00000101_11110010_11110111_0;
      patterns[1525] = 25'b00000101_11110011_11111000_0;
      patterns[1526] = 25'b00000101_11110100_11111001_0;
      patterns[1527] = 25'b00000101_11110101_11111010_0;
      patterns[1528] = 25'b00000101_11110110_11111011_0;
      patterns[1529] = 25'b00000101_11110111_11111100_0;
      patterns[1530] = 25'b00000101_11111000_11111101_0;
      patterns[1531] = 25'b00000101_11111001_11111110_0;
      patterns[1532] = 25'b00000101_11111010_11111111_0;
      patterns[1533] = 25'b00000101_11111011_00000000_1;
      patterns[1534] = 25'b00000101_11111100_00000001_1;
      patterns[1535] = 25'b00000101_11111101_00000010_1;
      patterns[1536] = 25'b00000101_11111110_00000011_1;
      patterns[1537] = 25'b00000101_11111111_00000100_1;
      patterns[1538] = 25'b00000110_00000000_00000110_0;
      patterns[1539] = 25'b00000110_00000001_00000111_0;
      patterns[1540] = 25'b00000110_00000010_00001000_0;
      patterns[1541] = 25'b00000110_00000011_00001001_0;
      patterns[1542] = 25'b00000110_00000100_00001010_0;
      patterns[1543] = 25'b00000110_00000101_00001011_0;
      patterns[1544] = 25'b00000110_00000110_00001100_0;
      patterns[1545] = 25'b00000110_00000111_00001101_0;
      patterns[1546] = 25'b00000110_00001000_00001110_0;
      patterns[1547] = 25'b00000110_00001001_00001111_0;
      patterns[1548] = 25'b00000110_00001010_00010000_0;
      patterns[1549] = 25'b00000110_00001011_00010001_0;
      patterns[1550] = 25'b00000110_00001100_00010010_0;
      patterns[1551] = 25'b00000110_00001101_00010011_0;
      patterns[1552] = 25'b00000110_00001110_00010100_0;
      patterns[1553] = 25'b00000110_00001111_00010101_0;
      patterns[1554] = 25'b00000110_00010000_00010110_0;
      patterns[1555] = 25'b00000110_00010001_00010111_0;
      patterns[1556] = 25'b00000110_00010010_00011000_0;
      patterns[1557] = 25'b00000110_00010011_00011001_0;
      patterns[1558] = 25'b00000110_00010100_00011010_0;
      patterns[1559] = 25'b00000110_00010101_00011011_0;
      patterns[1560] = 25'b00000110_00010110_00011100_0;
      patterns[1561] = 25'b00000110_00010111_00011101_0;
      patterns[1562] = 25'b00000110_00011000_00011110_0;
      patterns[1563] = 25'b00000110_00011001_00011111_0;
      patterns[1564] = 25'b00000110_00011010_00100000_0;
      patterns[1565] = 25'b00000110_00011011_00100001_0;
      patterns[1566] = 25'b00000110_00011100_00100010_0;
      patterns[1567] = 25'b00000110_00011101_00100011_0;
      patterns[1568] = 25'b00000110_00011110_00100100_0;
      patterns[1569] = 25'b00000110_00011111_00100101_0;
      patterns[1570] = 25'b00000110_00100000_00100110_0;
      patterns[1571] = 25'b00000110_00100001_00100111_0;
      patterns[1572] = 25'b00000110_00100010_00101000_0;
      patterns[1573] = 25'b00000110_00100011_00101001_0;
      patterns[1574] = 25'b00000110_00100100_00101010_0;
      patterns[1575] = 25'b00000110_00100101_00101011_0;
      patterns[1576] = 25'b00000110_00100110_00101100_0;
      patterns[1577] = 25'b00000110_00100111_00101101_0;
      patterns[1578] = 25'b00000110_00101000_00101110_0;
      patterns[1579] = 25'b00000110_00101001_00101111_0;
      patterns[1580] = 25'b00000110_00101010_00110000_0;
      patterns[1581] = 25'b00000110_00101011_00110001_0;
      patterns[1582] = 25'b00000110_00101100_00110010_0;
      patterns[1583] = 25'b00000110_00101101_00110011_0;
      patterns[1584] = 25'b00000110_00101110_00110100_0;
      patterns[1585] = 25'b00000110_00101111_00110101_0;
      patterns[1586] = 25'b00000110_00110000_00110110_0;
      patterns[1587] = 25'b00000110_00110001_00110111_0;
      patterns[1588] = 25'b00000110_00110010_00111000_0;
      patterns[1589] = 25'b00000110_00110011_00111001_0;
      patterns[1590] = 25'b00000110_00110100_00111010_0;
      patterns[1591] = 25'b00000110_00110101_00111011_0;
      patterns[1592] = 25'b00000110_00110110_00111100_0;
      patterns[1593] = 25'b00000110_00110111_00111101_0;
      patterns[1594] = 25'b00000110_00111000_00111110_0;
      patterns[1595] = 25'b00000110_00111001_00111111_0;
      patterns[1596] = 25'b00000110_00111010_01000000_0;
      patterns[1597] = 25'b00000110_00111011_01000001_0;
      patterns[1598] = 25'b00000110_00111100_01000010_0;
      patterns[1599] = 25'b00000110_00111101_01000011_0;
      patterns[1600] = 25'b00000110_00111110_01000100_0;
      patterns[1601] = 25'b00000110_00111111_01000101_0;
      patterns[1602] = 25'b00000110_01000000_01000110_0;
      patterns[1603] = 25'b00000110_01000001_01000111_0;
      patterns[1604] = 25'b00000110_01000010_01001000_0;
      patterns[1605] = 25'b00000110_01000011_01001001_0;
      patterns[1606] = 25'b00000110_01000100_01001010_0;
      patterns[1607] = 25'b00000110_01000101_01001011_0;
      patterns[1608] = 25'b00000110_01000110_01001100_0;
      patterns[1609] = 25'b00000110_01000111_01001101_0;
      patterns[1610] = 25'b00000110_01001000_01001110_0;
      patterns[1611] = 25'b00000110_01001001_01001111_0;
      patterns[1612] = 25'b00000110_01001010_01010000_0;
      patterns[1613] = 25'b00000110_01001011_01010001_0;
      patterns[1614] = 25'b00000110_01001100_01010010_0;
      patterns[1615] = 25'b00000110_01001101_01010011_0;
      patterns[1616] = 25'b00000110_01001110_01010100_0;
      patterns[1617] = 25'b00000110_01001111_01010101_0;
      patterns[1618] = 25'b00000110_01010000_01010110_0;
      patterns[1619] = 25'b00000110_01010001_01010111_0;
      patterns[1620] = 25'b00000110_01010010_01011000_0;
      patterns[1621] = 25'b00000110_01010011_01011001_0;
      patterns[1622] = 25'b00000110_01010100_01011010_0;
      patterns[1623] = 25'b00000110_01010101_01011011_0;
      patterns[1624] = 25'b00000110_01010110_01011100_0;
      patterns[1625] = 25'b00000110_01010111_01011101_0;
      patterns[1626] = 25'b00000110_01011000_01011110_0;
      patterns[1627] = 25'b00000110_01011001_01011111_0;
      patterns[1628] = 25'b00000110_01011010_01100000_0;
      patterns[1629] = 25'b00000110_01011011_01100001_0;
      patterns[1630] = 25'b00000110_01011100_01100010_0;
      patterns[1631] = 25'b00000110_01011101_01100011_0;
      patterns[1632] = 25'b00000110_01011110_01100100_0;
      patterns[1633] = 25'b00000110_01011111_01100101_0;
      patterns[1634] = 25'b00000110_01100000_01100110_0;
      patterns[1635] = 25'b00000110_01100001_01100111_0;
      patterns[1636] = 25'b00000110_01100010_01101000_0;
      patterns[1637] = 25'b00000110_01100011_01101001_0;
      patterns[1638] = 25'b00000110_01100100_01101010_0;
      patterns[1639] = 25'b00000110_01100101_01101011_0;
      patterns[1640] = 25'b00000110_01100110_01101100_0;
      patterns[1641] = 25'b00000110_01100111_01101101_0;
      patterns[1642] = 25'b00000110_01101000_01101110_0;
      patterns[1643] = 25'b00000110_01101001_01101111_0;
      patterns[1644] = 25'b00000110_01101010_01110000_0;
      patterns[1645] = 25'b00000110_01101011_01110001_0;
      patterns[1646] = 25'b00000110_01101100_01110010_0;
      patterns[1647] = 25'b00000110_01101101_01110011_0;
      patterns[1648] = 25'b00000110_01101110_01110100_0;
      patterns[1649] = 25'b00000110_01101111_01110101_0;
      patterns[1650] = 25'b00000110_01110000_01110110_0;
      patterns[1651] = 25'b00000110_01110001_01110111_0;
      patterns[1652] = 25'b00000110_01110010_01111000_0;
      patterns[1653] = 25'b00000110_01110011_01111001_0;
      patterns[1654] = 25'b00000110_01110100_01111010_0;
      patterns[1655] = 25'b00000110_01110101_01111011_0;
      patterns[1656] = 25'b00000110_01110110_01111100_0;
      patterns[1657] = 25'b00000110_01110111_01111101_0;
      patterns[1658] = 25'b00000110_01111000_01111110_0;
      patterns[1659] = 25'b00000110_01111001_01111111_0;
      patterns[1660] = 25'b00000110_01111010_10000000_0;
      patterns[1661] = 25'b00000110_01111011_10000001_0;
      patterns[1662] = 25'b00000110_01111100_10000010_0;
      patterns[1663] = 25'b00000110_01111101_10000011_0;
      patterns[1664] = 25'b00000110_01111110_10000100_0;
      patterns[1665] = 25'b00000110_01111111_10000101_0;
      patterns[1666] = 25'b00000110_10000000_10000110_0;
      patterns[1667] = 25'b00000110_10000001_10000111_0;
      patterns[1668] = 25'b00000110_10000010_10001000_0;
      patterns[1669] = 25'b00000110_10000011_10001001_0;
      patterns[1670] = 25'b00000110_10000100_10001010_0;
      patterns[1671] = 25'b00000110_10000101_10001011_0;
      patterns[1672] = 25'b00000110_10000110_10001100_0;
      patterns[1673] = 25'b00000110_10000111_10001101_0;
      patterns[1674] = 25'b00000110_10001000_10001110_0;
      patterns[1675] = 25'b00000110_10001001_10001111_0;
      patterns[1676] = 25'b00000110_10001010_10010000_0;
      patterns[1677] = 25'b00000110_10001011_10010001_0;
      patterns[1678] = 25'b00000110_10001100_10010010_0;
      patterns[1679] = 25'b00000110_10001101_10010011_0;
      patterns[1680] = 25'b00000110_10001110_10010100_0;
      patterns[1681] = 25'b00000110_10001111_10010101_0;
      patterns[1682] = 25'b00000110_10010000_10010110_0;
      patterns[1683] = 25'b00000110_10010001_10010111_0;
      patterns[1684] = 25'b00000110_10010010_10011000_0;
      patterns[1685] = 25'b00000110_10010011_10011001_0;
      patterns[1686] = 25'b00000110_10010100_10011010_0;
      patterns[1687] = 25'b00000110_10010101_10011011_0;
      patterns[1688] = 25'b00000110_10010110_10011100_0;
      patterns[1689] = 25'b00000110_10010111_10011101_0;
      patterns[1690] = 25'b00000110_10011000_10011110_0;
      patterns[1691] = 25'b00000110_10011001_10011111_0;
      patterns[1692] = 25'b00000110_10011010_10100000_0;
      patterns[1693] = 25'b00000110_10011011_10100001_0;
      patterns[1694] = 25'b00000110_10011100_10100010_0;
      patterns[1695] = 25'b00000110_10011101_10100011_0;
      patterns[1696] = 25'b00000110_10011110_10100100_0;
      patterns[1697] = 25'b00000110_10011111_10100101_0;
      patterns[1698] = 25'b00000110_10100000_10100110_0;
      patterns[1699] = 25'b00000110_10100001_10100111_0;
      patterns[1700] = 25'b00000110_10100010_10101000_0;
      patterns[1701] = 25'b00000110_10100011_10101001_0;
      patterns[1702] = 25'b00000110_10100100_10101010_0;
      patterns[1703] = 25'b00000110_10100101_10101011_0;
      patterns[1704] = 25'b00000110_10100110_10101100_0;
      patterns[1705] = 25'b00000110_10100111_10101101_0;
      patterns[1706] = 25'b00000110_10101000_10101110_0;
      patterns[1707] = 25'b00000110_10101001_10101111_0;
      patterns[1708] = 25'b00000110_10101010_10110000_0;
      patterns[1709] = 25'b00000110_10101011_10110001_0;
      patterns[1710] = 25'b00000110_10101100_10110010_0;
      patterns[1711] = 25'b00000110_10101101_10110011_0;
      patterns[1712] = 25'b00000110_10101110_10110100_0;
      patterns[1713] = 25'b00000110_10101111_10110101_0;
      patterns[1714] = 25'b00000110_10110000_10110110_0;
      patterns[1715] = 25'b00000110_10110001_10110111_0;
      patterns[1716] = 25'b00000110_10110010_10111000_0;
      patterns[1717] = 25'b00000110_10110011_10111001_0;
      patterns[1718] = 25'b00000110_10110100_10111010_0;
      patterns[1719] = 25'b00000110_10110101_10111011_0;
      patterns[1720] = 25'b00000110_10110110_10111100_0;
      patterns[1721] = 25'b00000110_10110111_10111101_0;
      patterns[1722] = 25'b00000110_10111000_10111110_0;
      patterns[1723] = 25'b00000110_10111001_10111111_0;
      patterns[1724] = 25'b00000110_10111010_11000000_0;
      patterns[1725] = 25'b00000110_10111011_11000001_0;
      patterns[1726] = 25'b00000110_10111100_11000010_0;
      patterns[1727] = 25'b00000110_10111101_11000011_0;
      patterns[1728] = 25'b00000110_10111110_11000100_0;
      patterns[1729] = 25'b00000110_10111111_11000101_0;
      patterns[1730] = 25'b00000110_11000000_11000110_0;
      patterns[1731] = 25'b00000110_11000001_11000111_0;
      patterns[1732] = 25'b00000110_11000010_11001000_0;
      patterns[1733] = 25'b00000110_11000011_11001001_0;
      patterns[1734] = 25'b00000110_11000100_11001010_0;
      patterns[1735] = 25'b00000110_11000101_11001011_0;
      patterns[1736] = 25'b00000110_11000110_11001100_0;
      patterns[1737] = 25'b00000110_11000111_11001101_0;
      patterns[1738] = 25'b00000110_11001000_11001110_0;
      patterns[1739] = 25'b00000110_11001001_11001111_0;
      patterns[1740] = 25'b00000110_11001010_11010000_0;
      patterns[1741] = 25'b00000110_11001011_11010001_0;
      patterns[1742] = 25'b00000110_11001100_11010010_0;
      patterns[1743] = 25'b00000110_11001101_11010011_0;
      patterns[1744] = 25'b00000110_11001110_11010100_0;
      patterns[1745] = 25'b00000110_11001111_11010101_0;
      patterns[1746] = 25'b00000110_11010000_11010110_0;
      patterns[1747] = 25'b00000110_11010001_11010111_0;
      patterns[1748] = 25'b00000110_11010010_11011000_0;
      patterns[1749] = 25'b00000110_11010011_11011001_0;
      patterns[1750] = 25'b00000110_11010100_11011010_0;
      patterns[1751] = 25'b00000110_11010101_11011011_0;
      patterns[1752] = 25'b00000110_11010110_11011100_0;
      patterns[1753] = 25'b00000110_11010111_11011101_0;
      patterns[1754] = 25'b00000110_11011000_11011110_0;
      patterns[1755] = 25'b00000110_11011001_11011111_0;
      patterns[1756] = 25'b00000110_11011010_11100000_0;
      patterns[1757] = 25'b00000110_11011011_11100001_0;
      patterns[1758] = 25'b00000110_11011100_11100010_0;
      patterns[1759] = 25'b00000110_11011101_11100011_0;
      patterns[1760] = 25'b00000110_11011110_11100100_0;
      patterns[1761] = 25'b00000110_11011111_11100101_0;
      patterns[1762] = 25'b00000110_11100000_11100110_0;
      patterns[1763] = 25'b00000110_11100001_11100111_0;
      patterns[1764] = 25'b00000110_11100010_11101000_0;
      patterns[1765] = 25'b00000110_11100011_11101001_0;
      patterns[1766] = 25'b00000110_11100100_11101010_0;
      patterns[1767] = 25'b00000110_11100101_11101011_0;
      patterns[1768] = 25'b00000110_11100110_11101100_0;
      patterns[1769] = 25'b00000110_11100111_11101101_0;
      patterns[1770] = 25'b00000110_11101000_11101110_0;
      patterns[1771] = 25'b00000110_11101001_11101111_0;
      patterns[1772] = 25'b00000110_11101010_11110000_0;
      patterns[1773] = 25'b00000110_11101011_11110001_0;
      patterns[1774] = 25'b00000110_11101100_11110010_0;
      patterns[1775] = 25'b00000110_11101101_11110011_0;
      patterns[1776] = 25'b00000110_11101110_11110100_0;
      patterns[1777] = 25'b00000110_11101111_11110101_0;
      patterns[1778] = 25'b00000110_11110000_11110110_0;
      patterns[1779] = 25'b00000110_11110001_11110111_0;
      patterns[1780] = 25'b00000110_11110010_11111000_0;
      patterns[1781] = 25'b00000110_11110011_11111001_0;
      patterns[1782] = 25'b00000110_11110100_11111010_0;
      patterns[1783] = 25'b00000110_11110101_11111011_0;
      patterns[1784] = 25'b00000110_11110110_11111100_0;
      patterns[1785] = 25'b00000110_11110111_11111101_0;
      patterns[1786] = 25'b00000110_11111000_11111110_0;
      patterns[1787] = 25'b00000110_11111001_11111111_0;
      patterns[1788] = 25'b00000110_11111010_00000000_1;
      patterns[1789] = 25'b00000110_11111011_00000001_1;
      patterns[1790] = 25'b00000110_11111100_00000010_1;
      patterns[1791] = 25'b00000110_11111101_00000011_1;
      patterns[1792] = 25'b00000110_11111110_00000100_1;
      patterns[1793] = 25'b00000110_11111111_00000101_1;
      patterns[1794] = 25'b00000111_00000000_00000111_0;
      patterns[1795] = 25'b00000111_00000001_00001000_0;
      patterns[1796] = 25'b00000111_00000010_00001001_0;
      patterns[1797] = 25'b00000111_00000011_00001010_0;
      patterns[1798] = 25'b00000111_00000100_00001011_0;
      patterns[1799] = 25'b00000111_00000101_00001100_0;
      patterns[1800] = 25'b00000111_00000110_00001101_0;
      patterns[1801] = 25'b00000111_00000111_00001110_0;
      patterns[1802] = 25'b00000111_00001000_00001111_0;
      patterns[1803] = 25'b00000111_00001001_00010000_0;
      patterns[1804] = 25'b00000111_00001010_00010001_0;
      patterns[1805] = 25'b00000111_00001011_00010010_0;
      patterns[1806] = 25'b00000111_00001100_00010011_0;
      patterns[1807] = 25'b00000111_00001101_00010100_0;
      patterns[1808] = 25'b00000111_00001110_00010101_0;
      patterns[1809] = 25'b00000111_00001111_00010110_0;
      patterns[1810] = 25'b00000111_00010000_00010111_0;
      patterns[1811] = 25'b00000111_00010001_00011000_0;
      patterns[1812] = 25'b00000111_00010010_00011001_0;
      patterns[1813] = 25'b00000111_00010011_00011010_0;
      patterns[1814] = 25'b00000111_00010100_00011011_0;
      patterns[1815] = 25'b00000111_00010101_00011100_0;
      patterns[1816] = 25'b00000111_00010110_00011101_0;
      patterns[1817] = 25'b00000111_00010111_00011110_0;
      patterns[1818] = 25'b00000111_00011000_00011111_0;
      patterns[1819] = 25'b00000111_00011001_00100000_0;
      patterns[1820] = 25'b00000111_00011010_00100001_0;
      patterns[1821] = 25'b00000111_00011011_00100010_0;
      patterns[1822] = 25'b00000111_00011100_00100011_0;
      patterns[1823] = 25'b00000111_00011101_00100100_0;
      patterns[1824] = 25'b00000111_00011110_00100101_0;
      patterns[1825] = 25'b00000111_00011111_00100110_0;
      patterns[1826] = 25'b00000111_00100000_00100111_0;
      patterns[1827] = 25'b00000111_00100001_00101000_0;
      patterns[1828] = 25'b00000111_00100010_00101001_0;
      patterns[1829] = 25'b00000111_00100011_00101010_0;
      patterns[1830] = 25'b00000111_00100100_00101011_0;
      patterns[1831] = 25'b00000111_00100101_00101100_0;
      patterns[1832] = 25'b00000111_00100110_00101101_0;
      patterns[1833] = 25'b00000111_00100111_00101110_0;
      patterns[1834] = 25'b00000111_00101000_00101111_0;
      patterns[1835] = 25'b00000111_00101001_00110000_0;
      patterns[1836] = 25'b00000111_00101010_00110001_0;
      patterns[1837] = 25'b00000111_00101011_00110010_0;
      patterns[1838] = 25'b00000111_00101100_00110011_0;
      patterns[1839] = 25'b00000111_00101101_00110100_0;
      patterns[1840] = 25'b00000111_00101110_00110101_0;
      patterns[1841] = 25'b00000111_00101111_00110110_0;
      patterns[1842] = 25'b00000111_00110000_00110111_0;
      patterns[1843] = 25'b00000111_00110001_00111000_0;
      patterns[1844] = 25'b00000111_00110010_00111001_0;
      patterns[1845] = 25'b00000111_00110011_00111010_0;
      patterns[1846] = 25'b00000111_00110100_00111011_0;
      patterns[1847] = 25'b00000111_00110101_00111100_0;
      patterns[1848] = 25'b00000111_00110110_00111101_0;
      patterns[1849] = 25'b00000111_00110111_00111110_0;
      patterns[1850] = 25'b00000111_00111000_00111111_0;
      patterns[1851] = 25'b00000111_00111001_01000000_0;
      patterns[1852] = 25'b00000111_00111010_01000001_0;
      patterns[1853] = 25'b00000111_00111011_01000010_0;
      patterns[1854] = 25'b00000111_00111100_01000011_0;
      patterns[1855] = 25'b00000111_00111101_01000100_0;
      patterns[1856] = 25'b00000111_00111110_01000101_0;
      patterns[1857] = 25'b00000111_00111111_01000110_0;
      patterns[1858] = 25'b00000111_01000000_01000111_0;
      patterns[1859] = 25'b00000111_01000001_01001000_0;
      patterns[1860] = 25'b00000111_01000010_01001001_0;
      patterns[1861] = 25'b00000111_01000011_01001010_0;
      patterns[1862] = 25'b00000111_01000100_01001011_0;
      patterns[1863] = 25'b00000111_01000101_01001100_0;
      patterns[1864] = 25'b00000111_01000110_01001101_0;
      patterns[1865] = 25'b00000111_01000111_01001110_0;
      patterns[1866] = 25'b00000111_01001000_01001111_0;
      patterns[1867] = 25'b00000111_01001001_01010000_0;
      patterns[1868] = 25'b00000111_01001010_01010001_0;
      patterns[1869] = 25'b00000111_01001011_01010010_0;
      patterns[1870] = 25'b00000111_01001100_01010011_0;
      patterns[1871] = 25'b00000111_01001101_01010100_0;
      patterns[1872] = 25'b00000111_01001110_01010101_0;
      patterns[1873] = 25'b00000111_01001111_01010110_0;
      patterns[1874] = 25'b00000111_01010000_01010111_0;
      patterns[1875] = 25'b00000111_01010001_01011000_0;
      patterns[1876] = 25'b00000111_01010010_01011001_0;
      patterns[1877] = 25'b00000111_01010011_01011010_0;
      patterns[1878] = 25'b00000111_01010100_01011011_0;
      patterns[1879] = 25'b00000111_01010101_01011100_0;
      patterns[1880] = 25'b00000111_01010110_01011101_0;
      patterns[1881] = 25'b00000111_01010111_01011110_0;
      patterns[1882] = 25'b00000111_01011000_01011111_0;
      patterns[1883] = 25'b00000111_01011001_01100000_0;
      patterns[1884] = 25'b00000111_01011010_01100001_0;
      patterns[1885] = 25'b00000111_01011011_01100010_0;
      patterns[1886] = 25'b00000111_01011100_01100011_0;
      patterns[1887] = 25'b00000111_01011101_01100100_0;
      patterns[1888] = 25'b00000111_01011110_01100101_0;
      patterns[1889] = 25'b00000111_01011111_01100110_0;
      patterns[1890] = 25'b00000111_01100000_01100111_0;
      patterns[1891] = 25'b00000111_01100001_01101000_0;
      patterns[1892] = 25'b00000111_01100010_01101001_0;
      patterns[1893] = 25'b00000111_01100011_01101010_0;
      patterns[1894] = 25'b00000111_01100100_01101011_0;
      patterns[1895] = 25'b00000111_01100101_01101100_0;
      patterns[1896] = 25'b00000111_01100110_01101101_0;
      patterns[1897] = 25'b00000111_01100111_01101110_0;
      patterns[1898] = 25'b00000111_01101000_01101111_0;
      patterns[1899] = 25'b00000111_01101001_01110000_0;
      patterns[1900] = 25'b00000111_01101010_01110001_0;
      patterns[1901] = 25'b00000111_01101011_01110010_0;
      patterns[1902] = 25'b00000111_01101100_01110011_0;
      patterns[1903] = 25'b00000111_01101101_01110100_0;
      patterns[1904] = 25'b00000111_01101110_01110101_0;
      patterns[1905] = 25'b00000111_01101111_01110110_0;
      patterns[1906] = 25'b00000111_01110000_01110111_0;
      patterns[1907] = 25'b00000111_01110001_01111000_0;
      patterns[1908] = 25'b00000111_01110010_01111001_0;
      patterns[1909] = 25'b00000111_01110011_01111010_0;
      patterns[1910] = 25'b00000111_01110100_01111011_0;
      patterns[1911] = 25'b00000111_01110101_01111100_0;
      patterns[1912] = 25'b00000111_01110110_01111101_0;
      patterns[1913] = 25'b00000111_01110111_01111110_0;
      patterns[1914] = 25'b00000111_01111000_01111111_0;
      patterns[1915] = 25'b00000111_01111001_10000000_0;
      patterns[1916] = 25'b00000111_01111010_10000001_0;
      patterns[1917] = 25'b00000111_01111011_10000010_0;
      patterns[1918] = 25'b00000111_01111100_10000011_0;
      patterns[1919] = 25'b00000111_01111101_10000100_0;
      patterns[1920] = 25'b00000111_01111110_10000101_0;
      patterns[1921] = 25'b00000111_01111111_10000110_0;
      patterns[1922] = 25'b00000111_10000000_10000111_0;
      patterns[1923] = 25'b00000111_10000001_10001000_0;
      patterns[1924] = 25'b00000111_10000010_10001001_0;
      patterns[1925] = 25'b00000111_10000011_10001010_0;
      patterns[1926] = 25'b00000111_10000100_10001011_0;
      patterns[1927] = 25'b00000111_10000101_10001100_0;
      patterns[1928] = 25'b00000111_10000110_10001101_0;
      patterns[1929] = 25'b00000111_10000111_10001110_0;
      patterns[1930] = 25'b00000111_10001000_10001111_0;
      patterns[1931] = 25'b00000111_10001001_10010000_0;
      patterns[1932] = 25'b00000111_10001010_10010001_0;
      patterns[1933] = 25'b00000111_10001011_10010010_0;
      patterns[1934] = 25'b00000111_10001100_10010011_0;
      patterns[1935] = 25'b00000111_10001101_10010100_0;
      patterns[1936] = 25'b00000111_10001110_10010101_0;
      patterns[1937] = 25'b00000111_10001111_10010110_0;
      patterns[1938] = 25'b00000111_10010000_10010111_0;
      patterns[1939] = 25'b00000111_10010001_10011000_0;
      patterns[1940] = 25'b00000111_10010010_10011001_0;
      patterns[1941] = 25'b00000111_10010011_10011010_0;
      patterns[1942] = 25'b00000111_10010100_10011011_0;
      patterns[1943] = 25'b00000111_10010101_10011100_0;
      patterns[1944] = 25'b00000111_10010110_10011101_0;
      patterns[1945] = 25'b00000111_10010111_10011110_0;
      patterns[1946] = 25'b00000111_10011000_10011111_0;
      patterns[1947] = 25'b00000111_10011001_10100000_0;
      patterns[1948] = 25'b00000111_10011010_10100001_0;
      patterns[1949] = 25'b00000111_10011011_10100010_0;
      patterns[1950] = 25'b00000111_10011100_10100011_0;
      patterns[1951] = 25'b00000111_10011101_10100100_0;
      patterns[1952] = 25'b00000111_10011110_10100101_0;
      patterns[1953] = 25'b00000111_10011111_10100110_0;
      patterns[1954] = 25'b00000111_10100000_10100111_0;
      patterns[1955] = 25'b00000111_10100001_10101000_0;
      patterns[1956] = 25'b00000111_10100010_10101001_0;
      patterns[1957] = 25'b00000111_10100011_10101010_0;
      patterns[1958] = 25'b00000111_10100100_10101011_0;
      patterns[1959] = 25'b00000111_10100101_10101100_0;
      patterns[1960] = 25'b00000111_10100110_10101101_0;
      patterns[1961] = 25'b00000111_10100111_10101110_0;
      patterns[1962] = 25'b00000111_10101000_10101111_0;
      patterns[1963] = 25'b00000111_10101001_10110000_0;
      patterns[1964] = 25'b00000111_10101010_10110001_0;
      patterns[1965] = 25'b00000111_10101011_10110010_0;
      patterns[1966] = 25'b00000111_10101100_10110011_0;
      patterns[1967] = 25'b00000111_10101101_10110100_0;
      patterns[1968] = 25'b00000111_10101110_10110101_0;
      patterns[1969] = 25'b00000111_10101111_10110110_0;
      patterns[1970] = 25'b00000111_10110000_10110111_0;
      patterns[1971] = 25'b00000111_10110001_10111000_0;
      patterns[1972] = 25'b00000111_10110010_10111001_0;
      patterns[1973] = 25'b00000111_10110011_10111010_0;
      patterns[1974] = 25'b00000111_10110100_10111011_0;
      patterns[1975] = 25'b00000111_10110101_10111100_0;
      patterns[1976] = 25'b00000111_10110110_10111101_0;
      patterns[1977] = 25'b00000111_10110111_10111110_0;
      patterns[1978] = 25'b00000111_10111000_10111111_0;
      patterns[1979] = 25'b00000111_10111001_11000000_0;
      patterns[1980] = 25'b00000111_10111010_11000001_0;
      patterns[1981] = 25'b00000111_10111011_11000010_0;
      patterns[1982] = 25'b00000111_10111100_11000011_0;
      patterns[1983] = 25'b00000111_10111101_11000100_0;
      patterns[1984] = 25'b00000111_10111110_11000101_0;
      patterns[1985] = 25'b00000111_10111111_11000110_0;
      patterns[1986] = 25'b00000111_11000000_11000111_0;
      patterns[1987] = 25'b00000111_11000001_11001000_0;
      patterns[1988] = 25'b00000111_11000010_11001001_0;
      patterns[1989] = 25'b00000111_11000011_11001010_0;
      patterns[1990] = 25'b00000111_11000100_11001011_0;
      patterns[1991] = 25'b00000111_11000101_11001100_0;
      patterns[1992] = 25'b00000111_11000110_11001101_0;
      patterns[1993] = 25'b00000111_11000111_11001110_0;
      patterns[1994] = 25'b00000111_11001000_11001111_0;
      patterns[1995] = 25'b00000111_11001001_11010000_0;
      patterns[1996] = 25'b00000111_11001010_11010001_0;
      patterns[1997] = 25'b00000111_11001011_11010010_0;
      patterns[1998] = 25'b00000111_11001100_11010011_0;
      patterns[1999] = 25'b00000111_11001101_11010100_0;
      patterns[2000] = 25'b00000111_11001110_11010101_0;
      patterns[2001] = 25'b00000111_11001111_11010110_0;
      patterns[2002] = 25'b00000111_11010000_11010111_0;
      patterns[2003] = 25'b00000111_11010001_11011000_0;
      patterns[2004] = 25'b00000111_11010010_11011001_0;
      patterns[2005] = 25'b00000111_11010011_11011010_0;
      patterns[2006] = 25'b00000111_11010100_11011011_0;
      patterns[2007] = 25'b00000111_11010101_11011100_0;
      patterns[2008] = 25'b00000111_11010110_11011101_0;
      patterns[2009] = 25'b00000111_11010111_11011110_0;
      patterns[2010] = 25'b00000111_11011000_11011111_0;
      patterns[2011] = 25'b00000111_11011001_11100000_0;
      patterns[2012] = 25'b00000111_11011010_11100001_0;
      patterns[2013] = 25'b00000111_11011011_11100010_0;
      patterns[2014] = 25'b00000111_11011100_11100011_0;
      patterns[2015] = 25'b00000111_11011101_11100100_0;
      patterns[2016] = 25'b00000111_11011110_11100101_0;
      patterns[2017] = 25'b00000111_11011111_11100110_0;
      patterns[2018] = 25'b00000111_11100000_11100111_0;
      patterns[2019] = 25'b00000111_11100001_11101000_0;
      patterns[2020] = 25'b00000111_11100010_11101001_0;
      patterns[2021] = 25'b00000111_11100011_11101010_0;
      patterns[2022] = 25'b00000111_11100100_11101011_0;
      patterns[2023] = 25'b00000111_11100101_11101100_0;
      patterns[2024] = 25'b00000111_11100110_11101101_0;
      patterns[2025] = 25'b00000111_11100111_11101110_0;
      patterns[2026] = 25'b00000111_11101000_11101111_0;
      patterns[2027] = 25'b00000111_11101001_11110000_0;
      patterns[2028] = 25'b00000111_11101010_11110001_0;
      patterns[2029] = 25'b00000111_11101011_11110010_0;
      patterns[2030] = 25'b00000111_11101100_11110011_0;
      patterns[2031] = 25'b00000111_11101101_11110100_0;
      patterns[2032] = 25'b00000111_11101110_11110101_0;
      patterns[2033] = 25'b00000111_11101111_11110110_0;
      patterns[2034] = 25'b00000111_11110000_11110111_0;
      patterns[2035] = 25'b00000111_11110001_11111000_0;
      patterns[2036] = 25'b00000111_11110010_11111001_0;
      patterns[2037] = 25'b00000111_11110011_11111010_0;
      patterns[2038] = 25'b00000111_11110100_11111011_0;
      patterns[2039] = 25'b00000111_11110101_11111100_0;
      patterns[2040] = 25'b00000111_11110110_11111101_0;
      patterns[2041] = 25'b00000111_11110111_11111110_0;
      patterns[2042] = 25'b00000111_11111000_11111111_0;
      patterns[2043] = 25'b00000111_11111001_00000000_1;
      patterns[2044] = 25'b00000111_11111010_00000001_1;
      patterns[2045] = 25'b00000111_11111011_00000010_1;
      patterns[2046] = 25'b00000111_11111100_00000011_1;
      patterns[2047] = 25'b00000111_11111101_00000100_1;
      patterns[2048] = 25'b00000111_11111110_00000101_1;
      patterns[2049] = 25'b00000111_11111111_00000110_1;
      patterns[2050] = 25'b00001000_00000000_00001000_0;
      patterns[2051] = 25'b00001000_00000001_00001001_0;
      patterns[2052] = 25'b00001000_00000010_00001010_0;
      patterns[2053] = 25'b00001000_00000011_00001011_0;
      patterns[2054] = 25'b00001000_00000100_00001100_0;
      patterns[2055] = 25'b00001000_00000101_00001101_0;
      patterns[2056] = 25'b00001000_00000110_00001110_0;
      patterns[2057] = 25'b00001000_00000111_00001111_0;
      patterns[2058] = 25'b00001000_00001000_00010000_0;
      patterns[2059] = 25'b00001000_00001001_00010001_0;
      patterns[2060] = 25'b00001000_00001010_00010010_0;
      patterns[2061] = 25'b00001000_00001011_00010011_0;
      patterns[2062] = 25'b00001000_00001100_00010100_0;
      patterns[2063] = 25'b00001000_00001101_00010101_0;
      patterns[2064] = 25'b00001000_00001110_00010110_0;
      patterns[2065] = 25'b00001000_00001111_00010111_0;
      patterns[2066] = 25'b00001000_00010000_00011000_0;
      patterns[2067] = 25'b00001000_00010001_00011001_0;
      patterns[2068] = 25'b00001000_00010010_00011010_0;
      patterns[2069] = 25'b00001000_00010011_00011011_0;
      patterns[2070] = 25'b00001000_00010100_00011100_0;
      patterns[2071] = 25'b00001000_00010101_00011101_0;
      patterns[2072] = 25'b00001000_00010110_00011110_0;
      patterns[2073] = 25'b00001000_00010111_00011111_0;
      patterns[2074] = 25'b00001000_00011000_00100000_0;
      patterns[2075] = 25'b00001000_00011001_00100001_0;
      patterns[2076] = 25'b00001000_00011010_00100010_0;
      patterns[2077] = 25'b00001000_00011011_00100011_0;
      patterns[2078] = 25'b00001000_00011100_00100100_0;
      patterns[2079] = 25'b00001000_00011101_00100101_0;
      patterns[2080] = 25'b00001000_00011110_00100110_0;
      patterns[2081] = 25'b00001000_00011111_00100111_0;
      patterns[2082] = 25'b00001000_00100000_00101000_0;
      patterns[2083] = 25'b00001000_00100001_00101001_0;
      patterns[2084] = 25'b00001000_00100010_00101010_0;
      patterns[2085] = 25'b00001000_00100011_00101011_0;
      patterns[2086] = 25'b00001000_00100100_00101100_0;
      patterns[2087] = 25'b00001000_00100101_00101101_0;
      patterns[2088] = 25'b00001000_00100110_00101110_0;
      patterns[2089] = 25'b00001000_00100111_00101111_0;
      patterns[2090] = 25'b00001000_00101000_00110000_0;
      patterns[2091] = 25'b00001000_00101001_00110001_0;
      patterns[2092] = 25'b00001000_00101010_00110010_0;
      patterns[2093] = 25'b00001000_00101011_00110011_0;
      patterns[2094] = 25'b00001000_00101100_00110100_0;
      patterns[2095] = 25'b00001000_00101101_00110101_0;
      patterns[2096] = 25'b00001000_00101110_00110110_0;
      patterns[2097] = 25'b00001000_00101111_00110111_0;
      patterns[2098] = 25'b00001000_00110000_00111000_0;
      patterns[2099] = 25'b00001000_00110001_00111001_0;
      patterns[2100] = 25'b00001000_00110010_00111010_0;
      patterns[2101] = 25'b00001000_00110011_00111011_0;
      patterns[2102] = 25'b00001000_00110100_00111100_0;
      patterns[2103] = 25'b00001000_00110101_00111101_0;
      patterns[2104] = 25'b00001000_00110110_00111110_0;
      patterns[2105] = 25'b00001000_00110111_00111111_0;
      patterns[2106] = 25'b00001000_00111000_01000000_0;
      patterns[2107] = 25'b00001000_00111001_01000001_0;
      patterns[2108] = 25'b00001000_00111010_01000010_0;
      patterns[2109] = 25'b00001000_00111011_01000011_0;
      patterns[2110] = 25'b00001000_00111100_01000100_0;
      patterns[2111] = 25'b00001000_00111101_01000101_0;
      patterns[2112] = 25'b00001000_00111110_01000110_0;
      patterns[2113] = 25'b00001000_00111111_01000111_0;
      patterns[2114] = 25'b00001000_01000000_01001000_0;
      patterns[2115] = 25'b00001000_01000001_01001001_0;
      patterns[2116] = 25'b00001000_01000010_01001010_0;
      patterns[2117] = 25'b00001000_01000011_01001011_0;
      patterns[2118] = 25'b00001000_01000100_01001100_0;
      patterns[2119] = 25'b00001000_01000101_01001101_0;
      patterns[2120] = 25'b00001000_01000110_01001110_0;
      patterns[2121] = 25'b00001000_01000111_01001111_0;
      patterns[2122] = 25'b00001000_01001000_01010000_0;
      patterns[2123] = 25'b00001000_01001001_01010001_0;
      patterns[2124] = 25'b00001000_01001010_01010010_0;
      patterns[2125] = 25'b00001000_01001011_01010011_0;
      patterns[2126] = 25'b00001000_01001100_01010100_0;
      patterns[2127] = 25'b00001000_01001101_01010101_0;
      patterns[2128] = 25'b00001000_01001110_01010110_0;
      patterns[2129] = 25'b00001000_01001111_01010111_0;
      patterns[2130] = 25'b00001000_01010000_01011000_0;
      patterns[2131] = 25'b00001000_01010001_01011001_0;
      patterns[2132] = 25'b00001000_01010010_01011010_0;
      patterns[2133] = 25'b00001000_01010011_01011011_0;
      patterns[2134] = 25'b00001000_01010100_01011100_0;
      patterns[2135] = 25'b00001000_01010101_01011101_0;
      patterns[2136] = 25'b00001000_01010110_01011110_0;
      patterns[2137] = 25'b00001000_01010111_01011111_0;
      patterns[2138] = 25'b00001000_01011000_01100000_0;
      patterns[2139] = 25'b00001000_01011001_01100001_0;
      patterns[2140] = 25'b00001000_01011010_01100010_0;
      patterns[2141] = 25'b00001000_01011011_01100011_0;
      patterns[2142] = 25'b00001000_01011100_01100100_0;
      patterns[2143] = 25'b00001000_01011101_01100101_0;
      patterns[2144] = 25'b00001000_01011110_01100110_0;
      patterns[2145] = 25'b00001000_01011111_01100111_0;
      patterns[2146] = 25'b00001000_01100000_01101000_0;
      patterns[2147] = 25'b00001000_01100001_01101001_0;
      patterns[2148] = 25'b00001000_01100010_01101010_0;
      patterns[2149] = 25'b00001000_01100011_01101011_0;
      patterns[2150] = 25'b00001000_01100100_01101100_0;
      patterns[2151] = 25'b00001000_01100101_01101101_0;
      patterns[2152] = 25'b00001000_01100110_01101110_0;
      patterns[2153] = 25'b00001000_01100111_01101111_0;
      patterns[2154] = 25'b00001000_01101000_01110000_0;
      patterns[2155] = 25'b00001000_01101001_01110001_0;
      patterns[2156] = 25'b00001000_01101010_01110010_0;
      patterns[2157] = 25'b00001000_01101011_01110011_0;
      patterns[2158] = 25'b00001000_01101100_01110100_0;
      patterns[2159] = 25'b00001000_01101101_01110101_0;
      patterns[2160] = 25'b00001000_01101110_01110110_0;
      patterns[2161] = 25'b00001000_01101111_01110111_0;
      patterns[2162] = 25'b00001000_01110000_01111000_0;
      patterns[2163] = 25'b00001000_01110001_01111001_0;
      patterns[2164] = 25'b00001000_01110010_01111010_0;
      patterns[2165] = 25'b00001000_01110011_01111011_0;
      patterns[2166] = 25'b00001000_01110100_01111100_0;
      patterns[2167] = 25'b00001000_01110101_01111101_0;
      patterns[2168] = 25'b00001000_01110110_01111110_0;
      patterns[2169] = 25'b00001000_01110111_01111111_0;
      patterns[2170] = 25'b00001000_01111000_10000000_0;
      patterns[2171] = 25'b00001000_01111001_10000001_0;
      patterns[2172] = 25'b00001000_01111010_10000010_0;
      patterns[2173] = 25'b00001000_01111011_10000011_0;
      patterns[2174] = 25'b00001000_01111100_10000100_0;
      patterns[2175] = 25'b00001000_01111101_10000101_0;
      patterns[2176] = 25'b00001000_01111110_10000110_0;
      patterns[2177] = 25'b00001000_01111111_10000111_0;
      patterns[2178] = 25'b00001000_10000000_10001000_0;
      patterns[2179] = 25'b00001000_10000001_10001001_0;
      patterns[2180] = 25'b00001000_10000010_10001010_0;
      patterns[2181] = 25'b00001000_10000011_10001011_0;
      patterns[2182] = 25'b00001000_10000100_10001100_0;
      patterns[2183] = 25'b00001000_10000101_10001101_0;
      patterns[2184] = 25'b00001000_10000110_10001110_0;
      patterns[2185] = 25'b00001000_10000111_10001111_0;
      patterns[2186] = 25'b00001000_10001000_10010000_0;
      patterns[2187] = 25'b00001000_10001001_10010001_0;
      patterns[2188] = 25'b00001000_10001010_10010010_0;
      patterns[2189] = 25'b00001000_10001011_10010011_0;
      patterns[2190] = 25'b00001000_10001100_10010100_0;
      patterns[2191] = 25'b00001000_10001101_10010101_0;
      patterns[2192] = 25'b00001000_10001110_10010110_0;
      patterns[2193] = 25'b00001000_10001111_10010111_0;
      patterns[2194] = 25'b00001000_10010000_10011000_0;
      patterns[2195] = 25'b00001000_10010001_10011001_0;
      patterns[2196] = 25'b00001000_10010010_10011010_0;
      patterns[2197] = 25'b00001000_10010011_10011011_0;
      patterns[2198] = 25'b00001000_10010100_10011100_0;
      patterns[2199] = 25'b00001000_10010101_10011101_0;
      patterns[2200] = 25'b00001000_10010110_10011110_0;
      patterns[2201] = 25'b00001000_10010111_10011111_0;
      patterns[2202] = 25'b00001000_10011000_10100000_0;
      patterns[2203] = 25'b00001000_10011001_10100001_0;
      patterns[2204] = 25'b00001000_10011010_10100010_0;
      patterns[2205] = 25'b00001000_10011011_10100011_0;
      patterns[2206] = 25'b00001000_10011100_10100100_0;
      patterns[2207] = 25'b00001000_10011101_10100101_0;
      patterns[2208] = 25'b00001000_10011110_10100110_0;
      patterns[2209] = 25'b00001000_10011111_10100111_0;
      patterns[2210] = 25'b00001000_10100000_10101000_0;
      patterns[2211] = 25'b00001000_10100001_10101001_0;
      patterns[2212] = 25'b00001000_10100010_10101010_0;
      patterns[2213] = 25'b00001000_10100011_10101011_0;
      patterns[2214] = 25'b00001000_10100100_10101100_0;
      patterns[2215] = 25'b00001000_10100101_10101101_0;
      patterns[2216] = 25'b00001000_10100110_10101110_0;
      patterns[2217] = 25'b00001000_10100111_10101111_0;
      patterns[2218] = 25'b00001000_10101000_10110000_0;
      patterns[2219] = 25'b00001000_10101001_10110001_0;
      patterns[2220] = 25'b00001000_10101010_10110010_0;
      patterns[2221] = 25'b00001000_10101011_10110011_0;
      patterns[2222] = 25'b00001000_10101100_10110100_0;
      patterns[2223] = 25'b00001000_10101101_10110101_0;
      patterns[2224] = 25'b00001000_10101110_10110110_0;
      patterns[2225] = 25'b00001000_10101111_10110111_0;
      patterns[2226] = 25'b00001000_10110000_10111000_0;
      patterns[2227] = 25'b00001000_10110001_10111001_0;
      patterns[2228] = 25'b00001000_10110010_10111010_0;
      patterns[2229] = 25'b00001000_10110011_10111011_0;
      patterns[2230] = 25'b00001000_10110100_10111100_0;
      patterns[2231] = 25'b00001000_10110101_10111101_0;
      patterns[2232] = 25'b00001000_10110110_10111110_0;
      patterns[2233] = 25'b00001000_10110111_10111111_0;
      patterns[2234] = 25'b00001000_10111000_11000000_0;
      patterns[2235] = 25'b00001000_10111001_11000001_0;
      patterns[2236] = 25'b00001000_10111010_11000010_0;
      patterns[2237] = 25'b00001000_10111011_11000011_0;
      patterns[2238] = 25'b00001000_10111100_11000100_0;
      patterns[2239] = 25'b00001000_10111101_11000101_0;
      patterns[2240] = 25'b00001000_10111110_11000110_0;
      patterns[2241] = 25'b00001000_10111111_11000111_0;
      patterns[2242] = 25'b00001000_11000000_11001000_0;
      patterns[2243] = 25'b00001000_11000001_11001001_0;
      patterns[2244] = 25'b00001000_11000010_11001010_0;
      patterns[2245] = 25'b00001000_11000011_11001011_0;
      patterns[2246] = 25'b00001000_11000100_11001100_0;
      patterns[2247] = 25'b00001000_11000101_11001101_0;
      patterns[2248] = 25'b00001000_11000110_11001110_0;
      patterns[2249] = 25'b00001000_11000111_11001111_0;
      patterns[2250] = 25'b00001000_11001000_11010000_0;
      patterns[2251] = 25'b00001000_11001001_11010001_0;
      patterns[2252] = 25'b00001000_11001010_11010010_0;
      patterns[2253] = 25'b00001000_11001011_11010011_0;
      patterns[2254] = 25'b00001000_11001100_11010100_0;
      patterns[2255] = 25'b00001000_11001101_11010101_0;
      patterns[2256] = 25'b00001000_11001110_11010110_0;
      patterns[2257] = 25'b00001000_11001111_11010111_0;
      patterns[2258] = 25'b00001000_11010000_11011000_0;
      patterns[2259] = 25'b00001000_11010001_11011001_0;
      patterns[2260] = 25'b00001000_11010010_11011010_0;
      patterns[2261] = 25'b00001000_11010011_11011011_0;
      patterns[2262] = 25'b00001000_11010100_11011100_0;
      patterns[2263] = 25'b00001000_11010101_11011101_0;
      patterns[2264] = 25'b00001000_11010110_11011110_0;
      patterns[2265] = 25'b00001000_11010111_11011111_0;
      patterns[2266] = 25'b00001000_11011000_11100000_0;
      patterns[2267] = 25'b00001000_11011001_11100001_0;
      patterns[2268] = 25'b00001000_11011010_11100010_0;
      patterns[2269] = 25'b00001000_11011011_11100011_0;
      patterns[2270] = 25'b00001000_11011100_11100100_0;
      patterns[2271] = 25'b00001000_11011101_11100101_0;
      patterns[2272] = 25'b00001000_11011110_11100110_0;
      patterns[2273] = 25'b00001000_11011111_11100111_0;
      patterns[2274] = 25'b00001000_11100000_11101000_0;
      patterns[2275] = 25'b00001000_11100001_11101001_0;
      patterns[2276] = 25'b00001000_11100010_11101010_0;
      patterns[2277] = 25'b00001000_11100011_11101011_0;
      patterns[2278] = 25'b00001000_11100100_11101100_0;
      patterns[2279] = 25'b00001000_11100101_11101101_0;
      patterns[2280] = 25'b00001000_11100110_11101110_0;
      patterns[2281] = 25'b00001000_11100111_11101111_0;
      patterns[2282] = 25'b00001000_11101000_11110000_0;
      patterns[2283] = 25'b00001000_11101001_11110001_0;
      patterns[2284] = 25'b00001000_11101010_11110010_0;
      patterns[2285] = 25'b00001000_11101011_11110011_0;
      patterns[2286] = 25'b00001000_11101100_11110100_0;
      patterns[2287] = 25'b00001000_11101101_11110101_0;
      patterns[2288] = 25'b00001000_11101110_11110110_0;
      patterns[2289] = 25'b00001000_11101111_11110111_0;
      patterns[2290] = 25'b00001000_11110000_11111000_0;
      patterns[2291] = 25'b00001000_11110001_11111001_0;
      patterns[2292] = 25'b00001000_11110010_11111010_0;
      patterns[2293] = 25'b00001000_11110011_11111011_0;
      patterns[2294] = 25'b00001000_11110100_11111100_0;
      patterns[2295] = 25'b00001000_11110101_11111101_0;
      patterns[2296] = 25'b00001000_11110110_11111110_0;
      patterns[2297] = 25'b00001000_11110111_11111111_0;
      patterns[2298] = 25'b00001000_11111000_00000000_1;
      patterns[2299] = 25'b00001000_11111001_00000001_1;
      patterns[2300] = 25'b00001000_11111010_00000010_1;
      patterns[2301] = 25'b00001000_11111011_00000011_1;
      patterns[2302] = 25'b00001000_11111100_00000100_1;
      patterns[2303] = 25'b00001000_11111101_00000101_1;
      patterns[2304] = 25'b00001000_11111110_00000110_1;
      patterns[2305] = 25'b00001000_11111111_00000111_1;
      patterns[2306] = 25'b00001001_00000000_00001001_0;
      patterns[2307] = 25'b00001001_00000001_00001010_0;
      patterns[2308] = 25'b00001001_00000010_00001011_0;
      patterns[2309] = 25'b00001001_00000011_00001100_0;
      patterns[2310] = 25'b00001001_00000100_00001101_0;
      patterns[2311] = 25'b00001001_00000101_00001110_0;
      patterns[2312] = 25'b00001001_00000110_00001111_0;
      patterns[2313] = 25'b00001001_00000111_00010000_0;
      patterns[2314] = 25'b00001001_00001000_00010001_0;
      patterns[2315] = 25'b00001001_00001001_00010010_0;
      patterns[2316] = 25'b00001001_00001010_00010011_0;
      patterns[2317] = 25'b00001001_00001011_00010100_0;
      patterns[2318] = 25'b00001001_00001100_00010101_0;
      patterns[2319] = 25'b00001001_00001101_00010110_0;
      patterns[2320] = 25'b00001001_00001110_00010111_0;
      patterns[2321] = 25'b00001001_00001111_00011000_0;
      patterns[2322] = 25'b00001001_00010000_00011001_0;
      patterns[2323] = 25'b00001001_00010001_00011010_0;
      patterns[2324] = 25'b00001001_00010010_00011011_0;
      patterns[2325] = 25'b00001001_00010011_00011100_0;
      patterns[2326] = 25'b00001001_00010100_00011101_0;
      patterns[2327] = 25'b00001001_00010101_00011110_0;
      patterns[2328] = 25'b00001001_00010110_00011111_0;
      patterns[2329] = 25'b00001001_00010111_00100000_0;
      patterns[2330] = 25'b00001001_00011000_00100001_0;
      patterns[2331] = 25'b00001001_00011001_00100010_0;
      patterns[2332] = 25'b00001001_00011010_00100011_0;
      patterns[2333] = 25'b00001001_00011011_00100100_0;
      patterns[2334] = 25'b00001001_00011100_00100101_0;
      patterns[2335] = 25'b00001001_00011101_00100110_0;
      patterns[2336] = 25'b00001001_00011110_00100111_0;
      patterns[2337] = 25'b00001001_00011111_00101000_0;
      patterns[2338] = 25'b00001001_00100000_00101001_0;
      patterns[2339] = 25'b00001001_00100001_00101010_0;
      patterns[2340] = 25'b00001001_00100010_00101011_0;
      patterns[2341] = 25'b00001001_00100011_00101100_0;
      patterns[2342] = 25'b00001001_00100100_00101101_0;
      patterns[2343] = 25'b00001001_00100101_00101110_0;
      patterns[2344] = 25'b00001001_00100110_00101111_0;
      patterns[2345] = 25'b00001001_00100111_00110000_0;
      patterns[2346] = 25'b00001001_00101000_00110001_0;
      patterns[2347] = 25'b00001001_00101001_00110010_0;
      patterns[2348] = 25'b00001001_00101010_00110011_0;
      patterns[2349] = 25'b00001001_00101011_00110100_0;
      patterns[2350] = 25'b00001001_00101100_00110101_0;
      patterns[2351] = 25'b00001001_00101101_00110110_0;
      patterns[2352] = 25'b00001001_00101110_00110111_0;
      patterns[2353] = 25'b00001001_00101111_00111000_0;
      patterns[2354] = 25'b00001001_00110000_00111001_0;
      patterns[2355] = 25'b00001001_00110001_00111010_0;
      patterns[2356] = 25'b00001001_00110010_00111011_0;
      patterns[2357] = 25'b00001001_00110011_00111100_0;
      patterns[2358] = 25'b00001001_00110100_00111101_0;
      patterns[2359] = 25'b00001001_00110101_00111110_0;
      patterns[2360] = 25'b00001001_00110110_00111111_0;
      patterns[2361] = 25'b00001001_00110111_01000000_0;
      patterns[2362] = 25'b00001001_00111000_01000001_0;
      patterns[2363] = 25'b00001001_00111001_01000010_0;
      patterns[2364] = 25'b00001001_00111010_01000011_0;
      patterns[2365] = 25'b00001001_00111011_01000100_0;
      patterns[2366] = 25'b00001001_00111100_01000101_0;
      patterns[2367] = 25'b00001001_00111101_01000110_0;
      patterns[2368] = 25'b00001001_00111110_01000111_0;
      patterns[2369] = 25'b00001001_00111111_01001000_0;
      patterns[2370] = 25'b00001001_01000000_01001001_0;
      patterns[2371] = 25'b00001001_01000001_01001010_0;
      patterns[2372] = 25'b00001001_01000010_01001011_0;
      patterns[2373] = 25'b00001001_01000011_01001100_0;
      patterns[2374] = 25'b00001001_01000100_01001101_0;
      patterns[2375] = 25'b00001001_01000101_01001110_0;
      patterns[2376] = 25'b00001001_01000110_01001111_0;
      patterns[2377] = 25'b00001001_01000111_01010000_0;
      patterns[2378] = 25'b00001001_01001000_01010001_0;
      patterns[2379] = 25'b00001001_01001001_01010010_0;
      patterns[2380] = 25'b00001001_01001010_01010011_0;
      patterns[2381] = 25'b00001001_01001011_01010100_0;
      patterns[2382] = 25'b00001001_01001100_01010101_0;
      patterns[2383] = 25'b00001001_01001101_01010110_0;
      patterns[2384] = 25'b00001001_01001110_01010111_0;
      patterns[2385] = 25'b00001001_01001111_01011000_0;
      patterns[2386] = 25'b00001001_01010000_01011001_0;
      patterns[2387] = 25'b00001001_01010001_01011010_0;
      patterns[2388] = 25'b00001001_01010010_01011011_0;
      patterns[2389] = 25'b00001001_01010011_01011100_0;
      patterns[2390] = 25'b00001001_01010100_01011101_0;
      patterns[2391] = 25'b00001001_01010101_01011110_0;
      patterns[2392] = 25'b00001001_01010110_01011111_0;
      patterns[2393] = 25'b00001001_01010111_01100000_0;
      patterns[2394] = 25'b00001001_01011000_01100001_0;
      patterns[2395] = 25'b00001001_01011001_01100010_0;
      patterns[2396] = 25'b00001001_01011010_01100011_0;
      patterns[2397] = 25'b00001001_01011011_01100100_0;
      patterns[2398] = 25'b00001001_01011100_01100101_0;
      patterns[2399] = 25'b00001001_01011101_01100110_0;
      patterns[2400] = 25'b00001001_01011110_01100111_0;
      patterns[2401] = 25'b00001001_01011111_01101000_0;
      patterns[2402] = 25'b00001001_01100000_01101001_0;
      patterns[2403] = 25'b00001001_01100001_01101010_0;
      patterns[2404] = 25'b00001001_01100010_01101011_0;
      patterns[2405] = 25'b00001001_01100011_01101100_0;
      patterns[2406] = 25'b00001001_01100100_01101101_0;
      patterns[2407] = 25'b00001001_01100101_01101110_0;
      patterns[2408] = 25'b00001001_01100110_01101111_0;
      patterns[2409] = 25'b00001001_01100111_01110000_0;
      patterns[2410] = 25'b00001001_01101000_01110001_0;
      patterns[2411] = 25'b00001001_01101001_01110010_0;
      patterns[2412] = 25'b00001001_01101010_01110011_0;
      patterns[2413] = 25'b00001001_01101011_01110100_0;
      patterns[2414] = 25'b00001001_01101100_01110101_0;
      patterns[2415] = 25'b00001001_01101101_01110110_0;
      patterns[2416] = 25'b00001001_01101110_01110111_0;
      patterns[2417] = 25'b00001001_01101111_01111000_0;
      patterns[2418] = 25'b00001001_01110000_01111001_0;
      patterns[2419] = 25'b00001001_01110001_01111010_0;
      patterns[2420] = 25'b00001001_01110010_01111011_0;
      patterns[2421] = 25'b00001001_01110011_01111100_0;
      patterns[2422] = 25'b00001001_01110100_01111101_0;
      patterns[2423] = 25'b00001001_01110101_01111110_0;
      patterns[2424] = 25'b00001001_01110110_01111111_0;
      patterns[2425] = 25'b00001001_01110111_10000000_0;
      patterns[2426] = 25'b00001001_01111000_10000001_0;
      patterns[2427] = 25'b00001001_01111001_10000010_0;
      patterns[2428] = 25'b00001001_01111010_10000011_0;
      patterns[2429] = 25'b00001001_01111011_10000100_0;
      patterns[2430] = 25'b00001001_01111100_10000101_0;
      patterns[2431] = 25'b00001001_01111101_10000110_0;
      patterns[2432] = 25'b00001001_01111110_10000111_0;
      patterns[2433] = 25'b00001001_01111111_10001000_0;
      patterns[2434] = 25'b00001001_10000000_10001001_0;
      patterns[2435] = 25'b00001001_10000001_10001010_0;
      patterns[2436] = 25'b00001001_10000010_10001011_0;
      patterns[2437] = 25'b00001001_10000011_10001100_0;
      patterns[2438] = 25'b00001001_10000100_10001101_0;
      patterns[2439] = 25'b00001001_10000101_10001110_0;
      patterns[2440] = 25'b00001001_10000110_10001111_0;
      patterns[2441] = 25'b00001001_10000111_10010000_0;
      patterns[2442] = 25'b00001001_10001000_10010001_0;
      patterns[2443] = 25'b00001001_10001001_10010010_0;
      patterns[2444] = 25'b00001001_10001010_10010011_0;
      patterns[2445] = 25'b00001001_10001011_10010100_0;
      patterns[2446] = 25'b00001001_10001100_10010101_0;
      patterns[2447] = 25'b00001001_10001101_10010110_0;
      patterns[2448] = 25'b00001001_10001110_10010111_0;
      patterns[2449] = 25'b00001001_10001111_10011000_0;
      patterns[2450] = 25'b00001001_10010000_10011001_0;
      patterns[2451] = 25'b00001001_10010001_10011010_0;
      patterns[2452] = 25'b00001001_10010010_10011011_0;
      patterns[2453] = 25'b00001001_10010011_10011100_0;
      patterns[2454] = 25'b00001001_10010100_10011101_0;
      patterns[2455] = 25'b00001001_10010101_10011110_0;
      patterns[2456] = 25'b00001001_10010110_10011111_0;
      patterns[2457] = 25'b00001001_10010111_10100000_0;
      patterns[2458] = 25'b00001001_10011000_10100001_0;
      patterns[2459] = 25'b00001001_10011001_10100010_0;
      patterns[2460] = 25'b00001001_10011010_10100011_0;
      patterns[2461] = 25'b00001001_10011011_10100100_0;
      patterns[2462] = 25'b00001001_10011100_10100101_0;
      patterns[2463] = 25'b00001001_10011101_10100110_0;
      patterns[2464] = 25'b00001001_10011110_10100111_0;
      patterns[2465] = 25'b00001001_10011111_10101000_0;
      patterns[2466] = 25'b00001001_10100000_10101001_0;
      patterns[2467] = 25'b00001001_10100001_10101010_0;
      patterns[2468] = 25'b00001001_10100010_10101011_0;
      patterns[2469] = 25'b00001001_10100011_10101100_0;
      patterns[2470] = 25'b00001001_10100100_10101101_0;
      patterns[2471] = 25'b00001001_10100101_10101110_0;
      patterns[2472] = 25'b00001001_10100110_10101111_0;
      patterns[2473] = 25'b00001001_10100111_10110000_0;
      patterns[2474] = 25'b00001001_10101000_10110001_0;
      patterns[2475] = 25'b00001001_10101001_10110010_0;
      patterns[2476] = 25'b00001001_10101010_10110011_0;
      patterns[2477] = 25'b00001001_10101011_10110100_0;
      patterns[2478] = 25'b00001001_10101100_10110101_0;
      patterns[2479] = 25'b00001001_10101101_10110110_0;
      patterns[2480] = 25'b00001001_10101110_10110111_0;
      patterns[2481] = 25'b00001001_10101111_10111000_0;
      patterns[2482] = 25'b00001001_10110000_10111001_0;
      patterns[2483] = 25'b00001001_10110001_10111010_0;
      patterns[2484] = 25'b00001001_10110010_10111011_0;
      patterns[2485] = 25'b00001001_10110011_10111100_0;
      patterns[2486] = 25'b00001001_10110100_10111101_0;
      patterns[2487] = 25'b00001001_10110101_10111110_0;
      patterns[2488] = 25'b00001001_10110110_10111111_0;
      patterns[2489] = 25'b00001001_10110111_11000000_0;
      patterns[2490] = 25'b00001001_10111000_11000001_0;
      patterns[2491] = 25'b00001001_10111001_11000010_0;
      patterns[2492] = 25'b00001001_10111010_11000011_0;
      patterns[2493] = 25'b00001001_10111011_11000100_0;
      patterns[2494] = 25'b00001001_10111100_11000101_0;
      patterns[2495] = 25'b00001001_10111101_11000110_0;
      patterns[2496] = 25'b00001001_10111110_11000111_0;
      patterns[2497] = 25'b00001001_10111111_11001000_0;
      patterns[2498] = 25'b00001001_11000000_11001001_0;
      patterns[2499] = 25'b00001001_11000001_11001010_0;
      patterns[2500] = 25'b00001001_11000010_11001011_0;
      patterns[2501] = 25'b00001001_11000011_11001100_0;
      patterns[2502] = 25'b00001001_11000100_11001101_0;
      patterns[2503] = 25'b00001001_11000101_11001110_0;
      patterns[2504] = 25'b00001001_11000110_11001111_0;
      patterns[2505] = 25'b00001001_11000111_11010000_0;
      patterns[2506] = 25'b00001001_11001000_11010001_0;
      patterns[2507] = 25'b00001001_11001001_11010010_0;
      patterns[2508] = 25'b00001001_11001010_11010011_0;
      patterns[2509] = 25'b00001001_11001011_11010100_0;
      patterns[2510] = 25'b00001001_11001100_11010101_0;
      patterns[2511] = 25'b00001001_11001101_11010110_0;
      patterns[2512] = 25'b00001001_11001110_11010111_0;
      patterns[2513] = 25'b00001001_11001111_11011000_0;
      patterns[2514] = 25'b00001001_11010000_11011001_0;
      patterns[2515] = 25'b00001001_11010001_11011010_0;
      patterns[2516] = 25'b00001001_11010010_11011011_0;
      patterns[2517] = 25'b00001001_11010011_11011100_0;
      patterns[2518] = 25'b00001001_11010100_11011101_0;
      patterns[2519] = 25'b00001001_11010101_11011110_0;
      patterns[2520] = 25'b00001001_11010110_11011111_0;
      patterns[2521] = 25'b00001001_11010111_11100000_0;
      patterns[2522] = 25'b00001001_11011000_11100001_0;
      patterns[2523] = 25'b00001001_11011001_11100010_0;
      patterns[2524] = 25'b00001001_11011010_11100011_0;
      patterns[2525] = 25'b00001001_11011011_11100100_0;
      patterns[2526] = 25'b00001001_11011100_11100101_0;
      patterns[2527] = 25'b00001001_11011101_11100110_0;
      patterns[2528] = 25'b00001001_11011110_11100111_0;
      patterns[2529] = 25'b00001001_11011111_11101000_0;
      patterns[2530] = 25'b00001001_11100000_11101001_0;
      patterns[2531] = 25'b00001001_11100001_11101010_0;
      patterns[2532] = 25'b00001001_11100010_11101011_0;
      patterns[2533] = 25'b00001001_11100011_11101100_0;
      patterns[2534] = 25'b00001001_11100100_11101101_0;
      patterns[2535] = 25'b00001001_11100101_11101110_0;
      patterns[2536] = 25'b00001001_11100110_11101111_0;
      patterns[2537] = 25'b00001001_11100111_11110000_0;
      patterns[2538] = 25'b00001001_11101000_11110001_0;
      patterns[2539] = 25'b00001001_11101001_11110010_0;
      patterns[2540] = 25'b00001001_11101010_11110011_0;
      patterns[2541] = 25'b00001001_11101011_11110100_0;
      patterns[2542] = 25'b00001001_11101100_11110101_0;
      patterns[2543] = 25'b00001001_11101101_11110110_0;
      patterns[2544] = 25'b00001001_11101110_11110111_0;
      patterns[2545] = 25'b00001001_11101111_11111000_0;
      patterns[2546] = 25'b00001001_11110000_11111001_0;
      patterns[2547] = 25'b00001001_11110001_11111010_0;
      patterns[2548] = 25'b00001001_11110010_11111011_0;
      patterns[2549] = 25'b00001001_11110011_11111100_0;
      patterns[2550] = 25'b00001001_11110100_11111101_0;
      patterns[2551] = 25'b00001001_11110101_11111110_0;
      patterns[2552] = 25'b00001001_11110110_11111111_0;
      patterns[2553] = 25'b00001001_11110111_00000000_1;
      patterns[2554] = 25'b00001001_11111000_00000001_1;
      patterns[2555] = 25'b00001001_11111001_00000010_1;
      patterns[2556] = 25'b00001001_11111010_00000011_1;
      patterns[2557] = 25'b00001001_11111011_00000100_1;
      patterns[2558] = 25'b00001001_11111100_00000101_1;
      patterns[2559] = 25'b00001001_11111101_00000110_1;
      patterns[2560] = 25'b00001001_11111110_00000111_1;
      patterns[2561] = 25'b00001001_11111111_00001000_1;
      patterns[2562] = 25'b00001010_00000000_00001010_0;
      patterns[2563] = 25'b00001010_00000001_00001011_0;
      patterns[2564] = 25'b00001010_00000010_00001100_0;
      patterns[2565] = 25'b00001010_00000011_00001101_0;
      patterns[2566] = 25'b00001010_00000100_00001110_0;
      patterns[2567] = 25'b00001010_00000101_00001111_0;
      patterns[2568] = 25'b00001010_00000110_00010000_0;
      patterns[2569] = 25'b00001010_00000111_00010001_0;
      patterns[2570] = 25'b00001010_00001000_00010010_0;
      patterns[2571] = 25'b00001010_00001001_00010011_0;
      patterns[2572] = 25'b00001010_00001010_00010100_0;
      patterns[2573] = 25'b00001010_00001011_00010101_0;
      patterns[2574] = 25'b00001010_00001100_00010110_0;
      patterns[2575] = 25'b00001010_00001101_00010111_0;
      patterns[2576] = 25'b00001010_00001110_00011000_0;
      patterns[2577] = 25'b00001010_00001111_00011001_0;
      patterns[2578] = 25'b00001010_00010000_00011010_0;
      patterns[2579] = 25'b00001010_00010001_00011011_0;
      patterns[2580] = 25'b00001010_00010010_00011100_0;
      patterns[2581] = 25'b00001010_00010011_00011101_0;
      patterns[2582] = 25'b00001010_00010100_00011110_0;
      patterns[2583] = 25'b00001010_00010101_00011111_0;
      patterns[2584] = 25'b00001010_00010110_00100000_0;
      patterns[2585] = 25'b00001010_00010111_00100001_0;
      patterns[2586] = 25'b00001010_00011000_00100010_0;
      patterns[2587] = 25'b00001010_00011001_00100011_0;
      patterns[2588] = 25'b00001010_00011010_00100100_0;
      patterns[2589] = 25'b00001010_00011011_00100101_0;
      patterns[2590] = 25'b00001010_00011100_00100110_0;
      patterns[2591] = 25'b00001010_00011101_00100111_0;
      patterns[2592] = 25'b00001010_00011110_00101000_0;
      patterns[2593] = 25'b00001010_00011111_00101001_0;
      patterns[2594] = 25'b00001010_00100000_00101010_0;
      patterns[2595] = 25'b00001010_00100001_00101011_0;
      patterns[2596] = 25'b00001010_00100010_00101100_0;
      patterns[2597] = 25'b00001010_00100011_00101101_0;
      patterns[2598] = 25'b00001010_00100100_00101110_0;
      patterns[2599] = 25'b00001010_00100101_00101111_0;
      patterns[2600] = 25'b00001010_00100110_00110000_0;
      patterns[2601] = 25'b00001010_00100111_00110001_0;
      patterns[2602] = 25'b00001010_00101000_00110010_0;
      patterns[2603] = 25'b00001010_00101001_00110011_0;
      patterns[2604] = 25'b00001010_00101010_00110100_0;
      patterns[2605] = 25'b00001010_00101011_00110101_0;
      patterns[2606] = 25'b00001010_00101100_00110110_0;
      patterns[2607] = 25'b00001010_00101101_00110111_0;
      patterns[2608] = 25'b00001010_00101110_00111000_0;
      patterns[2609] = 25'b00001010_00101111_00111001_0;
      patterns[2610] = 25'b00001010_00110000_00111010_0;
      patterns[2611] = 25'b00001010_00110001_00111011_0;
      patterns[2612] = 25'b00001010_00110010_00111100_0;
      patterns[2613] = 25'b00001010_00110011_00111101_0;
      patterns[2614] = 25'b00001010_00110100_00111110_0;
      patterns[2615] = 25'b00001010_00110101_00111111_0;
      patterns[2616] = 25'b00001010_00110110_01000000_0;
      patterns[2617] = 25'b00001010_00110111_01000001_0;
      patterns[2618] = 25'b00001010_00111000_01000010_0;
      patterns[2619] = 25'b00001010_00111001_01000011_0;
      patterns[2620] = 25'b00001010_00111010_01000100_0;
      patterns[2621] = 25'b00001010_00111011_01000101_0;
      patterns[2622] = 25'b00001010_00111100_01000110_0;
      patterns[2623] = 25'b00001010_00111101_01000111_0;
      patterns[2624] = 25'b00001010_00111110_01001000_0;
      patterns[2625] = 25'b00001010_00111111_01001001_0;
      patterns[2626] = 25'b00001010_01000000_01001010_0;
      patterns[2627] = 25'b00001010_01000001_01001011_0;
      patterns[2628] = 25'b00001010_01000010_01001100_0;
      patterns[2629] = 25'b00001010_01000011_01001101_0;
      patterns[2630] = 25'b00001010_01000100_01001110_0;
      patterns[2631] = 25'b00001010_01000101_01001111_0;
      patterns[2632] = 25'b00001010_01000110_01010000_0;
      patterns[2633] = 25'b00001010_01000111_01010001_0;
      patterns[2634] = 25'b00001010_01001000_01010010_0;
      patterns[2635] = 25'b00001010_01001001_01010011_0;
      patterns[2636] = 25'b00001010_01001010_01010100_0;
      patterns[2637] = 25'b00001010_01001011_01010101_0;
      patterns[2638] = 25'b00001010_01001100_01010110_0;
      patterns[2639] = 25'b00001010_01001101_01010111_0;
      patterns[2640] = 25'b00001010_01001110_01011000_0;
      patterns[2641] = 25'b00001010_01001111_01011001_0;
      patterns[2642] = 25'b00001010_01010000_01011010_0;
      patterns[2643] = 25'b00001010_01010001_01011011_0;
      patterns[2644] = 25'b00001010_01010010_01011100_0;
      patterns[2645] = 25'b00001010_01010011_01011101_0;
      patterns[2646] = 25'b00001010_01010100_01011110_0;
      patterns[2647] = 25'b00001010_01010101_01011111_0;
      patterns[2648] = 25'b00001010_01010110_01100000_0;
      patterns[2649] = 25'b00001010_01010111_01100001_0;
      patterns[2650] = 25'b00001010_01011000_01100010_0;
      patterns[2651] = 25'b00001010_01011001_01100011_0;
      patterns[2652] = 25'b00001010_01011010_01100100_0;
      patterns[2653] = 25'b00001010_01011011_01100101_0;
      patterns[2654] = 25'b00001010_01011100_01100110_0;
      patterns[2655] = 25'b00001010_01011101_01100111_0;
      patterns[2656] = 25'b00001010_01011110_01101000_0;
      patterns[2657] = 25'b00001010_01011111_01101001_0;
      patterns[2658] = 25'b00001010_01100000_01101010_0;
      patterns[2659] = 25'b00001010_01100001_01101011_0;
      patterns[2660] = 25'b00001010_01100010_01101100_0;
      patterns[2661] = 25'b00001010_01100011_01101101_0;
      patterns[2662] = 25'b00001010_01100100_01101110_0;
      patterns[2663] = 25'b00001010_01100101_01101111_0;
      patterns[2664] = 25'b00001010_01100110_01110000_0;
      patterns[2665] = 25'b00001010_01100111_01110001_0;
      patterns[2666] = 25'b00001010_01101000_01110010_0;
      patterns[2667] = 25'b00001010_01101001_01110011_0;
      patterns[2668] = 25'b00001010_01101010_01110100_0;
      patterns[2669] = 25'b00001010_01101011_01110101_0;
      patterns[2670] = 25'b00001010_01101100_01110110_0;
      patterns[2671] = 25'b00001010_01101101_01110111_0;
      patterns[2672] = 25'b00001010_01101110_01111000_0;
      patterns[2673] = 25'b00001010_01101111_01111001_0;
      patterns[2674] = 25'b00001010_01110000_01111010_0;
      patterns[2675] = 25'b00001010_01110001_01111011_0;
      patterns[2676] = 25'b00001010_01110010_01111100_0;
      patterns[2677] = 25'b00001010_01110011_01111101_0;
      patterns[2678] = 25'b00001010_01110100_01111110_0;
      patterns[2679] = 25'b00001010_01110101_01111111_0;
      patterns[2680] = 25'b00001010_01110110_10000000_0;
      patterns[2681] = 25'b00001010_01110111_10000001_0;
      patterns[2682] = 25'b00001010_01111000_10000010_0;
      patterns[2683] = 25'b00001010_01111001_10000011_0;
      patterns[2684] = 25'b00001010_01111010_10000100_0;
      patterns[2685] = 25'b00001010_01111011_10000101_0;
      patterns[2686] = 25'b00001010_01111100_10000110_0;
      patterns[2687] = 25'b00001010_01111101_10000111_0;
      patterns[2688] = 25'b00001010_01111110_10001000_0;
      patterns[2689] = 25'b00001010_01111111_10001001_0;
      patterns[2690] = 25'b00001010_10000000_10001010_0;
      patterns[2691] = 25'b00001010_10000001_10001011_0;
      patterns[2692] = 25'b00001010_10000010_10001100_0;
      patterns[2693] = 25'b00001010_10000011_10001101_0;
      patterns[2694] = 25'b00001010_10000100_10001110_0;
      patterns[2695] = 25'b00001010_10000101_10001111_0;
      patterns[2696] = 25'b00001010_10000110_10010000_0;
      patterns[2697] = 25'b00001010_10000111_10010001_0;
      patterns[2698] = 25'b00001010_10001000_10010010_0;
      patterns[2699] = 25'b00001010_10001001_10010011_0;
      patterns[2700] = 25'b00001010_10001010_10010100_0;
      patterns[2701] = 25'b00001010_10001011_10010101_0;
      patterns[2702] = 25'b00001010_10001100_10010110_0;
      patterns[2703] = 25'b00001010_10001101_10010111_0;
      patterns[2704] = 25'b00001010_10001110_10011000_0;
      patterns[2705] = 25'b00001010_10001111_10011001_0;
      patterns[2706] = 25'b00001010_10010000_10011010_0;
      patterns[2707] = 25'b00001010_10010001_10011011_0;
      patterns[2708] = 25'b00001010_10010010_10011100_0;
      patterns[2709] = 25'b00001010_10010011_10011101_0;
      patterns[2710] = 25'b00001010_10010100_10011110_0;
      patterns[2711] = 25'b00001010_10010101_10011111_0;
      patterns[2712] = 25'b00001010_10010110_10100000_0;
      patterns[2713] = 25'b00001010_10010111_10100001_0;
      patterns[2714] = 25'b00001010_10011000_10100010_0;
      patterns[2715] = 25'b00001010_10011001_10100011_0;
      patterns[2716] = 25'b00001010_10011010_10100100_0;
      patterns[2717] = 25'b00001010_10011011_10100101_0;
      patterns[2718] = 25'b00001010_10011100_10100110_0;
      patterns[2719] = 25'b00001010_10011101_10100111_0;
      patterns[2720] = 25'b00001010_10011110_10101000_0;
      patterns[2721] = 25'b00001010_10011111_10101001_0;
      patterns[2722] = 25'b00001010_10100000_10101010_0;
      patterns[2723] = 25'b00001010_10100001_10101011_0;
      patterns[2724] = 25'b00001010_10100010_10101100_0;
      patterns[2725] = 25'b00001010_10100011_10101101_0;
      patterns[2726] = 25'b00001010_10100100_10101110_0;
      patterns[2727] = 25'b00001010_10100101_10101111_0;
      patterns[2728] = 25'b00001010_10100110_10110000_0;
      patterns[2729] = 25'b00001010_10100111_10110001_0;
      patterns[2730] = 25'b00001010_10101000_10110010_0;
      patterns[2731] = 25'b00001010_10101001_10110011_0;
      patterns[2732] = 25'b00001010_10101010_10110100_0;
      patterns[2733] = 25'b00001010_10101011_10110101_0;
      patterns[2734] = 25'b00001010_10101100_10110110_0;
      patterns[2735] = 25'b00001010_10101101_10110111_0;
      patterns[2736] = 25'b00001010_10101110_10111000_0;
      patterns[2737] = 25'b00001010_10101111_10111001_0;
      patterns[2738] = 25'b00001010_10110000_10111010_0;
      patterns[2739] = 25'b00001010_10110001_10111011_0;
      patterns[2740] = 25'b00001010_10110010_10111100_0;
      patterns[2741] = 25'b00001010_10110011_10111101_0;
      patterns[2742] = 25'b00001010_10110100_10111110_0;
      patterns[2743] = 25'b00001010_10110101_10111111_0;
      patterns[2744] = 25'b00001010_10110110_11000000_0;
      patterns[2745] = 25'b00001010_10110111_11000001_0;
      patterns[2746] = 25'b00001010_10111000_11000010_0;
      patterns[2747] = 25'b00001010_10111001_11000011_0;
      patterns[2748] = 25'b00001010_10111010_11000100_0;
      patterns[2749] = 25'b00001010_10111011_11000101_0;
      patterns[2750] = 25'b00001010_10111100_11000110_0;
      patterns[2751] = 25'b00001010_10111101_11000111_0;
      patterns[2752] = 25'b00001010_10111110_11001000_0;
      patterns[2753] = 25'b00001010_10111111_11001001_0;
      patterns[2754] = 25'b00001010_11000000_11001010_0;
      patterns[2755] = 25'b00001010_11000001_11001011_0;
      patterns[2756] = 25'b00001010_11000010_11001100_0;
      patterns[2757] = 25'b00001010_11000011_11001101_0;
      patterns[2758] = 25'b00001010_11000100_11001110_0;
      patterns[2759] = 25'b00001010_11000101_11001111_0;
      patterns[2760] = 25'b00001010_11000110_11010000_0;
      patterns[2761] = 25'b00001010_11000111_11010001_0;
      patterns[2762] = 25'b00001010_11001000_11010010_0;
      patterns[2763] = 25'b00001010_11001001_11010011_0;
      patterns[2764] = 25'b00001010_11001010_11010100_0;
      patterns[2765] = 25'b00001010_11001011_11010101_0;
      patterns[2766] = 25'b00001010_11001100_11010110_0;
      patterns[2767] = 25'b00001010_11001101_11010111_0;
      patterns[2768] = 25'b00001010_11001110_11011000_0;
      patterns[2769] = 25'b00001010_11001111_11011001_0;
      patterns[2770] = 25'b00001010_11010000_11011010_0;
      patterns[2771] = 25'b00001010_11010001_11011011_0;
      patterns[2772] = 25'b00001010_11010010_11011100_0;
      patterns[2773] = 25'b00001010_11010011_11011101_0;
      patterns[2774] = 25'b00001010_11010100_11011110_0;
      patterns[2775] = 25'b00001010_11010101_11011111_0;
      patterns[2776] = 25'b00001010_11010110_11100000_0;
      patterns[2777] = 25'b00001010_11010111_11100001_0;
      patterns[2778] = 25'b00001010_11011000_11100010_0;
      patterns[2779] = 25'b00001010_11011001_11100011_0;
      patterns[2780] = 25'b00001010_11011010_11100100_0;
      patterns[2781] = 25'b00001010_11011011_11100101_0;
      patterns[2782] = 25'b00001010_11011100_11100110_0;
      patterns[2783] = 25'b00001010_11011101_11100111_0;
      patterns[2784] = 25'b00001010_11011110_11101000_0;
      patterns[2785] = 25'b00001010_11011111_11101001_0;
      patterns[2786] = 25'b00001010_11100000_11101010_0;
      patterns[2787] = 25'b00001010_11100001_11101011_0;
      patterns[2788] = 25'b00001010_11100010_11101100_0;
      patterns[2789] = 25'b00001010_11100011_11101101_0;
      patterns[2790] = 25'b00001010_11100100_11101110_0;
      patterns[2791] = 25'b00001010_11100101_11101111_0;
      patterns[2792] = 25'b00001010_11100110_11110000_0;
      patterns[2793] = 25'b00001010_11100111_11110001_0;
      patterns[2794] = 25'b00001010_11101000_11110010_0;
      patterns[2795] = 25'b00001010_11101001_11110011_0;
      patterns[2796] = 25'b00001010_11101010_11110100_0;
      patterns[2797] = 25'b00001010_11101011_11110101_0;
      patterns[2798] = 25'b00001010_11101100_11110110_0;
      patterns[2799] = 25'b00001010_11101101_11110111_0;
      patterns[2800] = 25'b00001010_11101110_11111000_0;
      patterns[2801] = 25'b00001010_11101111_11111001_0;
      patterns[2802] = 25'b00001010_11110000_11111010_0;
      patterns[2803] = 25'b00001010_11110001_11111011_0;
      patterns[2804] = 25'b00001010_11110010_11111100_0;
      patterns[2805] = 25'b00001010_11110011_11111101_0;
      patterns[2806] = 25'b00001010_11110100_11111110_0;
      patterns[2807] = 25'b00001010_11110101_11111111_0;
      patterns[2808] = 25'b00001010_11110110_00000000_1;
      patterns[2809] = 25'b00001010_11110111_00000001_1;
      patterns[2810] = 25'b00001010_11111000_00000010_1;
      patterns[2811] = 25'b00001010_11111001_00000011_1;
      patterns[2812] = 25'b00001010_11111010_00000100_1;
      patterns[2813] = 25'b00001010_11111011_00000101_1;
      patterns[2814] = 25'b00001010_11111100_00000110_1;
      patterns[2815] = 25'b00001010_11111101_00000111_1;
      patterns[2816] = 25'b00001010_11111110_00001000_1;
      patterns[2817] = 25'b00001010_11111111_00001001_1;
      patterns[2818] = 25'b00001011_00000000_00001011_0;
      patterns[2819] = 25'b00001011_00000001_00001100_0;
      patterns[2820] = 25'b00001011_00000010_00001101_0;
      patterns[2821] = 25'b00001011_00000011_00001110_0;
      patterns[2822] = 25'b00001011_00000100_00001111_0;
      patterns[2823] = 25'b00001011_00000101_00010000_0;
      patterns[2824] = 25'b00001011_00000110_00010001_0;
      patterns[2825] = 25'b00001011_00000111_00010010_0;
      patterns[2826] = 25'b00001011_00001000_00010011_0;
      patterns[2827] = 25'b00001011_00001001_00010100_0;
      patterns[2828] = 25'b00001011_00001010_00010101_0;
      patterns[2829] = 25'b00001011_00001011_00010110_0;
      patterns[2830] = 25'b00001011_00001100_00010111_0;
      patterns[2831] = 25'b00001011_00001101_00011000_0;
      patterns[2832] = 25'b00001011_00001110_00011001_0;
      patterns[2833] = 25'b00001011_00001111_00011010_0;
      patterns[2834] = 25'b00001011_00010000_00011011_0;
      patterns[2835] = 25'b00001011_00010001_00011100_0;
      patterns[2836] = 25'b00001011_00010010_00011101_0;
      patterns[2837] = 25'b00001011_00010011_00011110_0;
      patterns[2838] = 25'b00001011_00010100_00011111_0;
      patterns[2839] = 25'b00001011_00010101_00100000_0;
      patterns[2840] = 25'b00001011_00010110_00100001_0;
      patterns[2841] = 25'b00001011_00010111_00100010_0;
      patterns[2842] = 25'b00001011_00011000_00100011_0;
      patterns[2843] = 25'b00001011_00011001_00100100_0;
      patterns[2844] = 25'b00001011_00011010_00100101_0;
      patterns[2845] = 25'b00001011_00011011_00100110_0;
      patterns[2846] = 25'b00001011_00011100_00100111_0;
      patterns[2847] = 25'b00001011_00011101_00101000_0;
      patterns[2848] = 25'b00001011_00011110_00101001_0;
      patterns[2849] = 25'b00001011_00011111_00101010_0;
      patterns[2850] = 25'b00001011_00100000_00101011_0;
      patterns[2851] = 25'b00001011_00100001_00101100_0;
      patterns[2852] = 25'b00001011_00100010_00101101_0;
      patterns[2853] = 25'b00001011_00100011_00101110_0;
      patterns[2854] = 25'b00001011_00100100_00101111_0;
      patterns[2855] = 25'b00001011_00100101_00110000_0;
      patterns[2856] = 25'b00001011_00100110_00110001_0;
      patterns[2857] = 25'b00001011_00100111_00110010_0;
      patterns[2858] = 25'b00001011_00101000_00110011_0;
      patterns[2859] = 25'b00001011_00101001_00110100_0;
      patterns[2860] = 25'b00001011_00101010_00110101_0;
      patterns[2861] = 25'b00001011_00101011_00110110_0;
      patterns[2862] = 25'b00001011_00101100_00110111_0;
      patterns[2863] = 25'b00001011_00101101_00111000_0;
      patterns[2864] = 25'b00001011_00101110_00111001_0;
      patterns[2865] = 25'b00001011_00101111_00111010_0;
      patterns[2866] = 25'b00001011_00110000_00111011_0;
      patterns[2867] = 25'b00001011_00110001_00111100_0;
      patterns[2868] = 25'b00001011_00110010_00111101_0;
      patterns[2869] = 25'b00001011_00110011_00111110_0;
      patterns[2870] = 25'b00001011_00110100_00111111_0;
      patterns[2871] = 25'b00001011_00110101_01000000_0;
      patterns[2872] = 25'b00001011_00110110_01000001_0;
      patterns[2873] = 25'b00001011_00110111_01000010_0;
      patterns[2874] = 25'b00001011_00111000_01000011_0;
      patterns[2875] = 25'b00001011_00111001_01000100_0;
      patterns[2876] = 25'b00001011_00111010_01000101_0;
      patterns[2877] = 25'b00001011_00111011_01000110_0;
      patterns[2878] = 25'b00001011_00111100_01000111_0;
      patterns[2879] = 25'b00001011_00111101_01001000_0;
      patterns[2880] = 25'b00001011_00111110_01001001_0;
      patterns[2881] = 25'b00001011_00111111_01001010_0;
      patterns[2882] = 25'b00001011_01000000_01001011_0;
      patterns[2883] = 25'b00001011_01000001_01001100_0;
      patterns[2884] = 25'b00001011_01000010_01001101_0;
      patterns[2885] = 25'b00001011_01000011_01001110_0;
      patterns[2886] = 25'b00001011_01000100_01001111_0;
      patterns[2887] = 25'b00001011_01000101_01010000_0;
      patterns[2888] = 25'b00001011_01000110_01010001_0;
      patterns[2889] = 25'b00001011_01000111_01010010_0;
      patterns[2890] = 25'b00001011_01001000_01010011_0;
      patterns[2891] = 25'b00001011_01001001_01010100_0;
      patterns[2892] = 25'b00001011_01001010_01010101_0;
      patterns[2893] = 25'b00001011_01001011_01010110_0;
      patterns[2894] = 25'b00001011_01001100_01010111_0;
      patterns[2895] = 25'b00001011_01001101_01011000_0;
      patterns[2896] = 25'b00001011_01001110_01011001_0;
      patterns[2897] = 25'b00001011_01001111_01011010_0;
      patterns[2898] = 25'b00001011_01010000_01011011_0;
      patterns[2899] = 25'b00001011_01010001_01011100_0;
      patterns[2900] = 25'b00001011_01010010_01011101_0;
      patterns[2901] = 25'b00001011_01010011_01011110_0;
      patterns[2902] = 25'b00001011_01010100_01011111_0;
      patterns[2903] = 25'b00001011_01010101_01100000_0;
      patterns[2904] = 25'b00001011_01010110_01100001_0;
      patterns[2905] = 25'b00001011_01010111_01100010_0;
      patterns[2906] = 25'b00001011_01011000_01100011_0;
      patterns[2907] = 25'b00001011_01011001_01100100_0;
      patterns[2908] = 25'b00001011_01011010_01100101_0;
      patterns[2909] = 25'b00001011_01011011_01100110_0;
      patterns[2910] = 25'b00001011_01011100_01100111_0;
      patterns[2911] = 25'b00001011_01011101_01101000_0;
      patterns[2912] = 25'b00001011_01011110_01101001_0;
      patterns[2913] = 25'b00001011_01011111_01101010_0;
      patterns[2914] = 25'b00001011_01100000_01101011_0;
      patterns[2915] = 25'b00001011_01100001_01101100_0;
      patterns[2916] = 25'b00001011_01100010_01101101_0;
      patterns[2917] = 25'b00001011_01100011_01101110_0;
      patterns[2918] = 25'b00001011_01100100_01101111_0;
      patterns[2919] = 25'b00001011_01100101_01110000_0;
      patterns[2920] = 25'b00001011_01100110_01110001_0;
      patterns[2921] = 25'b00001011_01100111_01110010_0;
      patterns[2922] = 25'b00001011_01101000_01110011_0;
      patterns[2923] = 25'b00001011_01101001_01110100_0;
      patterns[2924] = 25'b00001011_01101010_01110101_0;
      patterns[2925] = 25'b00001011_01101011_01110110_0;
      patterns[2926] = 25'b00001011_01101100_01110111_0;
      patterns[2927] = 25'b00001011_01101101_01111000_0;
      patterns[2928] = 25'b00001011_01101110_01111001_0;
      patterns[2929] = 25'b00001011_01101111_01111010_0;
      patterns[2930] = 25'b00001011_01110000_01111011_0;
      patterns[2931] = 25'b00001011_01110001_01111100_0;
      patterns[2932] = 25'b00001011_01110010_01111101_0;
      patterns[2933] = 25'b00001011_01110011_01111110_0;
      patterns[2934] = 25'b00001011_01110100_01111111_0;
      patterns[2935] = 25'b00001011_01110101_10000000_0;
      patterns[2936] = 25'b00001011_01110110_10000001_0;
      patterns[2937] = 25'b00001011_01110111_10000010_0;
      patterns[2938] = 25'b00001011_01111000_10000011_0;
      patterns[2939] = 25'b00001011_01111001_10000100_0;
      patterns[2940] = 25'b00001011_01111010_10000101_0;
      patterns[2941] = 25'b00001011_01111011_10000110_0;
      patterns[2942] = 25'b00001011_01111100_10000111_0;
      patterns[2943] = 25'b00001011_01111101_10001000_0;
      patterns[2944] = 25'b00001011_01111110_10001001_0;
      patterns[2945] = 25'b00001011_01111111_10001010_0;
      patterns[2946] = 25'b00001011_10000000_10001011_0;
      patterns[2947] = 25'b00001011_10000001_10001100_0;
      patterns[2948] = 25'b00001011_10000010_10001101_0;
      patterns[2949] = 25'b00001011_10000011_10001110_0;
      patterns[2950] = 25'b00001011_10000100_10001111_0;
      patterns[2951] = 25'b00001011_10000101_10010000_0;
      patterns[2952] = 25'b00001011_10000110_10010001_0;
      patterns[2953] = 25'b00001011_10000111_10010010_0;
      patterns[2954] = 25'b00001011_10001000_10010011_0;
      patterns[2955] = 25'b00001011_10001001_10010100_0;
      patterns[2956] = 25'b00001011_10001010_10010101_0;
      patterns[2957] = 25'b00001011_10001011_10010110_0;
      patterns[2958] = 25'b00001011_10001100_10010111_0;
      patterns[2959] = 25'b00001011_10001101_10011000_0;
      patterns[2960] = 25'b00001011_10001110_10011001_0;
      patterns[2961] = 25'b00001011_10001111_10011010_0;
      patterns[2962] = 25'b00001011_10010000_10011011_0;
      patterns[2963] = 25'b00001011_10010001_10011100_0;
      patterns[2964] = 25'b00001011_10010010_10011101_0;
      patterns[2965] = 25'b00001011_10010011_10011110_0;
      patterns[2966] = 25'b00001011_10010100_10011111_0;
      patterns[2967] = 25'b00001011_10010101_10100000_0;
      patterns[2968] = 25'b00001011_10010110_10100001_0;
      patterns[2969] = 25'b00001011_10010111_10100010_0;
      patterns[2970] = 25'b00001011_10011000_10100011_0;
      patterns[2971] = 25'b00001011_10011001_10100100_0;
      patterns[2972] = 25'b00001011_10011010_10100101_0;
      patterns[2973] = 25'b00001011_10011011_10100110_0;
      patterns[2974] = 25'b00001011_10011100_10100111_0;
      patterns[2975] = 25'b00001011_10011101_10101000_0;
      patterns[2976] = 25'b00001011_10011110_10101001_0;
      patterns[2977] = 25'b00001011_10011111_10101010_0;
      patterns[2978] = 25'b00001011_10100000_10101011_0;
      patterns[2979] = 25'b00001011_10100001_10101100_0;
      patterns[2980] = 25'b00001011_10100010_10101101_0;
      patterns[2981] = 25'b00001011_10100011_10101110_0;
      patterns[2982] = 25'b00001011_10100100_10101111_0;
      patterns[2983] = 25'b00001011_10100101_10110000_0;
      patterns[2984] = 25'b00001011_10100110_10110001_0;
      patterns[2985] = 25'b00001011_10100111_10110010_0;
      patterns[2986] = 25'b00001011_10101000_10110011_0;
      patterns[2987] = 25'b00001011_10101001_10110100_0;
      patterns[2988] = 25'b00001011_10101010_10110101_0;
      patterns[2989] = 25'b00001011_10101011_10110110_0;
      patterns[2990] = 25'b00001011_10101100_10110111_0;
      patterns[2991] = 25'b00001011_10101101_10111000_0;
      patterns[2992] = 25'b00001011_10101110_10111001_0;
      patterns[2993] = 25'b00001011_10101111_10111010_0;
      patterns[2994] = 25'b00001011_10110000_10111011_0;
      patterns[2995] = 25'b00001011_10110001_10111100_0;
      patterns[2996] = 25'b00001011_10110010_10111101_0;
      patterns[2997] = 25'b00001011_10110011_10111110_0;
      patterns[2998] = 25'b00001011_10110100_10111111_0;
      patterns[2999] = 25'b00001011_10110101_11000000_0;
      patterns[3000] = 25'b00001011_10110110_11000001_0;
      patterns[3001] = 25'b00001011_10110111_11000010_0;
      patterns[3002] = 25'b00001011_10111000_11000011_0;
      patterns[3003] = 25'b00001011_10111001_11000100_0;
      patterns[3004] = 25'b00001011_10111010_11000101_0;
      patterns[3005] = 25'b00001011_10111011_11000110_0;
      patterns[3006] = 25'b00001011_10111100_11000111_0;
      patterns[3007] = 25'b00001011_10111101_11001000_0;
      patterns[3008] = 25'b00001011_10111110_11001001_0;
      patterns[3009] = 25'b00001011_10111111_11001010_0;
      patterns[3010] = 25'b00001011_11000000_11001011_0;
      patterns[3011] = 25'b00001011_11000001_11001100_0;
      patterns[3012] = 25'b00001011_11000010_11001101_0;
      patterns[3013] = 25'b00001011_11000011_11001110_0;
      patterns[3014] = 25'b00001011_11000100_11001111_0;
      patterns[3015] = 25'b00001011_11000101_11010000_0;
      patterns[3016] = 25'b00001011_11000110_11010001_0;
      patterns[3017] = 25'b00001011_11000111_11010010_0;
      patterns[3018] = 25'b00001011_11001000_11010011_0;
      patterns[3019] = 25'b00001011_11001001_11010100_0;
      patterns[3020] = 25'b00001011_11001010_11010101_0;
      patterns[3021] = 25'b00001011_11001011_11010110_0;
      patterns[3022] = 25'b00001011_11001100_11010111_0;
      patterns[3023] = 25'b00001011_11001101_11011000_0;
      patterns[3024] = 25'b00001011_11001110_11011001_0;
      patterns[3025] = 25'b00001011_11001111_11011010_0;
      patterns[3026] = 25'b00001011_11010000_11011011_0;
      patterns[3027] = 25'b00001011_11010001_11011100_0;
      patterns[3028] = 25'b00001011_11010010_11011101_0;
      patterns[3029] = 25'b00001011_11010011_11011110_0;
      patterns[3030] = 25'b00001011_11010100_11011111_0;
      patterns[3031] = 25'b00001011_11010101_11100000_0;
      patterns[3032] = 25'b00001011_11010110_11100001_0;
      patterns[3033] = 25'b00001011_11010111_11100010_0;
      patterns[3034] = 25'b00001011_11011000_11100011_0;
      patterns[3035] = 25'b00001011_11011001_11100100_0;
      patterns[3036] = 25'b00001011_11011010_11100101_0;
      patterns[3037] = 25'b00001011_11011011_11100110_0;
      patterns[3038] = 25'b00001011_11011100_11100111_0;
      patterns[3039] = 25'b00001011_11011101_11101000_0;
      patterns[3040] = 25'b00001011_11011110_11101001_0;
      patterns[3041] = 25'b00001011_11011111_11101010_0;
      patterns[3042] = 25'b00001011_11100000_11101011_0;
      patterns[3043] = 25'b00001011_11100001_11101100_0;
      patterns[3044] = 25'b00001011_11100010_11101101_0;
      patterns[3045] = 25'b00001011_11100011_11101110_0;
      patterns[3046] = 25'b00001011_11100100_11101111_0;
      patterns[3047] = 25'b00001011_11100101_11110000_0;
      patterns[3048] = 25'b00001011_11100110_11110001_0;
      patterns[3049] = 25'b00001011_11100111_11110010_0;
      patterns[3050] = 25'b00001011_11101000_11110011_0;
      patterns[3051] = 25'b00001011_11101001_11110100_0;
      patterns[3052] = 25'b00001011_11101010_11110101_0;
      patterns[3053] = 25'b00001011_11101011_11110110_0;
      patterns[3054] = 25'b00001011_11101100_11110111_0;
      patterns[3055] = 25'b00001011_11101101_11111000_0;
      patterns[3056] = 25'b00001011_11101110_11111001_0;
      patterns[3057] = 25'b00001011_11101111_11111010_0;
      patterns[3058] = 25'b00001011_11110000_11111011_0;
      patterns[3059] = 25'b00001011_11110001_11111100_0;
      patterns[3060] = 25'b00001011_11110010_11111101_0;
      patterns[3061] = 25'b00001011_11110011_11111110_0;
      patterns[3062] = 25'b00001011_11110100_11111111_0;
      patterns[3063] = 25'b00001011_11110101_00000000_1;
      patterns[3064] = 25'b00001011_11110110_00000001_1;
      patterns[3065] = 25'b00001011_11110111_00000010_1;
      patterns[3066] = 25'b00001011_11111000_00000011_1;
      patterns[3067] = 25'b00001011_11111001_00000100_1;
      patterns[3068] = 25'b00001011_11111010_00000101_1;
      patterns[3069] = 25'b00001011_11111011_00000110_1;
      patterns[3070] = 25'b00001011_11111100_00000111_1;
      patterns[3071] = 25'b00001011_11111101_00001000_1;
      patterns[3072] = 25'b00001011_11111110_00001001_1;
      patterns[3073] = 25'b00001011_11111111_00001010_1;
      patterns[3074] = 25'b00001100_00000000_00001100_0;
      patterns[3075] = 25'b00001100_00000001_00001101_0;
      patterns[3076] = 25'b00001100_00000010_00001110_0;
      patterns[3077] = 25'b00001100_00000011_00001111_0;
      patterns[3078] = 25'b00001100_00000100_00010000_0;
      patterns[3079] = 25'b00001100_00000101_00010001_0;
      patterns[3080] = 25'b00001100_00000110_00010010_0;
      patterns[3081] = 25'b00001100_00000111_00010011_0;
      patterns[3082] = 25'b00001100_00001000_00010100_0;
      patterns[3083] = 25'b00001100_00001001_00010101_0;
      patterns[3084] = 25'b00001100_00001010_00010110_0;
      patterns[3085] = 25'b00001100_00001011_00010111_0;
      patterns[3086] = 25'b00001100_00001100_00011000_0;
      patterns[3087] = 25'b00001100_00001101_00011001_0;
      patterns[3088] = 25'b00001100_00001110_00011010_0;
      patterns[3089] = 25'b00001100_00001111_00011011_0;
      patterns[3090] = 25'b00001100_00010000_00011100_0;
      patterns[3091] = 25'b00001100_00010001_00011101_0;
      patterns[3092] = 25'b00001100_00010010_00011110_0;
      patterns[3093] = 25'b00001100_00010011_00011111_0;
      patterns[3094] = 25'b00001100_00010100_00100000_0;
      patterns[3095] = 25'b00001100_00010101_00100001_0;
      patterns[3096] = 25'b00001100_00010110_00100010_0;
      patterns[3097] = 25'b00001100_00010111_00100011_0;
      patterns[3098] = 25'b00001100_00011000_00100100_0;
      patterns[3099] = 25'b00001100_00011001_00100101_0;
      patterns[3100] = 25'b00001100_00011010_00100110_0;
      patterns[3101] = 25'b00001100_00011011_00100111_0;
      patterns[3102] = 25'b00001100_00011100_00101000_0;
      patterns[3103] = 25'b00001100_00011101_00101001_0;
      patterns[3104] = 25'b00001100_00011110_00101010_0;
      patterns[3105] = 25'b00001100_00011111_00101011_0;
      patterns[3106] = 25'b00001100_00100000_00101100_0;
      patterns[3107] = 25'b00001100_00100001_00101101_0;
      patterns[3108] = 25'b00001100_00100010_00101110_0;
      patterns[3109] = 25'b00001100_00100011_00101111_0;
      patterns[3110] = 25'b00001100_00100100_00110000_0;
      patterns[3111] = 25'b00001100_00100101_00110001_0;
      patterns[3112] = 25'b00001100_00100110_00110010_0;
      patterns[3113] = 25'b00001100_00100111_00110011_0;
      patterns[3114] = 25'b00001100_00101000_00110100_0;
      patterns[3115] = 25'b00001100_00101001_00110101_0;
      patterns[3116] = 25'b00001100_00101010_00110110_0;
      patterns[3117] = 25'b00001100_00101011_00110111_0;
      patterns[3118] = 25'b00001100_00101100_00111000_0;
      patterns[3119] = 25'b00001100_00101101_00111001_0;
      patterns[3120] = 25'b00001100_00101110_00111010_0;
      patterns[3121] = 25'b00001100_00101111_00111011_0;
      patterns[3122] = 25'b00001100_00110000_00111100_0;
      patterns[3123] = 25'b00001100_00110001_00111101_0;
      patterns[3124] = 25'b00001100_00110010_00111110_0;
      patterns[3125] = 25'b00001100_00110011_00111111_0;
      patterns[3126] = 25'b00001100_00110100_01000000_0;
      patterns[3127] = 25'b00001100_00110101_01000001_0;
      patterns[3128] = 25'b00001100_00110110_01000010_0;
      patterns[3129] = 25'b00001100_00110111_01000011_0;
      patterns[3130] = 25'b00001100_00111000_01000100_0;
      patterns[3131] = 25'b00001100_00111001_01000101_0;
      patterns[3132] = 25'b00001100_00111010_01000110_0;
      patterns[3133] = 25'b00001100_00111011_01000111_0;
      patterns[3134] = 25'b00001100_00111100_01001000_0;
      patterns[3135] = 25'b00001100_00111101_01001001_0;
      patterns[3136] = 25'b00001100_00111110_01001010_0;
      patterns[3137] = 25'b00001100_00111111_01001011_0;
      patterns[3138] = 25'b00001100_01000000_01001100_0;
      patterns[3139] = 25'b00001100_01000001_01001101_0;
      patterns[3140] = 25'b00001100_01000010_01001110_0;
      patterns[3141] = 25'b00001100_01000011_01001111_0;
      patterns[3142] = 25'b00001100_01000100_01010000_0;
      patterns[3143] = 25'b00001100_01000101_01010001_0;
      patterns[3144] = 25'b00001100_01000110_01010010_0;
      patterns[3145] = 25'b00001100_01000111_01010011_0;
      patterns[3146] = 25'b00001100_01001000_01010100_0;
      patterns[3147] = 25'b00001100_01001001_01010101_0;
      patterns[3148] = 25'b00001100_01001010_01010110_0;
      patterns[3149] = 25'b00001100_01001011_01010111_0;
      patterns[3150] = 25'b00001100_01001100_01011000_0;
      patterns[3151] = 25'b00001100_01001101_01011001_0;
      patterns[3152] = 25'b00001100_01001110_01011010_0;
      patterns[3153] = 25'b00001100_01001111_01011011_0;
      patterns[3154] = 25'b00001100_01010000_01011100_0;
      patterns[3155] = 25'b00001100_01010001_01011101_0;
      patterns[3156] = 25'b00001100_01010010_01011110_0;
      patterns[3157] = 25'b00001100_01010011_01011111_0;
      patterns[3158] = 25'b00001100_01010100_01100000_0;
      patterns[3159] = 25'b00001100_01010101_01100001_0;
      patterns[3160] = 25'b00001100_01010110_01100010_0;
      patterns[3161] = 25'b00001100_01010111_01100011_0;
      patterns[3162] = 25'b00001100_01011000_01100100_0;
      patterns[3163] = 25'b00001100_01011001_01100101_0;
      patterns[3164] = 25'b00001100_01011010_01100110_0;
      patterns[3165] = 25'b00001100_01011011_01100111_0;
      patterns[3166] = 25'b00001100_01011100_01101000_0;
      patterns[3167] = 25'b00001100_01011101_01101001_0;
      patterns[3168] = 25'b00001100_01011110_01101010_0;
      patterns[3169] = 25'b00001100_01011111_01101011_0;
      patterns[3170] = 25'b00001100_01100000_01101100_0;
      patterns[3171] = 25'b00001100_01100001_01101101_0;
      patterns[3172] = 25'b00001100_01100010_01101110_0;
      patterns[3173] = 25'b00001100_01100011_01101111_0;
      patterns[3174] = 25'b00001100_01100100_01110000_0;
      patterns[3175] = 25'b00001100_01100101_01110001_0;
      patterns[3176] = 25'b00001100_01100110_01110010_0;
      patterns[3177] = 25'b00001100_01100111_01110011_0;
      patterns[3178] = 25'b00001100_01101000_01110100_0;
      patterns[3179] = 25'b00001100_01101001_01110101_0;
      patterns[3180] = 25'b00001100_01101010_01110110_0;
      patterns[3181] = 25'b00001100_01101011_01110111_0;
      patterns[3182] = 25'b00001100_01101100_01111000_0;
      patterns[3183] = 25'b00001100_01101101_01111001_0;
      patterns[3184] = 25'b00001100_01101110_01111010_0;
      patterns[3185] = 25'b00001100_01101111_01111011_0;
      patterns[3186] = 25'b00001100_01110000_01111100_0;
      patterns[3187] = 25'b00001100_01110001_01111101_0;
      patterns[3188] = 25'b00001100_01110010_01111110_0;
      patterns[3189] = 25'b00001100_01110011_01111111_0;
      patterns[3190] = 25'b00001100_01110100_10000000_0;
      patterns[3191] = 25'b00001100_01110101_10000001_0;
      patterns[3192] = 25'b00001100_01110110_10000010_0;
      patterns[3193] = 25'b00001100_01110111_10000011_0;
      patterns[3194] = 25'b00001100_01111000_10000100_0;
      patterns[3195] = 25'b00001100_01111001_10000101_0;
      patterns[3196] = 25'b00001100_01111010_10000110_0;
      patterns[3197] = 25'b00001100_01111011_10000111_0;
      patterns[3198] = 25'b00001100_01111100_10001000_0;
      patterns[3199] = 25'b00001100_01111101_10001001_0;
      patterns[3200] = 25'b00001100_01111110_10001010_0;
      patterns[3201] = 25'b00001100_01111111_10001011_0;
      patterns[3202] = 25'b00001100_10000000_10001100_0;
      patterns[3203] = 25'b00001100_10000001_10001101_0;
      patterns[3204] = 25'b00001100_10000010_10001110_0;
      patterns[3205] = 25'b00001100_10000011_10001111_0;
      patterns[3206] = 25'b00001100_10000100_10010000_0;
      patterns[3207] = 25'b00001100_10000101_10010001_0;
      patterns[3208] = 25'b00001100_10000110_10010010_0;
      patterns[3209] = 25'b00001100_10000111_10010011_0;
      patterns[3210] = 25'b00001100_10001000_10010100_0;
      patterns[3211] = 25'b00001100_10001001_10010101_0;
      patterns[3212] = 25'b00001100_10001010_10010110_0;
      patterns[3213] = 25'b00001100_10001011_10010111_0;
      patterns[3214] = 25'b00001100_10001100_10011000_0;
      patterns[3215] = 25'b00001100_10001101_10011001_0;
      patterns[3216] = 25'b00001100_10001110_10011010_0;
      patterns[3217] = 25'b00001100_10001111_10011011_0;
      patterns[3218] = 25'b00001100_10010000_10011100_0;
      patterns[3219] = 25'b00001100_10010001_10011101_0;
      patterns[3220] = 25'b00001100_10010010_10011110_0;
      patterns[3221] = 25'b00001100_10010011_10011111_0;
      patterns[3222] = 25'b00001100_10010100_10100000_0;
      patterns[3223] = 25'b00001100_10010101_10100001_0;
      patterns[3224] = 25'b00001100_10010110_10100010_0;
      patterns[3225] = 25'b00001100_10010111_10100011_0;
      patterns[3226] = 25'b00001100_10011000_10100100_0;
      patterns[3227] = 25'b00001100_10011001_10100101_0;
      patterns[3228] = 25'b00001100_10011010_10100110_0;
      patterns[3229] = 25'b00001100_10011011_10100111_0;
      patterns[3230] = 25'b00001100_10011100_10101000_0;
      patterns[3231] = 25'b00001100_10011101_10101001_0;
      patterns[3232] = 25'b00001100_10011110_10101010_0;
      patterns[3233] = 25'b00001100_10011111_10101011_0;
      patterns[3234] = 25'b00001100_10100000_10101100_0;
      patterns[3235] = 25'b00001100_10100001_10101101_0;
      patterns[3236] = 25'b00001100_10100010_10101110_0;
      patterns[3237] = 25'b00001100_10100011_10101111_0;
      patterns[3238] = 25'b00001100_10100100_10110000_0;
      patterns[3239] = 25'b00001100_10100101_10110001_0;
      patterns[3240] = 25'b00001100_10100110_10110010_0;
      patterns[3241] = 25'b00001100_10100111_10110011_0;
      patterns[3242] = 25'b00001100_10101000_10110100_0;
      patterns[3243] = 25'b00001100_10101001_10110101_0;
      patterns[3244] = 25'b00001100_10101010_10110110_0;
      patterns[3245] = 25'b00001100_10101011_10110111_0;
      patterns[3246] = 25'b00001100_10101100_10111000_0;
      patterns[3247] = 25'b00001100_10101101_10111001_0;
      patterns[3248] = 25'b00001100_10101110_10111010_0;
      patterns[3249] = 25'b00001100_10101111_10111011_0;
      patterns[3250] = 25'b00001100_10110000_10111100_0;
      patterns[3251] = 25'b00001100_10110001_10111101_0;
      patterns[3252] = 25'b00001100_10110010_10111110_0;
      patterns[3253] = 25'b00001100_10110011_10111111_0;
      patterns[3254] = 25'b00001100_10110100_11000000_0;
      patterns[3255] = 25'b00001100_10110101_11000001_0;
      patterns[3256] = 25'b00001100_10110110_11000010_0;
      patterns[3257] = 25'b00001100_10110111_11000011_0;
      patterns[3258] = 25'b00001100_10111000_11000100_0;
      patterns[3259] = 25'b00001100_10111001_11000101_0;
      patterns[3260] = 25'b00001100_10111010_11000110_0;
      patterns[3261] = 25'b00001100_10111011_11000111_0;
      patterns[3262] = 25'b00001100_10111100_11001000_0;
      patterns[3263] = 25'b00001100_10111101_11001001_0;
      patterns[3264] = 25'b00001100_10111110_11001010_0;
      patterns[3265] = 25'b00001100_10111111_11001011_0;
      patterns[3266] = 25'b00001100_11000000_11001100_0;
      patterns[3267] = 25'b00001100_11000001_11001101_0;
      patterns[3268] = 25'b00001100_11000010_11001110_0;
      patterns[3269] = 25'b00001100_11000011_11001111_0;
      patterns[3270] = 25'b00001100_11000100_11010000_0;
      patterns[3271] = 25'b00001100_11000101_11010001_0;
      patterns[3272] = 25'b00001100_11000110_11010010_0;
      patterns[3273] = 25'b00001100_11000111_11010011_0;
      patterns[3274] = 25'b00001100_11001000_11010100_0;
      patterns[3275] = 25'b00001100_11001001_11010101_0;
      patterns[3276] = 25'b00001100_11001010_11010110_0;
      patterns[3277] = 25'b00001100_11001011_11010111_0;
      patterns[3278] = 25'b00001100_11001100_11011000_0;
      patterns[3279] = 25'b00001100_11001101_11011001_0;
      patterns[3280] = 25'b00001100_11001110_11011010_0;
      patterns[3281] = 25'b00001100_11001111_11011011_0;
      patterns[3282] = 25'b00001100_11010000_11011100_0;
      patterns[3283] = 25'b00001100_11010001_11011101_0;
      patterns[3284] = 25'b00001100_11010010_11011110_0;
      patterns[3285] = 25'b00001100_11010011_11011111_0;
      patterns[3286] = 25'b00001100_11010100_11100000_0;
      patterns[3287] = 25'b00001100_11010101_11100001_0;
      patterns[3288] = 25'b00001100_11010110_11100010_0;
      patterns[3289] = 25'b00001100_11010111_11100011_0;
      patterns[3290] = 25'b00001100_11011000_11100100_0;
      patterns[3291] = 25'b00001100_11011001_11100101_0;
      patterns[3292] = 25'b00001100_11011010_11100110_0;
      patterns[3293] = 25'b00001100_11011011_11100111_0;
      patterns[3294] = 25'b00001100_11011100_11101000_0;
      patterns[3295] = 25'b00001100_11011101_11101001_0;
      patterns[3296] = 25'b00001100_11011110_11101010_0;
      patterns[3297] = 25'b00001100_11011111_11101011_0;
      patterns[3298] = 25'b00001100_11100000_11101100_0;
      patterns[3299] = 25'b00001100_11100001_11101101_0;
      patterns[3300] = 25'b00001100_11100010_11101110_0;
      patterns[3301] = 25'b00001100_11100011_11101111_0;
      patterns[3302] = 25'b00001100_11100100_11110000_0;
      patterns[3303] = 25'b00001100_11100101_11110001_0;
      patterns[3304] = 25'b00001100_11100110_11110010_0;
      patterns[3305] = 25'b00001100_11100111_11110011_0;
      patterns[3306] = 25'b00001100_11101000_11110100_0;
      patterns[3307] = 25'b00001100_11101001_11110101_0;
      patterns[3308] = 25'b00001100_11101010_11110110_0;
      patterns[3309] = 25'b00001100_11101011_11110111_0;
      patterns[3310] = 25'b00001100_11101100_11111000_0;
      patterns[3311] = 25'b00001100_11101101_11111001_0;
      patterns[3312] = 25'b00001100_11101110_11111010_0;
      patterns[3313] = 25'b00001100_11101111_11111011_0;
      patterns[3314] = 25'b00001100_11110000_11111100_0;
      patterns[3315] = 25'b00001100_11110001_11111101_0;
      patterns[3316] = 25'b00001100_11110010_11111110_0;
      patterns[3317] = 25'b00001100_11110011_11111111_0;
      patterns[3318] = 25'b00001100_11110100_00000000_1;
      patterns[3319] = 25'b00001100_11110101_00000001_1;
      patterns[3320] = 25'b00001100_11110110_00000010_1;
      patterns[3321] = 25'b00001100_11110111_00000011_1;
      patterns[3322] = 25'b00001100_11111000_00000100_1;
      patterns[3323] = 25'b00001100_11111001_00000101_1;
      patterns[3324] = 25'b00001100_11111010_00000110_1;
      patterns[3325] = 25'b00001100_11111011_00000111_1;
      patterns[3326] = 25'b00001100_11111100_00001000_1;
      patterns[3327] = 25'b00001100_11111101_00001001_1;
      patterns[3328] = 25'b00001100_11111110_00001010_1;
      patterns[3329] = 25'b00001100_11111111_00001011_1;
      patterns[3330] = 25'b00001101_00000000_00001101_0;
      patterns[3331] = 25'b00001101_00000001_00001110_0;
      patterns[3332] = 25'b00001101_00000010_00001111_0;
      patterns[3333] = 25'b00001101_00000011_00010000_0;
      patterns[3334] = 25'b00001101_00000100_00010001_0;
      patterns[3335] = 25'b00001101_00000101_00010010_0;
      patterns[3336] = 25'b00001101_00000110_00010011_0;
      patterns[3337] = 25'b00001101_00000111_00010100_0;
      patterns[3338] = 25'b00001101_00001000_00010101_0;
      patterns[3339] = 25'b00001101_00001001_00010110_0;
      patterns[3340] = 25'b00001101_00001010_00010111_0;
      patterns[3341] = 25'b00001101_00001011_00011000_0;
      patterns[3342] = 25'b00001101_00001100_00011001_0;
      patterns[3343] = 25'b00001101_00001101_00011010_0;
      patterns[3344] = 25'b00001101_00001110_00011011_0;
      patterns[3345] = 25'b00001101_00001111_00011100_0;
      patterns[3346] = 25'b00001101_00010000_00011101_0;
      patterns[3347] = 25'b00001101_00010001_00011110_0;
      patterns[3348] = 25'b00001101_00010010_00011111_0;
      patterns[3349] = 25'b00001101_00010011_00100000_0;
      patterns[3350] = 25'b00001101_00010100_00100001_0;
      patterns[3351] = 25'b00001101_00010101_00100010_0;
      patterns[3352] = 25'b00001101_00010110_00100011_0;
      patterns[3353] = 25'b00001101_00010111_00100100_0;
      patterns[3354] = 25'b00001101_00011000_00100101_0;
      patterns[3355] = 25'b00001101_00011001_00100110_0;
      patterns[3356] = 25'b00001101_00011010_00100111_0;
      patterns[3357] = 25'b00001101_00011011_00101000_0;
      patterns[3358] = 25'b00001101_00011100_00101001_0;
      patterns[3359] = 25'b00001101_00011101_00101010_0;
      patterns[3360] = 25'b00001101_00011110_00101011_0;
      patterns[3361] = 25'b00001101_00011111_00101100_0;
      patterns[3362] = 25'b00001101_00100000_00101101_0;
      patterns[3363] = 25'b00001101_00100001_00101110_0;
      patterns[3364] = 25'b00001101_00100010_00101111_0;
      patterns[3365] = 25'b00001101_00100011_00110000_0;
      patterns[3366] = 25'b00001101_00100100_00110001_0;
      patterns[3367] = 25'b00001101_00100101_00110010_0;
      patterns[3368] = 25'b00001101_00100110_00110011_0;
      patterns[3369] = 25'b00001101_00100111_00110100_0;
      patterns[3370] = 25'b00001101_00101000_00110101_0;
      patterns[3371] = 25'b00001101_00101001_00110110_0;
      patterns[3372] = 25'b00001101_00101010_00110111_0;
      patterns[3373] = 25'b00001101_00101011_00111000_0;
      patterns[3374] = 25'b00001101_00101100_00111001_0;
      patterns[3375] = 25'b00001101_00101101_00111010_0;
      patterns[3376] = 25'b00001101_00101110_00111011_0;
      patterns[3377] = 25'b00001101_00101111_00111100_0;
      patterns[3378] = 25'b00001101_00110000_00111101_0;
      patterns[3379] = 25'b00001101_00110001_00111110_0;
      patterns[3380] = 25'b00001101_00110010_00111111_0;
      patterns[3381] = 25'b00001101_00110011_01000000_0;
      patterns[3382] = 25'b00001101_00110100_01000001_0;
      patterns[3383] = 25'b00001101_00110101_01000010_0;
      patterns[3384] = 25'b00001101_00110110_01000011_0;
      patterns[3385] = 25'b00001101_00110111_01000100_0;
      patterns[3386] = 25'b00001101_00111000_01000101_0;
      patterns[3387] = 25'b00001101_00111001_01000110_0;
      patterns[3388] = 25'b00001101_00111010_01000111_0;
      patterns[3389] = 25'b00001101_00111011_01001000_0;
      patterns[3390] = 25'b00001101_00111100_01001001_0;
      patterns[3391] = 25'b00001101_00111101_01001010_0;
      patterns[3392] = 25'b00001101_00111110_01001011_0;
      patterns[3393] = 25'b00001101_00111111_01001100_0;
      patterns[3394] = 25'b00001101_01000000_01001101_0;
      patterns[3395] = 25'b00001101_01000001_01001110_0;
      patterns[3396] = 25'b00001101_01000010_01001111_0;
      patterns[3397] = 25'b00001101_01000011_01010000_0;
      patterns[3398] = 25'b00001101_01000100_01010001_0;
      patterns[3399] = 25'b00001101_01000101_01010010_0;
      patterns[3400] = 25'b00001101_01000110_01010011_0;
      patterns[3401] = 25'b00001101_01000111_01010100_0;
      patterns[3402] = 25'b00001101_01001000_01010101_0;
      patterns[3403] = 25'b00001101_01001001_01010110_0;
      patterns[3404] = 25'b00001101_01001010_01010111_0;
      patterns[3405] = 25'b00001101_01001011_01011000_0;
      patterns[3406] = 25'b00001101_01001100_01011001_0;
      patterns[3407] = 25'b00001101_01001101_01011010_0;
      patterns[3408] = 25'b00001101_01001110_01011011_0;
      patterns[3409] = 25'b00001101_01001111_01011100_0;
      patterns[3410] = 25'b00001101_01010000_01011101_0;
      patterns[3411] = 25'b00001101_01010001_01011110_0;
      patterns[3412] = 25'b00001101_01010010_01011111_0;
      patterns[3413] = 25'b00001101_01010011_01100000_0;
      patterns[3414] = 25'b00001101_01010100_01100001_0;
      patterns[3415] = 25'b00001101_01010101_01100010_0;
      patterns[3416] = 25'b00001101_01010110_01100011_0;
      patterns[3417] = 25'b00001101_01010111_01100100_0;
      patterns[3418] = 25'b00001101_01011000_01100101_0;
      patterns[3419] = 25'b00001101_01011001_01100110_0;
      patterns[3420] = 25'b00001101_01011010_01100111_0;
      patterns[3421] = 25'b00001101_01011011_01101000_0;
      patterns[3422] = 25'b00001101_01011100_01101001_0;
      patterns[3423] = 25'b00001101_01011101_01101010_0;
      patterns[3424] = 25'b00001101_01011110_01101011_0;
      patterns[3425] = 25'b00001101_01011111_01101100_0;
      patterns[3426] = 25'b00001101_01100000_01101101_0;
      patterns[3427] = 25'b00001101_01100001_01101110_0;
      patterns[3428] = 25'b00001101_01100010_01101111_0;
      patterns[3429] = 25'b00001101_01100011_01110000_0;
      patterns[3430] = 25'b00001101_01100100_01110001_0;
      patterns[3431] = 25'b00001101_01100101_01110010_0;
      patterns[3432] = 25'b00001101_01100110_01110011_0;
      patterns[3433] = 25'b00001101_01100111_01110100_0;
      patterns[3434] = 25'b00001101_01101000_01110101_0;
      patterns[3435] = 25'b00001101_01101001_01110110_0;
      patterns[3436] = 25'b00001101_01101010_01110111_0;
      patterns[3437] = 25'b00001101_01101011_01111000_0;
      patterns[3438] = 25'b00001101_01101100_01111001_0;
      patterns[3439] = 25'b00001101_01101101_01111010_0;
      patterns[3440] = 25'b00001101_01101110_01111011_0;
      patterns[3441] = 25'b00001101_01101111_01111100_0;
      patterns[3442] = 25'b00001101_01110000_01111101_0;
      patterns[3443] = 25'b00001101_01110001_01111110_0;
      patterns[3444] = 25'b00001101_01110010_01111111_0;
      patterns[3445] = 25'b00001101_01110011_10000000_0;
      patterns[3446] = 25'b00001101_01110100_10000001_0;
      patterns[3447] = 25'b00001101_01110101_10000010_0;
      patterns[3448] = 25'b00001101_01110110_10000011_0;
      patterns[3449] = 25'b00001101_01110111_10000100_0;
      patterns[3450] = 25'b00001101_01111000_10000101_0;
      patterns[3451] = 25'b00001101_01111001_10000110_0;
      patterns[3452] = 25'b00001101_01111010_10000111_0;
      patterns[3453] = 25'b00001101_01111011_10001000_0;
      patterns[3454] = 25'b00001101_01111100_10001001_0;
      patterns[3455] = 25'b00001101_01111101_10001010_0;
      patterns[3456] = 25'b00001101_01111110_10001011_0;
      patterns[3457] = 25'b00001101_01111111_10001100_0;
      patterns[3458] = 25'b00001101_10000000_10001101_0;
      patterns[3459] = 25'b00001101_10000001_10001110_0;
      patterns[3460] = 25'b00001101_10000010_10001111_0;
      patterns[3461] = 25'b00001101_10000011_10010000_0;
      patterns[3462] = 25'b00001101_10000100_10010001_0;
      patterns[3463] = 25'b00001101_10000101_10010010_0;
      patterns[3464] = 25'b00001101_10000110_10010011_0;
      patterns[3465] = 25'b00001101_10000111_10010100_0;
      patterns[3466] = 25'b00001101_10001000_10010101_0;
      patterns[3467] = 25'b00001101_10001001_10010110_0;
      patterns[3468] = 25'b00001101_10001010_10010111_0;
      patterns[3469] = 25'b00001101_10001011_10011000_0;
      patterns[3470] = 25'b00001101_10001100_10011001_0;
      patterns[3471] = 25'b00001101_10001101_10011010_0;
      patterns[3472] = 25'b00001101_10001110_10011011_0;
      patterns[3473] = 25'b00001101_10001111_10011100_0;
      patterns[3474] = 25'b00001101_10010000_10011101_0;
      patterns[3475] = 25'b00001101_10010001_10011110_0;
      patterns[3476] = 25'b00001101_10010010_10011111_0;
      patterns[3477] = 25'b00001101_10010011_10100000_0;
      patterns[3478] = 25'b00001101_10010100_10100001_0;
      patterns[3479] = 25'b00001101_10010101_10100010_0;
      patterns[3480] = 25'b00001101_10010110_10100011_0;
      patterns[3481] = 25'b00001101_10010111_10100100_0;
      patterns[3482] = 25'b00001101_10011000_10100101_0;
      patterns[3483] = 25'b00001101_10011001_10100110_0;
      patterns[3484] = 25'b00001101_10011010_10100111_0;
      patterns[3485] = 25'b00001101_10011011_10101000_0;
      patterns[3486] = 25'b00001101_10011100_10101001_0;
      patterns[3487] = 25'b00001101_10011101_10101010_0;
      patterns[3488] = 25'b00001101_10011110_10101011_0;
      patterns[3489] = 25'b00001101_10011111_10101100_0;
      patterns[3490] = 25'b00001101_10100000_10101101_0;
      patterns[3491] = 25'b00001101_10100001_10101110_0;
      patterns[3492] = 25'b00001101_10100010_10101111_0;
      patterns[3493] = 25'b00001101_10100011_10110000_0;
      patterns[3494] = 25'b00001101_10100100_10110001_0;
      patterns[3495] = 25'b00001101_10100101_10110010_0;
      patterns[3496] = 25'b00001101_10100110_10110011_0;
      patterns[3497] = 25'b00001101_10100111_10110100_0;
      patterns[3498] = 25'b00001101_10101000_10110101_0;
      patterns[3499] = 25'b00001101_10101001_10110110_0;
      patterns[3500] = 25'b00001101_10101010_10110111_0;
      patterns[3501] = 25'b00001101_10101011_10111000_0;
      patterns[3502] = 25'b00001101_10101100_10111001_0;
      patterns[3503] = 25'b00001101_10101101_10111010_0;
      patterns[3504] = 25'b00001101_10101110_10111011_0;
      patterns[3505] = 25'b00001101_10101111_10111100_0;
      patterns[3506] = 25'b00001101_10110000_10111101_0;
      patterns[3507] = 25'b00001101_10110001_10111110_0;
      patterns[3508] = 25'b00001101_10110010_10111111_0;
      patterns[3509] = 25'b00001101_10110011_11000000_0;
      patterns[3510] = 25'b00001101_10110100_11000001_0;
      patterns[3511] = 25'b00001101_10110101_11000010_0;
      patterns[3512] = 25'b00001101_10110110_11000011_0;
      patterns[3513] = 25'b00001101_10110111_11000100_0;
      patterns[3514] = 25'b00001101_10111000_11000101_0;
      patterns[3515] = 25'b00001101_10111001_11000110_0;
      patterns[3516] = 25'b00001101_10111010_11000111_0;
      patterns[3517] = 25'b00001101_10111011_11001000_0;
      patterns[3518] = 25'b00001101_10111100_11001001_0;
      patterns[3519] = 25'b00001101_10111101_11001010_0;
      patterns[3520] = 25'b00001101_10111110_11001011_0;
      patterns[3521] = 25'b00001101_10111111_11001100_0;
      patterns[3522] = 25'b00001101_11000000_11001101_0;
      patterns[3523] = 25'b00001101_11000001_11001110_0;
      patterns[3524] = 25'b00001101_11000010_11001111_0;
      patterns[3525] = 25'b00001101_11000011_11010000_0;
      patterns[3526] = 25'b00001101_11000100_11010001_0;
      patterns[3527] = 25'b00001101_11000101_11010010_0;
      patterns[3528] = 25'b00001101_11000110_11010011_0;
      patterns[3529] = 25'b00001101_11000111_11010100_0;
      patterns[3530] = 25'b00001101_11001000_11010101_0;
      patterns[3531] = 25'b00001101_11001001_11010110_0;
      patterns[3532] = 25'b00001101_11001010_11010111_0;
      patterns[3533] = 25'b00001101_11001011_11011000_0;
      patterns[3534] = 25'b00001101_11001100_11011001_0;
      patterns[3535] = 25'b00001101_11001101_11011010_0;
      patterns[3536] = 25'b00001101_11001110_11011011_0;
      patterns[3537] = 25'b00001101_11001111_11011100_0;
      patterns[3538] = 25'b00001101_11010000_11011101_0;
      patterns[3539] = 25'b00001101_11010001_11011110_0;
      patterns[3540] = 25'b00001101_11010010_11011111_0;
      patterns[3541] = 25'b00001101_11010011_11100000_0;
      patterns[3542] = 25'b00001101_11010100_11100001_0;
      patterns[3543] = 25'b00001101_11010101_11100010_0;
      patterns[3544] = 25'b00001101_11010110_11100011_0;
      patterns[3545] = 25'b00001101_11010111_11100100_0;
      patterns[3546] = 25'b00001101_11011000_11100101_0;
      patterns[3547] = 25'b00001101_11011001_11100110_0;
      patterns[3548] = 25'b00001101_11011010_11100111_0;
      patterns[3549] = 25'b00001101_11011011_11101000_0;
      patterns[3550] = 25'b00001101_11011100_11101001_0;
      patterns[3551] = 25'b00001101_11011101_11101010_0;
      patterns[3552] = 25'b00001101_11011110_11101011_0;
      patterns[3553] = 25'b00001101_11011111_11101100_0;
      patterns[3554] = 25'b00001101_11100000_11101101_0;
      patterns[3555] = 25'b00001101_11100001_11101110_0;
      patterns[3556] = 25'b00001101_11100010_11101111_0;
      patterns[3557] = 25'b00001101_11100011_11110000_0;
      patterns[3558] = 25'b00001101_11100100_11110001_0;
      patterns[3559] = 25'b00001101_11100101_11110010_0;
      patterns[3560] = 25'b00001101_11100110_11110011_0;
      patterns[3561] = 25'b00001101_11100111_11110100_0;
      patterns[3562] = 25'b00001101_11101000_11110101_0;
      patterns[3563] = 25'b00001101_11101001_11110110_0;
      patterns[3564] = 25'b00001101_11101010_11110111_0;
      patterns[3565] = 25'b00001101_11101011_11111000_0;
      patterns[3566] = 25'b00001101_11101100_11111001_0;
      patterns[3567] = 25'b00001101_11101101_11111010_0;
      patterns[3568] = 25'b00001101_11101110_11111011_0;
      patterns[3569] = 25'b00001101_11101111_11111100_0;
      patterns[3570] = 25'b00001101_11110000_11111101_0;
      patterns[3571] = 25'b00001101_11110001_11111110_0;
      patterns[3572] = 25'b00001101_11110010_11111111_0;
      patterns[3573] = 25'b00001101_11110011_00000000_1;
      patterns[3574] = 25'b00001101_11110100_00000001_1;
      patterns[3575] = 25'b00001101_11110101_00000010_1;
      patterns[3576] = 25'b00001101_11110110_00000011_1;
      patterns[3577] = 25'b00001101_11110111_00000100_1;
      patterns[3578] = 25'b00001101_11111000_00000101_1;
      patterns[3579] = 25'b00001101_11111001_00000110_1;
      patterns[3580] = 25'b00001101_11111010_00000111_1;
      patterns[3581] = 25'b00001101_11111011_00001000_1;
      patterns[3582] = 25'b00001101_11111100_00001001_1;
      patterns[3583] = 25'b00001101_11111101_00001010_1;
      patterns[3584] = 25'b00001101_11111110_00001011_1;
      patterns[3585] = 25'b00001101_11111111_00001100_1;
      patterns[3586] = 25'b00001110_00000000_00001110_0;
      patterns[3587] = 25'b00001110_00000001_00001111_0;
      patterns[3588] = 25'b00001110_00000010_00010000_0;
      patterns[3589] = 25'b00001110_00000011_00010001_0;
      patterns[3590] = 25'b00001110_00000100_00010010_0;
      patterns[3591] = 25'b00001110_00000101_00010011_0;
      patterns[3592] = 25'b00001110_00000110_00010100_0;
      patterns[3593] = 25'b00001110_00000111_00010101_0;
      patterns[3594] = 25'b00001110_00001000_00010110_0;
      patterns[3595] = 25'b00001110_00001001_00010111_0;
      patterns[3596] = 25'b00001110_00001010_00011000_0;
      patterns[3597] = 25'b00001110_00001011_00011001_0;
      patterns[3598] = 25'b00001110_00001100_00011010_0;
      patterns[3599] = 25'b00001110_00001101_00011011_0;
      patterns[3600] = 25'b00001110_00001110_00011100_0;
      patterns[3601] = 25'b00001110_00001111_00011101_0;
      patterns[3602] = 25'b00001110_00010000_00011110_0;
      patterns[3603] = 25'b00001110_00010001_00011111_0;
      patterns[3604] = 25'b00001110_00010010_00100000_0;
      patterns[3605] = 25'b00001110_00010011_00100001_0;
      patterns[3606] = 25'b00001110_00010100_00100010_0;
      patterns[3607] = 25'b00001110_00010101_00100011_0;
      patterns[3608] = 25'b00001110_00010110_00100100_0;
      patterns[3609] = 25'b00001110_00010111_00100101_0;
      patterns[3610] = 25'b00001110_00011000_00100110_0;
      patterns[3611] = 25'b00001110_00011001_00100111_0;
      patterns[3612] = 25'b00001110_00011010_00101000_0;
      patterns[3613] = 25'b00001110_00011011_00101001_0;
      patterns[3614] = 25'b00001110_00011100_00101010_0;
      patterns[3615] = 25'b00001110_00011101_00101011_0;
      patterns[3616] = 25'b00001110_00011110_00101100_0;
      patterns[3617] = 25'b00001110_00011111_00101101_0;
      patterns[3618] = 25'b00001110_00100000_00101110_0;
      patterns[3619] = 25'b00001110_00100001_00101111_0;
      patterns[3620] = 25'b00001110_00100010_00110000_0;
      patterns[3621] = 25'b00001110_00100011_00110001_0;
      patterns[3622] = 25'b00001110_00100100_00110010_0;
      patterns[3623] = 25'b00001110_00100101_00110011_0;
      patterns[3624] = 25'b00001110_00100110_00110100_0;
      patterns[3625] = 25'b00001110_00100111_00110101_0;
      patterns[3626] = 25'b00001110_00101000_00110110_0;
      patterns[3627] = 25'b00001110_00101001_00110111_0;
      patterns[3628] = 25'b00001110_00101010_00111000_0;
      patterns[3629] = 25'b00001110_00101011_00111001_0;
      patterns[3630] = 25'b00001110_00101100_00111010_0;
      patterns[3631] = 25'b00001110_00101101_00111011_0;
      patterns[3632] = 25'b00001110_00101110_00111100_0;
      patterns[3633] = 25'b00001110_00101111_00111101_0;
      patterns[3634] = 25'b00001110_00110000_00111110_0;
      patterns[3635] = 25'b00001110_00110001_00111111_0;
      patterns[3636] = 25'b00001110_00110010_01000000_0;
      patterns[3637] = 25'b00001110_00110011_01000001_0;
      patterns[3638] = 25'b00001110_00110100_01000010_0;
      patterns[3639] = 25'b00001110_00110101_01000011_0;
      patterns[3640] = 25'b00001110_00110110_01000100_0;
      patterns[3641] = 25'b00001110_00110111_01000101_0;
      patterns[3642] = 25'b00001110_00111000_01000110_0;
      patterns[3643] = 25'b00001110_00111001_01000111_0;
      patterns[3644] = 25'b00001110_00111010_01001000_0;
      patterns[3645] = 25'b00001110_00111011_01001001_0;
      patterns[3646] = 25'b00001110_00111100_01001010_0;
      patterns[3647] = 25'b00001110_00111101_01001011_0;
      patterns[3648] = 25'b00001110_00111110_01001100_0;
      patterns[3649] = 25'b00001110_00111111_01001101_0;
      patterns[3650] = 25'b00001110_01000000_01001110_0;
      patterns[3651] = 25'b00001110_01000001_01001111_0;
      patterns[3652] = 25'b00001110_01000010_01010000_0;
      patterns[3653] = 25'b00001110_01000011_01010001_0;
      patterns[3654] = 25'b00001110_01000100_01010010_0;
      patterns[3655] = 25'b00001110_01000101_01010011_0;
      patterns[3656] = 25'b00001110_01000110_01010100_0;
      patterns[3657] = 25'b00001110_01000111_01010101_0;
      patterns[3658] = 25'b00001110_01001000_01010110_0;
      patterns[3659] = 25'b00001110_01001001_01010111_0;
      patterns[3660] = 25'b00001110_01001010_01011000_0;
      patterns[3661] = 25'b00001110_01001011_01011001_0;
      patterns[3662] = 25'b00001110_01001100_01011010_0;
      patterns[3663] = 25'b00001110_01001101_01011011_0;
      patterns[3664] = 25'b00001110_01001110_01011100_0;
      patterns[3665] = 25'b00001110_01001111_01011101_0;
      patterns[3666] = 25'b00001110_01010000_01011110_0;
      patterns[3667] = 25'b00001110_01010001_01011111_0;
      patterns[3668] = 25'b00001110_01010010_01100000_0;
      patterns[3669] = 25'b00001110_01010011_01100001_0;
      patterns[3670] = 25'b00001110_01010100_01100010_0;
      patterns[3671] = 25'b00001110_01010101_01100011_0;
      patterns[3672] = 25'b00001110_01010110_01100100_0;
      patterns[3673] = 25'b00001110_01010111_01100101_0;
      patterns[3674] = 25'b00001110_01011000_01100110_0;
      patterns[3675] = 25'b00001110_01011001_01100111_0;
      patterns[3676] = 25'b00001110_01011010_01101000_0;
      patterns[3677] = 25'b00001110_01011011_01101001_0;
      patterns[3678] = 25'b00001110_01011100_01101010_0;
      patterns[3679] = 25'b00001110_01011101_01101011_0;
      patterns[3680] = 25'b00001110_01011110_01101100_0;
      patterns[3681] = 25'b00001110_01011111_01101101_0;
      patterns[3682] = 25'b00001110_01100000_01101110_0;
      patterns[3683] = 25'b00001110_01100001_01101111_0;
      patterns[3684] = 25'b00001110_01100010_01110000_0;
      patterns[3685] = 25'b00001110_01100011_01110001_0;
      patterns[3686] = 25'b00001110_01100100_01110010_0;
      patterns[3687] = 25'b00001110_01100101_01110011_0;
      patterns[3688] = 25'b00001110_01100110_01110100_0;
      patterns[3689] = 25'b00001110_01100111_01110101_0;
      patterns[3690] = 25'b00001110_01101000_01110110_0;
      patterns[3691] = 25'b00001110_01101001_01110111_0;
      patterns[3692] = 25'b00001110_01101010_01111000_0;
      patterns[3693] = 25'b00001110_01101011_01111001_0;
      patterns[3694] = 25'b00001110_01101100_01111010_0;
      patterns[3695] = 25'b00001110_01101101_01111011_0;
      patterns[3696] = 25'b00001110_01101110_01111100_0;
      patterns[3697] = 25'b00001110_01101111_01111101_0;
      patterns[3698] = 25'b00001110_01110000_01111110_0;
      patterns[3699] = 25'b00001110_01110001_01111111_0;
      patterns[3700] = 25'b00001110_01110010_10000000_0;
      patterns[3701] = 25'b00001110_01110011_10000001_0;
      patterns[3702] = 25'b00001110_01110100_10000010_0;
      patterns[3703] = 25'b00001110_01110101_10000011_0;
      patterns[3704] = 25'b00001110_01110110_10000100_0;
      patterns[3705] = 25'b00001110_01110111_10000101_0;
      patterns[3706] = 25'b00001110_01111000_10000110_0;
      patterns[3707] = 25'b00001110_01111001_10000111_0;
      patterns[3708] = 25'b00001110_01111010_10001000_0;
      patterns[3709] = 25'b00001110_01111011_10001001_0;
      patterns[3710] = 25'b00001110_01111100_10001010_0;
      patterns[3711] = 25'b00001110_01111101_10001011_0;
      patterns[3712] = 25'b00001110_01111110_10001100_0;
      patterns[3713] = 25'b00001110_01111111_10001101_0;
      patterns[3714] = 25'b00001110_10000000_10001110_0;
      patterns[3715] = 25'b00001110_10000001_10001111_0;
      patterns[3716] = 25'b00001110_10000010_10010000_0;
      patterns[3717] = 25'b00001110_10000011_10010001_0;
      patterns[3718] = 25'b00001110_10000100_10010010_0;
      patterns[3719] = 25'b00001110_10000101_10010011_0;
      patterns[3720] = 25'b00001110_10000110_10010100_0;
      patterns[3721] = 25'b00001110_10000111_10010101_0;
      patterns[3722] = 25'b00001110_10001000_10010110_0;
      patterns[3723] = 25'b00001110_10001001_10010111_0;
      patterns[3724] = 25'b00001110_10001010_10011000_0;
      patterns[3725] = 25'b00001110_10001011_10011001_0;
      patterns[3726] = 25'b00001110_10001100_10011010_0;
      patterns[3727] = 25'b00001110_10001101_10011011_0;
      patterns[3728] = 25'b00001110_10001110_10011100_0;
      patterns[3729] = 25'b00001110_10001111_10011101_0;
      patterns[3730] = 25'b00001110_10010000_10011110_0;
      patterns[3731] = 25'b00001110_10010001_10011111_0;
      patterns[3732] = 25'b00001110_10010010_10100000_0;
      patterns[3733] = 25'b00001110_10010011_10100001_0;
      patterns[3734] = 25'b00001110_10010100_10100010_0;
      patterns[3735] = 25'b00001110_10010101_10100011_0;
      patterns[3736] = 25'b00001110_10010110_10100100_0;
      patterns[3737] = 25'b00001110_10010111_10100101_0;
      patterns[3738] = 25'b00001110_10011000_10100110_0;
      patterns[3739] = 25'b00001110_10011001_10100111_0;
      patterns[3740] = 25'b00001110_10011010_10101000_0;
      patterns[3741] = 25'b00001110_10011011_10101001_0;
      patterns[3742] = 25'b00001110_10011100_10101010_0;
      patterns[3743] = 25'b00001110_10011101_10101011_0;
      patterns[3744] = 25'b00001110_10011110_10101100_0;
      patterns[3745] = 25'b00001110_10011111_10101101_0;
      patterns[3746] = 25'b00001110_10100000_10101110_0;
      patterns[3747] = 25'b00001110_10100001_10101111_0;
      patterns[3748] = 25'b00001110_10100010_10110000_0;
      patterns[3749] = 25'b00001110_10100011_10110001_0;
      patterns[3750] = 25'b00001110_10100100_10110010_0;
      patterns[3751] = 25'b00001110_10100101_10110011_0;
      patterns[3752] = 25'b00001110_10100110_10110100_0;
      patterns[3753] = 25'b00001110_10100111_10110101_0;
      patterns[3754] = 25'b00001110_10101000_10110110_0;
      patterns[3755] = 25'b00001110_10101001_10110111_0;
      patterns[3756] = 25'b00001110_10101010_10111000_0;
      patterns[3757] = 25'b00001110_10101011_10111001_0;
      patterns[3758] = 25'b00001110_10101100_10111010_0;
      patterns[3759] = 25'b00001110_10101101_10111011_0;
      patterns[3760] = 25'b00001110_10101110_10111100_0;
      patterns[3761] = 25'b00001110_10101111_10111101_0;
      patterns[3762] = 25'b00001110_10110000_10111110_0;
      patterns[3763] = 25'b00001110_10110001_10111111_0;
      patterns[3764] = 25'b00001110_10110010_11000000_0;
      patterns[3765] = 25'b00001110_10110011_11000001_0;
      patterns[3766] = 25'b00001110_10110100_11000010_0;
      patterns[3767] = 25'b00001110_10110101_11000011_0;
      patterns[3768] = 25'b00001110_10110110_11000100_0;
      patterns[3769] = 25'b00001110_10110111_11000101_0;
      patterns[3770] = 25'b00001110_10111000_11000110_0;
      patterns[3771] = 25'b00001110_10111001_11000111_0;
      patterns[3772] = 25'b00001110_10111010_11001000_0;
      patterns[3773] = 25'b00001110_10111011_11001001_0;
      patterns[3774] = 25'b00001110_10111100_11001010_0;
      patterns[3775] = 25'b00001110_10111101_11001011_0;
      patterns[3776] = 25'b00001110_10111110_11001100_0;
      patterns[3777] = 25'b00001110_10111111_11001101_0;
      patterns[3778] = 25'b00001110_11000000_11001110_0;
      patterns[3779] = 25'b00001110_11000001_11001111_0;
      patterns[3780] = 25'b00001110_11000010_11010000_0;
      patterns[3781] = 25'b00001110_11000011_11010001_0;
      patterns[3782] = 25'b00001110_11000100_11010010_0;
      patterns[3783] = 25'b00001110_11000101_11010011_0;
      patterns[3784] = 25'b00001110_11000110_11010100_0;
      patterns[3785] = 25'b00001110_11000111_11010101_0;
      patterns[3786] = 25'b00001110_11001000_11010110_0;
      patterns[3787] = 25'b00001110_11001001_11010111_0;
      patterns[3788] = 25'b00001110_11001010_11011000_0;
      patterns[3789] = 25'b00001110_11001011_11011001_0;
      patterns[3790] = 25'b00001110_11001100_11011010_0;
      patterns[3791] = 25'b00001110_11001101_11011011_0;
      patterns[3792] = 25'b00001110_11001110_11011100_0;
      patterns[3793] = 25'b00001110_11001111_11011101_0;
      patterns[3794] = 25'b00001110_11010000_11011110_0;
      patterns[3795] = 25'b00001110_11010001_11011111_0;
      patterns[3796] = 25'b00001110_11010010_11100000_0;
      patterns[3797] = 25'b00001110_11010011_11100001_0;
      patterns[3798] = 25'b00001110_11010100_11100010_0;
      patterns[3799] = 25'b00001110_11010101_11100011_0;
      patterns[3800] = 25'b00001110_11010110_11100100_0;
      patterns[3801] = 25'b00001110_11010111_11100101_0;
      patterns[3802] = 25'b00001110_11011000_11100110_0;
      patterns[3803] = 25'b00001110_11011001_11100111_0;
      patterns[3804] = 25'b00001110_11011010_11101000_0;
      patterns[3805] = 25'b00001110_11011011_11101001_0;
      patterns[3806] = 25'b00001110_11011100_11101010_0;
      patterns[3807] = 25'b00001110_11011101_11101011_0;
      patterns[3808] = 25'b00001110_11011110_11101100_0;
      patterns[3809] = 25'b00001110_11011111_11101101_0;
      patterns[3810] = 25'b00001110_11100000_11101110_0;
      patterns[3811] = 25'b00001110_11100001_11101111_0;
      patterns[3812] = 25'b00001110_11100010_11110000_0;
      patterns[3813] = 25'b00001110_11100011_11110001_0;
      patterns[3814] = 25'b00001110_11100100_11110010_0;
      patterns[3815] = 25'b00001110_11100101_11110011_0;
      patterns[3816] = 25'b00001110_11100110_11110100_0;
      patterns[3817] = 25'b00001110_11100111_11110101_0;
      patterns[3818] = 25'b00001110_11101000_11110110_0;
      patterns[3819] = 25'b00001110_11101001_11110111_0;
      patterns[3820] = 25'b00001110_11101010_11111000_0;
      patterns[3821] = 25'b00001110_11101011_11111001_0;
      patterns[3822] = 25'b00001110_11101100_11111010_0;
      patterns[3823] = 25'b00001110_11101101_11111011_0;
      patterns[3824] = 25'b00001110_11101110_11111100_0;
      patterns[3825] = 25'b00001110_11101111_11111101_0;
      patterns[3826] = 25'b00001110_11110000_11111110_0;
      patterns[3827] = 25'b00001110_11110001_11111111_0;
      patterns[3828] = 25'b00001110_11110010_00000000_1;
      patterns[3829] = 25'b00001110_11110011_00000001_1;
      patterns[3830] = 25'b00001110_11110100_00000010_1;
      patterns[3831] = 25'b00001110_11110101_00000011_1;
      patterns[3832] = 25'b00001110_11110110_00000100_1;
      patterns[3833] = 25'b00001110_11110111_00000101_1;
      patterns[3834] = 25'b00001110_11111000_00000110_1;
      patterns[3835] = 25'b00001110_11111001_00000111_1;
      patterns[3836] = 25'b00001110_11111010_00001000_1;
      patterns[3837] = 25'b00001110_11111011_00001001_1;
      patterns[3838] = 25'b00001110_11111100_00001010_1;
      patterns[3839] = 25'b00001110_11111101_00001011_1;
      patterns[3840] = 25'b00001110_11111110_00001100_1;
      patterns[3841] = 25'b00001110_11111111_00001101_1;
      patterns[3842] = 25'b00001111_00000000_00001111_0;
      patterns[3843] = 25'b00001111_00000001_00010000_0;
      patterns[3844] = 25'b00001111_00000010_00010001_0;
      patterns[3845] = 25'b00001111_00000011_00010010_0;
      patterns[3846] = 25'b00001111_00000100_00010011_0;
      patterns[3847] = 25'b00001111_00000101_00010100_0;
      patterns[3848] = 25'b00001111_00000110_00010101_0;
      patterns[3849] = 25'b00001111_00000111_00010110_0;
      patterns[3850] = 25'b00001111_00001000_00010111_0;
      patterns[3851] = 25'b00001111_00001001_00011000_0;
      patterns[3852] = 25'b00001111_00001010_00011001_0;
      patterns[3853] = 25'b00001111_00001011_00011010_0;
      patterns[3854] = 25'b00001111_00001100_00011011_0;
      patterns[3855] = 25'b00001111_00001101_00011100_0;
      patterns[3856] = 25'b00001111_00001110_00011101_0;
      patterns[3857] = 25'b00001111_00001111_00011110_0;
      patterns[3858] = 25'b00001111_00010000_00011111_0;
      patterns[3859] = 25'b00001111_00010001_00100000_0;
      patterns[3860] = 25'b00001111_00010010_00100001_0;
      patterns[3861] = 25'b00001111_00010011_00100010_0;
      patterns[3862] = 25'b00001111_00010100_00100011_0;
      patterns[3863] = 25'b00001111_00010101_00100100_0;
      patterns[3864] = 25'b00001111_00010110_00100101_0;
      patterns[3865] = 25'b00001111_00010111_00100110_0;
      patterns[3866] = 25'b00001111_00011000_00100111_0;
      patterns[3867] = 25'b00001111_00011001_00101000_0;
      patterns[3868] = 25'b00001111_00011010_00101001_0;
      patterns[3869] = 25'b00001111_00011011_00101010_0;
      patterns[3870] = 25'b00001111_00011100_00101011_0;
      patterns[3871] = 25'b00001111_00011101_00101100_0;
      patterns[3872] = 25'b00001111_00011110_00101101_0;
      patterns[3873] = 25'b00001111_00011111_00101110_0;
      patterns[3874] = 25'b00001111_00100000_00101111_0;
      patterns[3875] = 25'b00001111_00100001_00110000_0;
      patterns[3876] = 25'b00001111_00100010_00110001_0;
      patterns[3877] = 25'b00001111_00100011_00110010_0;
      patterns[3878] = 25'b00001111_00100100_00110011_0;
      patterns[3879] = 25'b00001111_00100101_00110100_0;
      patterns[3880] = 25'b00001111_00100110_00110101_0;
      patterns[3881] = 25'b00001111_00100111_00110110_0;
      patterns[3882] = 25'b00001111_00101000_00110111_0;
      patterns[3883] = 25'b00001111_00101001_00111000_0;
      patterns[3884] = 25'b00001111_00101010_00111001_0;
      patterns[3885] = 25'b00001111_00101011_00111010_0;
      patterns[3886] = 25'b00001111_00101100_00111011_0;
      patterns[3887] = 25'b00001111_00101101_00111100_0;
      patterns[3888] = 25'b00001111_00101110_00111101_0;
      patterns[3889] = 25'b00001111_00101111_00111110_0;
      patterns[3890] = 25'b00001111_00110000_00111111_0;
      patterns[3891] = 25'b00001111_00110001_01000000_0;
      patterns[3892] = 25'b00001111_00110010_01000001_0;
      patterns[3893] = 25'b00001111_00110011_01000010_0;
      patterns[3894] = 25'b00001111_00110100_01000011_0;
      patterns[3895] = 25'b00001111_00110101_01000100_0;
      patterns[3896] = 25'b00001111_00110110_01000101_0;
      patterns[3897] = 25'b00001111_00110111_01000110_0;
      patterns[3898] = 25'b00001111_00111000_01000111_0;
      patterns[3899] = 25'b00001111_00111001_01001000_0;
      patterns[3900] = 25'b00001111_00111010_01001001_0;
      patterns[3901] = 25'b00001111_00111011_01001010_0;
      patterns[3902] = 25'b00001111_00111100_01001011_0;
      patterns[3903] = 25'b00001111_00111101_01001100_0;
      patterns[3904] = 25'b00001111_00111110_01001101_0;
      patterns[3905] = 25'b00001111_00111111_01001110_0;
      patterns[3906] = 25'b00001111_01000000_01001111_0;
      patterns[3907] = 25'b00001111_01000001_01010000_0;
      patterns[3908] = 25'b00001111_01000010_01010001_0;
      patterns[3909] = 25'b00001111_01000011_01010010_0;
      patterns[3910] = 25'b00001111_01000100_01010011_0;
      patterns[3911] = 25'b00001111_01000101_01010100_0;
      patterns[3912] = 25'b00001111_01000110_01010101_0;
      patterns[3913] = 25'b00001111_01000111_01010110_0;
      patterns[3914] = 25'b00001111_01001000_01010111_0;
      patterns[3915] = 25'b00001111_01001001_01011000_0;
      patterns[3916] = 25'b00001111_01001010_01011001_0;
      patterns[3917] = 25'b00001111_01001011_01011010_0;
      patterns[3918] = 25'b00001111_01001100_01011011_0;
      patterns[3919] = 25'b00001111_01001101_01011100_0;
      patterns[3920] = 25'b00001111_01001110_01011101_0;
      patterns[3921] = 25'b00001111_01001111_01011110_0;
      patterns[3922] = 25'b00001111_01010000_01011111_0;
      patterns[3923] = 25'b00001111_01010001_01100000_0;
      patterns[3924] = 25'b00001111_01010010_01100001_0;
      patterns[3925] = 25'b00001111_01010011_01100010_0;
      patterns[3926] = 25'b00001111_01010100_01100011_0;
      patterns[3927] = 25'b00001111_01010101_01100100_0;
      patterns[3928] = 25'b00001111_01010110_01100101_0;
      patterns[3929] = 25'b00001111_01010111_01100110_0;
      patterns[3930] = 25'b00001111_01011000_01100111_0;
      patterns[3931] = 25'b00001111_01011001_01101000_0;
      patterns[3932] = 25'b00001111_01011010_01101001_0;
      patterns[3933] = 25'b00001111_01011011_01101010_0;
      patterns[3934] = 25'b00001111_01011100_01101011_0;
      patterns[3935] = 25'b00001111_01011101_01101100_0;
      patterns[3936] = 25'b00001111_01011110_01101101_0;
      patterns[3937] = 25'b00001111_01011111_01101110_0;
      patterns[3938] = 25'b00001111_01100000_01101111_0;
      patterns[3939] = 25'b00001111_01100001_01110000_0;
      patterns[3940] = 25'b00001111_01100010_01110001_0;
      patterns[3941] = 25'b00001111_01100011_01110010_0;
      patterns[3942] = 25'b00001111_01100100_01110011_0;
      patterns[3943] = 25'b00001111_01100101_01110100_0;
      patterns[3944] = 25'b00001111_01100110_01110101_0;
      patterns[3945] = 25'b00001111_01100111_01110110_0;
      patterns[3946] = 25'b00001111_01101000_01110111_0;
      patterns[3947] = 25'b00001111_01101001_01111000_0;
      patterns[3948] = 25'b00001111_01101010_01111001_0;
      patterns[3949] = 25'b00001111_01101011_01111010_0;
      patterns[3950] = 25'b00001111_01101100_01111011_0;
      patterns[3951] = 25'b00001111_01101101_01111100_0;
      patterns[3952] = 25'b00001111_01101110_01111101_0;
      patterns[3953] = 25'b00001111_01101111_01111110_0;
      patterns[3954] = 25'b00001111_01110000_01111111_0;
      patterns[3955] = 25'b00001111_01110001_10000000_0;
      patterns[3956] = 25'b00001111_01110010_10000001_0;
      patterns[3957] = 25'b00001111_01110011_10000010_0;
      patterns[3958] = 25'b00001111_01110100_10000011_0;
      patterns[3959] = 25'b00001111_01110101_10000100_0;
      patterns[3960] = 25'b00001111_01110110_10000101_0;
      patterns[3961] = 25'b00001111_01110111_10000110_0;
      patterns[3962] = 25'b00001111_01111000_10000111_0;
      patterns[3963] = 25'b00001111_01111001_10001000_0;
      patterns[3964] = 25'b00001111_01111010_10001001_0;
      patterns[3965] = 25'b00001111_01111011_10001010_0;
      patterns[3966] = 25'b00001111_01111100_10001011_0;
      patterns[3967] = 25'b00001111_01111101_10001100_0;
      patterns[3968] = 25'b00001111_01111110_10001101_0;
      patterns[3969] = 25'b00001111_01111111_10001110_0;
      patterns[3970] = 25'b00001111_10000000_10001111_0;
      patterns[3971] = 25'b00001111_10000001_10010000_0;
      patterns[3972] = 25'b00001111_10000010_10010001_0;
      patterns[3973] = 25'b00001111_10000011_10010010_0;
      patterns[3974] = 25'b00001111_10000100_10010011_0;
      patterns[3975] = 25'b00001111_10000101_10010100_0;
      patterns[3976] = 25'b00001111_10000110_10010101_0;
      patterns[3977] = 25'b00001111_10000111_10010110_0;
      patterns[3978] = 25'b00001111_10001000_10010111_0;
      patterns[3979] = 25'b00001111_10001001_10011000_0;
      patterns[3980] = 25'b00001111_10001010_10011001_0;
      patterns[3981] = 25'b00001111_10001011_10011010_0;
      patterns[3982] = 25'b00001111_10001100_10011011_0;
      patterns[3983] = 25'b00001111_10001101_10011100_0;
      patterns[3984] = 25'b00001111_10001110_10011101_0;
      patterns[3985] = 25'b00001111_10001111_10011110_0;
      patterns[3986] = 25'b00001111_10010000_10011111_0;
      patterns[3987] = 25'b00001111_10010001_10100000_0;
      patterns[3988] = 25'b00001111_10010010_10100001_0;
      patterns[3989] = 25'b00001111_10010011_10100010_0;
      patterns[3990] = 25'b00001111_10010100_10100011_0;
      patterns[3991] = 25'b00001111_10010101_10100100_0;
      patterns[3992] = 25'b00001111_10010110_10100101_0;
      patterns[3993] = 25'b00001111_10010111_10100110_0;
      patterns[3994] = 25'b00001111_10011000_10100111_0;
      patterns[3995] = 25'b00001111_10011001_10101000_0;
      patterns[3996] = 25'b00001111_10011010_10101001_0;
      patterns[3997] = 25'b00001111_10011011_10101010_0;
      patterns[3998] = 25'b00001111_10011100_10101011_0;
      patterns[3999] = 25'b00001111_10011101_10101100_0;
      patterns[4000] = 25'b00001111_10011110_10101101_0;
      patterns[4001] = 25'b00001111_10011111_10101110_0;
      patterns[4002] = 25'b00001111_10100000_10101111_0;
      patterns[4003] = 25'b00001111_10100001_10110000_0;
      patterns[4004] = 25'b00001111_10100010_10110001_0;
      patterns[4005] = 25'b00001111_10100011_10110010_0;
      patterns[4006] = 25'b00001111_10100100_10110011_0;
      patterns[4007] = 25'b00001111_10100101_10110100_0;
      patterns[4008] = 25'b00001111_10100110_10110101_0;
      patterns[4009] = 25'b00001111_10100111_10110110_0;
      patterns[4010] = 25'b00001111_10101000_10110111_0;
      patterns[4011] = 25'b00001111_10101001_10111000_0;
      patterns[4012] = 25'b00001111_10101010_10111001_0;
      patterns[4013] = 25'b00001111_10101011_10111010_0;
      patterns[4014] = 25'b00001111_10101100_10111011_0;
      patterns[4015] = 25'b00001111_10101101_10111100_0;
      patterns[4016] = 25'b00001111_10101110_10111101_0;
      patterns[4017] = 25'b00001111_10101111_10111110_0;
      patterns[4018] = 25'b00001111_10110000_10111111_0;
      patterns[4019] = 25'b00001111_10110001_11000000_0;
      patterns[4020] = 25'b00001111_10110010_11000001_0;
      patterns[4021] = 25'b00001111_10110011_11000010_0;
      patterns[4022] = 25'b00001111_10110100_11000011_0;
      patterns[4023] = 25'b00001111_10110101_11000100_0;
      patterns[4024] = 25'b00001111_10110110_11000101_0;
      patterns[4025] = 25'b00001111_10110111_11000110_0;
      patterns[4026] = 25'b00001111_10111000_11000111_0;
      patterns[4027] = 25'b00001111_10111001_11001000_0;
      patterns[4028] = 25'b00001111_10111010_11001001_0;
      patterns[4029] = 25'b00001111_10111011_11001010_0;
      patterns[4030] = 25'b00001111_10111100_11001011_0;
      patterns[4031] = 25'b00001111_10111101_11001100_0;
      patterns[4032] = 25'b00001111_10111110_11001101_0;
      patterns[4033] = 25'b00001111_10111111_11001110_0;
      patterns[4034] = 25'b00001111_11000000_11001111_0;
      patterns[4035] = 25'b00001111_11000001_11010000_0;
      patterns[4036] = 25'b00001111_11000010_11010001_0;
      patterns[4037] = 25'b00001111_11000011_11010010_0;
      patterns[4038] = 25'b00001111_11000100_11010011_0;
      patterns[4039] = 25'b00001111_11000101_11010100_0;
      patterns[4040] = 25'b00001111_11000110_11010101_0;
      patterns[4041] = 25'b00001111_11000111_11010110_0;
      patterns[4042] = 25'b00001111_11001000_11010111_0;
      patterns[4043] = 25'b00001111_11001001_11011000_0;
      patterns[4044] = 25'b00001111_11001010_11011001_0;
      patterns[4045] = 25'b00001111_11001011_11011010_0;
      patterns[4046] = 25'b00001111_11001100_11011011_0;
      patterns[4047] = 25'b00001111_11001101_11011100_0;
      patterns[4048] = 25'b00001111_11001110_11011101_0;
      patterns[4049] = 25'b00001111_11001111_11011110_0;
      patterns[4050] = 25'b00001111_11010000_11011111_0;
      patterns[4051] = 25'b00001111_11010001_11100000_0;
      patterns[4052] = 25'b00001111_11010010_11100001_0;
      patterns[4053] = 25'b00001111_11010011_11100010_0;
      patterns[4054] = 25'b00001111_11010100_11100011_0;
      patterns[4055] = 25'b00001111_11010101_11100100_0;
      patterns[4056] = 25'b00001111_11010110_11100101_0;
      patterns[4057] = 25'b00001111_11010111_11100110_0;
      patterns[4058] = 25'b00001111_11011000_11100111_0;
      patterns[4059] = 25'b00001111_11011001_11101000_0;
      patterns[4060] = 25'b00001111_11011010_11101001_0;
      patterns[4061] = 25'b00001111_11011011_11101010_0;
      patterns[4062] = 25'b00001111_11011100_11101011_0;
      patterns[4063] = 25'b00001111_11011101_11101100_0;
      patterns[4064] = 25'b00001111_11011110_11101101_0;
      patterns[4065] = 25'b00001111_11011111_11101110_0;
      patterns[4066] = 25'b00001111_11100000_11101111_0;
      patterns[4067] = 25'b00001111_11100001_11110000_0;
      patterns[4068] = 25'b00001111_11100010_11110001_0;
      patterns[4069] = 25'b00001111_11100011_11110010_0;
      patterns[4070] = 25'b00001111_11100100_11110011_0;
      patterns[4071] = 25'b00001111_11100101_11110100_0;
      patterns[4072] = 25'b00001111_11100110_11110101_0;
      patterns[4073] = 25'b00001111_11100111_11110110_0;
      patterns[4074] = 25'b00001111_11101000_11110111_0;
      patterns[4075] = 25'b00001111_11101001_11111000_0;
      patterns[4076] = 25'b00001111_11101010_11111001_0;
      patterns[4077] = 25'b00001111_11101011_11111010_0;
      patterns[4078] = 25'b00001111_11101100_11111011_0;
      patterns[4079] = 25'b00001111_11101101_11111100_0;
      patterns[4080] = 25'b00001111_11101110_11111101_0;
      patterns[4081] = 25'b00001111_11101111_11111110_0;
      patterns[4082] = 25'b00001111_11110000_11111111_0;
      patterns[4083] = 25'b00001111_11110001_00000000_1;
      patterns[4084] = 25'b00001111_11110010_00000001_1;
      patterns[4085] = 25'b00001111_11110011_00000010_1;
      patterns[4086] = 25'b00001111_11110100_00000011_1;
      patterns[4087] = 25'b00001111_11110101_00000100_1;
      patterns[4088] = 25'b00001111_11110110_00000101_1;
      patterns[4089] = 25'b00001111_11110111_00000110_1;
      patterns[4090] = 25'b00001111_11111000_00000111_1;
      patterns[4091] = 25'b00001111_11111001_00001000_1;
      patterns[4092] = 25'b00001111_11111010_00001001_1;
      patterns[4093] = 25'b00001111_11111011_00001010_1;
      patterns[4094] = 25'b00001111_11111100_00001011_1;
      patterns[4095] = 25'b00001111_11111101_00001100_1;
      patterns[4096] = 25'b00001111_11111110_00001101_1;
      patterns[4097] = 25'b00001111_11111111_00001110_1;
      patterns[4098] = 25'b00010000_00000000_00010000_0;
      patterns[4099] = 25'b00010000_00000001_00010001_0;
      patterns[4100] = 25'b00010000_00000010_00010010_0;
      patterns[4101] = 25'b00010000_00000011_00010011_0;
      patterns[4102] = 25'b00010000_00000100_00010100_0;
      patterns[4103] = 25'b00010000_00000101_00010101_0;
      patterns[4104] = 25'b00010000_00000110_00010110_0;
      patterns[4105] = 25'b00010000_00000111_00010111_0;
      patterns[4106] = 25'b00010000_00001000_00011000_0;
      patterns[4107] = 25'b00010000_00001001_00011001_0;
      patterns[4108] = 25'b00010000_00001010_00011010_0;
      patterns[4109] = 25'b00010000_00001011_00011011_0;
      patterns[4110] = 25'b00010000_00001100_00011100_0;
      patterns[4111] = 25'b00010000_00001101_00011101_0;
      patterns[4112] = 25'b00010000_00001110_00011110_0;
      patterns[4113] = 25'b00010000_00001111_00011111_0;
      patterns[4114] = 25'b00010000_00010000_00100000_0;
      patterns[4115] = 25'b00010000_00010001_00100001_0;
      patterns[4116] = 25'b00010000_00010010_00100010_0;
      patterns[4117] = 25'b00010000_00010011_00100011_0;
      patterns[4118] = 25'b00010000_00010100_00100100_0;
      patterns[4119] = 25'b00010000_00010101_00100101_0;
      patterns[4120] = 25'b00010000_00010110_00100110_0;
      patterns[4121] = 25'b00010000_00010111_00100111_0;
      patterns[4122] = 25'b00010000_00011000_00101000_0;
      patterns[4123] = 25'b00010000_00011001_00101001_0;
      patterns[4124] = 25'b00010000_00011010_00101010_0;
      patterns[4125] = 25'b00010000_00011011_00101011_0;
      patterns[4126] = 25'b00010000_00011100_00101100_0;
      patterns[4127] = 25'b00010000_00011101_00101101_0;
      patterns[4128] = 25'b00010000_00011110_00101110_0;
      patterns[4129] = 25'b00010000_00011111_00101111_0;
      patterns[4130] = 25'b00010000_00100000_00110000_0;
      patterns[4131] = 25'b00010000_00100001_00110001_0;
      patterns[4132] = 25'b00010000_00100010_00110010_0;
      patterns[4133] = 25'b00010000_00100011_00110011_0;
      patterns[4134] = 25'b00010000_00100100_00110100_0;
      patterns[4135] = 25'b00010000_00100101_00110101_0;
      patterns[4136] = 25'b00010000_00100110_00110110_0;
      patterns[4137] = 25'b00010000_00100111_00110111_0;
      patterns[4138] = 25'b00010000_00101000_00111000_0;
      patterns[4139] = 25'b00010000_00101001_00111001_0;
      patterns[4140] = 25'b00010000_00101010_00111010_0;
      patterns[4141] = 25'b00010000_00101011_00111011_0;
      patterns[4142] = 25'b00010000_00101100_00111100_0;
      patterns[4143] = 25'b00010000_00101101_00111101_0;
      patterns[4144] = 25'b00010000_00101110_00111110_0;
      patterns[4145] = 25'b00010000_00101111_00111111_0;
      patterns[4146] = 25'b00010000_00110000_01000000_0;
      patterns[4147] = 25'b00010000_00110001_01000001_0;
      patterns[4148] = 25'b00010000_00110010_01000010_0;
      patterns[4149] = 25'b00010000_00110011_01000011_0;
      patterns[4150] = 25'b00010000_00110100_01000100_0;
      patterns[4151] = 25'b00010000_00110101_01000101_0;
      patterns[4152] = 25'b00010000_00110110_01000110_0;
      patterns[4153] = 25'b00010000_00110111_01000111_0;
      patterns[4154] = 25'b00010000_00111000_01001000_0;
      patterns[4155] = 25'b00010000_00111001_01001001_0;
      patterns[4156] = 25'b00010000_00111010_01001010_0;
      patterns[4157] = 25'b00010000_00111011_01001011_0;
      patterns[4158] = 25'b00010000_00111100_01001100_0;
      patterns[4159] = 25'b00010000_00111101_01001101_0;
      patterns[4160] = 25'b00010000_00111110_01001110_0;
      patterns[4161] = 25'b00010000_00111111_01001111_0;
      patterns[4162] = 25'b00010000_01000000_01010000_0;
      patterns[4163] = 25'b00010000_01000001_01010001_0;
      patterns[4164] = 25'b00010000_01000010_01010010_0;
      patterns[4165] = 25'b00010000_01000011_01010011_0;
      patterns[4166] = 25'b00010000_01000100_01010100_0;
      patterns[4167] = 25'b00010000_01000101_01010101_0;
      patterns[4168] = 25'b00010000_01000110_01010110_0;
      patterns[4169] = 25'b00010000_01000111_01010111_0;
      patterns[4170] = 25'b00010000_01001000_01011000_0;
      patterns[4171] = 25'b00010000_01001001_01011001_0;
      patterns[4172] = 25'b00010000_01001010_01011010_0;
      patterns[4173] = 25'b00010000_01001011_01011011_0;
      patterns[4174] = 25'b00010000_01001100_01011100_0;
      patterns[4175] = 25'b00010000_01001101_01011101_0;
      patterns[4176] = 25'b00010000_01001110_01011110_0;
      patterns[4177] = 25'b00010000_01001111_01011111_0;
      patterns[4178] = 25'b00010000_01010000_01100000_0;
      patterns[4179] = 25'b00010000_01010001_01100001_0;
      patterns[4180] = 25'b00010000_01010010_01100010_0;
      patterns[4181] = 25'b00010000_01010011_01100011_0;
      patterns[4182] = 25'b00010000_01010100_01100100_0;
      patterns[4183] = 25'b00010000_01010101_01100101_0;
      patterns[4184] = 25'b00010000_01010110_01100110_0;
      patterns[4185] = 25'b00010000_01010111_01100111_0;
      patterns[4186] = 25'b00010000_01011000_01101000_0;
      patterns[4187] = 25'b00010000_01011001_01101001_0;
      patterns[4188] = 25'b00010000_01011010_01101010_0;
      patterns[4189] = 25'b00010000_01011011_01101011_0;
      patterns[4190] = 25'b00010000_01011100_01101100_0;
      patterns[4191] = 25'b00010000_01011101_01101101_0;
      patterns[4192] = 25'b00010000_01011110_01101110_0;
      patterns[4193] = 25'b00010000_01011111_01101111_0;
      patterns[4194] = 25'b00010000_01100000_01110000_0;
      patterns[4195] = 25'b00010000_01100001_01110001_0;
      patterns[4196] = 25'b00010000_01100010_01110010_0;
      patterns[4197] = 25'b00010000_01100011_01110011_0;
      patterns[4198] = 25'b00010000_01100100_01110100_0;
      patterns[4199] = 25'b00010000_01100101_01110101_0;
      patterns[4200] = 25'b00010000_01100110_01110110_0;
      patterns[4201] = 25'b00010000_01100111_01110111_0;
      patterns[4202] = 25'b00010000_01101000_01111000_0;
      patterns[4203] = 25'b00010000_01101001_01111001_0;
      patterns[4204] = 25'b00010000_01101010_01111010_0;
      patterns[4205] = 25'b00010000_01101011_01111011_0;
      patterns[4206] = 25'b00010000_01101100_01111100_0;
      patterns[4207] = 25'b00010000_01101101_01111101_0;
      patterns[4208] = 25'b00010000_01101110_01111110_0;
      patterns[4209] = 25'b00010000_01101111_01111111_0;
      patterns[4210] = 25'b00010000_01110000_10000000_0;
      patterns[4211] = 25'b00010000_01110001_10000001_0;
      patterns[4212] = 25'b00010000_01110010_10000010_0;
      patterns[4213] = 25'b00010000_01110011_10000011_0;
      patterns[4214] = 25'b00010000_01110100_10000100_0;
      patterns[4215] = 25'b00010000_01110101_10000101_0;
      patterns[4216] = 25'b00010000_01110110_10000110_0;
      patterns[4217] = 25'b00010000_01110111_10000111_0;
      patterns[4218] = 25'b00010000_01111000_10001000_0;
      patterns[4219] = 25'b00010000_01111001_10001001_0;
      patterns[4220] = 25'b00010000_01111010_10001010_0;
      patterns[4221] = 25'b00010000_01111011_10001011_0;
      patterns[4222] = 25'b00010000_01111100_10001100_0;
      patterns[4223] = 25'b00010000_01111101_10001101_0;
      patterns[4224] = 25'b00010000_01111110_10001110_0;
      patterns[4225] = 25'b00010000_01111111_10001111_0;
      patterns[4226] = 25'b00010000_10000000_10010000_0;
      patterns[4227] = 25'b00010000_10000001_10010001_0;
      patterns[4228] = 25'b00010000_10000010_10010010_0;
      patterns[4229] = 25'b00010000_10000011_10010011_0;
      patterns[4230] = 25'b00010000_10000100_10010100_0;
      patterns[4231] = 25'b00010000_10000101_10010101_0;
      patterns[4232] = 25'b00010000_10000110_10010110_0;
      patterns[4233] = 25'b00010000_10000111_10010111_0;
      patterns[4234] = 25'b00010000_10001000_10011000_0;
      patterns[4235] = 25'b00010000_10001001_10011001_0;
      patterns[4236] = 25'b00010000_10001010_10011010_0;
      patterns[4237] = 25'b00010000_10001011_10011011_0;
      patterns[4238] = 25'b00010000_10001100_10011100_0;
      patterns[4239] = 25'b00010000_10001101_10011101_0;
      patterns[4240] = 25'b00010000_10001110_10011110_0;
      patterns[4241] = 25'b00010000_10001111_10011111_0;
      patterns[4242] = 25'b00010000_10010000_10100000_0;
      patterns[4243] = 25'b00010000_10010001_10100001_0;
      patterns[4244] = 25'b00010000_10010010_10100010_0;
      patterns[4245] = 25'b00010000_10010011_10100011_0;
      patterns[4246] = 25'b00010000_10010100_10100100_0;
      patterns[4247] = 25'b00010000_10010101_10100101_0;
      patterns[4248] = 25'b00010000_10010110_10100110_0;
      patterns[4249] = 25'b00010000_10010111_10100111_0;
      patterns[4250] = 25'b00010000_10011000_10101000_0;
      patterns[4251] = 25'b00010000_10011001_10101001_0;
      patterns[4252] = 25'b00010000_10011010_10101010_0;
      patterns[4253] = 25'b00010000_10011011_10101011_0;
      patterns[4254] = 25'b00010000_10011100_10101100_0;
      patterns[4255] = 25'b00010000_10011101_10101101_0;
      patterns[4256] = 25'b00010000_10011110_10101110_0;
      patterns[4257] = 25'b00010000_10011111_10101111_0;
      patterns[4258] = 25'b00010000_10100000_10110000_0;
      patterns[4259] = 25'b00010000_10100001_10110001_0;
      patterns[4260] = 25'b00010000_10100010_10110010_0;
      patterns[4261] = 25'b00010000_10100011_10110011_0;
      patterns[4262] = 25'b00010000_10100100_10110100_0;
      patterns[4263] = 25'b00010000_10100101_10110101_0;
      patterns[4264] = 25'b00010000_10100110_10110110_0;
      patterns[4265] = 25'b00010000_10100111_10110111_0;
      patterns[4266] = 25'b00010000_10101000_10111000_0;
      patterns[4267] = 25'b00010000_10101001_10111001_0;
      patterns[4268] = 25'b00010000_10101010_10111010_0;
      patterns[4269] = 25'b00010000_10101011_10111011_0;
      patterns[4270] = 25'b00010000_10101100_10111100_0;
      patterns[4271] = 25'b00010000_10101101_10111101_0;
      patterns[4272] = 25'b00010000_10101110_10111110_0;
      patterns[4273] = 25'b00010000_10101111_10111111_0;
      patterns[4274] = 25'b00010000_10110000_11000000_0;
      patterns[4275] = 25'b00010000_10110001_11000001_0;
      patterns[4276] = 25'b00010000_10110010_11000010_0;
      patterns[4277] = 25'b00010000_10110011_11000011_0;
      patterns[4278] = 25'b00010000_10110100_11000100_0;
      patterns[4279] = 25'b00010000_10110101_11000101_0;
      patterns[4280] = 25'b00010000_10110110_11000110_0;
      patterns[4281] = 25'b00010000_10110111_11000111_0;
      patterns[4282] = 25'b00010000_10111000_11001000_0;
      patterns[4283] = 25'b00010000_10111001_11001001_0;
      patterns[4284] = 25'b00010000_10111010_11001010_0;
      patterns[4285] = 25'b00010000_10111011_11001011_0;
      patterns[4286] = 25'b00010000_10111100_11001100_0;
      patterns[4287] = 25'b00010000_10111101_11001101_0;
      patterns[4288] = 25'b00010000_10111110_11001110_0;
      patterns[4289] = 25'b00010000_10111111_11001111_0;
      patterns[4290] = 25'b00010000_11000000_11010000_0;
      patterns[4291] = 25'b00010000_11000001_11010001_0;
      patterns[4292] = 25'b00010000_11000010_11010010_0;
      patterns[4293] = 25'b00010000_11000011_11010011_0;
      patterns[4294] = 25'b00010000_11000100_11010100_0;
      patterns[4295] = 25'b00010000_11000101_11010101_0;
      patterns[4296] = 25'b00010000_11000110_11010110_0;
      patterns[4297] = 25'b00010000_11000111_11010111_0;
      patterns[4298] = 25'b00010000_11001000_11011000_0;
      patterns[4299] = 25'b00010000_11001001_11011001_0;
      patterns[4300] = 25'b00010000_11001010_11011010_0;
      patterns[4301] = 25'b00010000_11001011_11011011_0;
      patterns[4302] = 25'b00010000_11001100_11011100_0;
      patterns[4303] = 25'b00010000_11001101_11011101_0;
      patterns[4304] = 25'b00010000_11001110_11011110_0;
      patterns[4305] = 25'b00010000_11001111_11011111_0;
      patterns[4306] = 25'b00010000_11010000_11100000_0;
      patterns[4307] = 25'b00010000_11010001_11100001_0;
      patterns[4308] = 25'b00010000_11010010_11100010_0;
      patterns[4309] = 25'b00010000_11010011_11100011_0;
      patterns[4310] = 25'b00010000_11010100_11100100_0;
      patterns[4311] = 25'b00010000_11010101_11100101_0;
      patterns[4312] = 25'b00010000_11010110_11100110_0;
      patterns[4313] = 25'b00010000_11010111_11100111_0;
      patterns[4314] = 25'b00010000_11011000_11101000_0;
      patterns[4315] = 25'b00010000_11011001_11101001_0;
      patterns[4316] = 25'b00010000_11011010_11101010_0;
      patterns[4317] = 25'b00010000_11011011_11101011_0;
      patterns[4318] = 25'b00010000_11011100_11101100_0;
      patterns[4319] = 25'b00010000_11011101_11101101_0;
      patterns[4320] = 25'b00010000_11011110_11101110_0;
      patterns[4321] = 25'b00010000_11011111_11101111_0;
      patterns[4322] = 25'b00010000_11100000_11110000_0;
      patterns[4323] = 25'b00010000_11100001_11110001_0;
      patterns[4324] = 25'b00010000_11100010_11110010_0;
      patterns[4325] = 25'b00010000_11100011_11110011_0;
      patterns[4326] = 25'b00010000_11100100_11110100_0;
      patterns[4327] = 25'b00010000_11100101_11110101_0;
      patterns[4328] = 25'b00010000_11100110_11110110_0;
      patterns[4329] = 25'b00010000_11100111_11110111_0;
      patterns[4330] = 25'b00010000_11101000_11111000_0;
      patterns[4331] = 25'b00010000_11101001_11111001_0;
      patterns[4332] = 25'b00010000_11101010_11111010_0;
      patterns[4333] = 25'b00010000_11101011_11111011_0;
      patterns[4334] = 25'b00010000_11101100_11111100_0;
      patterns[4335] = 25'b00010000_11101101_11111101_0;
      patterns[4336] = 25'b00010000_11101110_11111110_0;
      patterns[4337] = 25'b00010000_11101111_11111111_0;
      patterns[4338] = 25'b00010000_11110000_00000000_1;
      patterns[4339] = 25'b00010000_11110001_00000001_1;
      patterns[4340] = 25'b00010000_11110010_00000010_1;
      patterns[4341] = 25'b00010000_11110011_00000011_1;
      patterns[4342] = 25'b00010000_11110100_00000100_1;
      patterns[4343] = 25'b00010000_11110101_00000101_1;
      patterns[4344] = 25'b00010000_11110110_00000110_1;
      patterns[4345] = 25'b00010000_11110111_00000111_1;
      patterns[4346] = 25'b00010000_11111000_00001000_1;
      patterns[4347] = 25'b00010000_11111001_00001001_1;
      patterns[4348] = 25'b00010000_11111010_00001010_1;
      patterns[4349] = 25'b00010000_11111011_00001011_1;
      patterns[4350] = 25'b00010000_11111100_00001100_1;
      patterns[4351] = 25'b00010000_11111101_00001101_1;
      patterns[4352] = 25'b00010000_11111110_00001110_1;
      patterns[4353] = 25'b00010000_11111111_00001111_1;
      patterns[4354] = 25'b00010001_00000000_00010001_0;
      patterns[4355] = 25'b00010001_00000001_00010010_0;
      patterns[4356] = 25'b00010001_00000010_00010011_0;
      patterns[4357] = 25'b00010001_00000011_00010100_0;
      patterns[4358] = 25'b00010001_00000100_00010101_0;
      patterns[4359] = 25'b00010001_00000101_00010110_0;
      patterns[4360] = 25'b00010001_00000110_00010111_0;
      patterns[4361] = 25'b00010001_00000111_00011000_0;
      patterns[4362] = 25'b00010001_00001000_00011001_0;
      patterns[4363] = 25'b00010001_00001001_00011010_0;
      patterns[4364] = 25'b00010001_00001010_00011011_0;
      patterns[4365] = 25'b00010001_00001011_00011100_0;
      patterns[4366] = 25'b00010001_00001100_00011101_0;
      patterns[4367] = 25'b00010001_00001101_00011110_0;
      patterns[4368] = 25'b00010001_00001110_00011111_0;
      patterns[4369] = 25'b00010001_00001111_00100000_0;
      patterns[4370] = 25'b00010001_00010000_00100001_0;
      patterns[4371] = 25'b00010001_00010001_00100010_0;
      patterns[4372] = 25'b00010001_00010010_00100011_0;
      patterns[4373] = 25'b00010001_00010011_00100100_0;
      patterns[4374] = 25'b00010001_00010100_00100101_0;
      patterns[4375] = 25'b00010001_00010101_00100110_0;
      patterns[4376] = 25'b00010001_00010110_00100111_0;
      patterns[4377] = 25'b00010001_00010111_00101000_0;
      patterns[4378] = 25'b00010001_00011000_00101001_0;
      patterns[4379] = 25'b00010001_00011001_00101010_0;
      patterns[4380] = 25'b00010001_00011010_00101011_0;
      patterns[4381] = 25'b00010001_00011011_00101100_0;
      patterns[4382] = 25'b00010001_00011100_00101101_0;
      patterns[4383] = 25'b00010001_00011101_00101110_0;
      patterns[4384] = 25'b00010001_00011110_00101111_0;
      patterns[4385] = 25'b00010001_00011111_00110000_0;
      patterns[4386] = 25'b00010001_00100000_00110001_0;
      patterns[4387] = 25'b00010001_00100001_00110010_0;
      patterns[4388] = 25'b00010001_00100010_00110011_0;
      patterns[4389] = 25'b00010001_00100011_00110100_0;
      patterns[4390] = 25'b00010001_00100100_00110101_0;
      patterns[4391] = 25'b00010001_00100101_00110110_0;
      patterns[4392] = 25'b00010001_00100110_00110111_0;
      patterns[4393] = 25'b00010001_00100111_00111000_0;
      patterns[4394] = 25'b00010001_00101000_00111001_0;
      patterns[4395] = 25'b00010001_00101001_00111010_0;
      patterns[4396] = 25'b00010001_00101010_00111011_0;
      patterns[4397] = 25'b00010001_00101011_00111100_0;
      patterns[4398] = 25'b00010001_00101100_00111101_0;
      patterns[4399] = 25'b00010001_00101101_00111110_0;
      patterns[4400] = 25'b00010001_00101110_00111111_0;
      patterns[4401] = 25'b00010001_00101111_01000000_0;
      patterns[4402] = 25'b00010001_00110000_01000001_0;
      patterns[4403] = 25'b00010001_00110001_01000010_0;
      patterns[4404] = 25'b00010001_00110010_01000011_0;
      patterns[4405] = 25'b00010001_00110011_01000100_0;
      patterns[4406] = 25'b00010001_00110100_01000101_0;
      patterns[4407] = 25'b00010001_00110101_01000110_0;
      patterns[4408] = 25'b00010001_00110110_01000111_0;
      patterns[4409] = 25'b00010001_00110111_01001000_0;
      patterns[4410] = 25'b00010001_00111000_01001001_0;
      patterns[4411] = 25'b00010001_00111001_01001010_0;
      patterns[4412] = 25'b00010001_00111010_01001011_0;
      patterns[4413] = 25'b00010001_00111011_01001100_0;
      patterns[4414] = 25'b00010001_00111100_01001101_0;
      patterns[4415] = 25'b00010001_00111101_01001110_0;
      patterns[4416] = 25'b00010001_00111110_01001111_0;
      patterns[4417] = 25'b00010001_00111111_01010000_0;
      patterns[4418] = 25'b00010001_01000000_01010001_0;
      patterns[4419] = 25'b00010001_01000001_01010010_0;
      patterns[4420] = 25'b00010001_01000010_01010011_0;
      patterns[4421] = 25'b00010001_01000011_01010100_0;
      patterns[4422] = 25'b00010001_01000100_01010101_0;
      patterns[4423] = 25'b00010001_01000101_01010110_0;
      patterns[4424] = 25'b00010001_01000110_01010111_0;
      patterns[4425] = 25'b00010001_01000111_01011000_0;
      patterns[4426] = 25'b00010001_01001000_01011001_0;
      patterns[4427] = 25'b00010001_01001001_01011010_0;
      patterns[4428] = 25'b00010001_01001010_01011011_0;
      patterns[4429] = 25'b00010001_01001011_01011100_0;
      patterns[4430] = 25'b00010001_01001100_01011101_0;
      patterns[4431] = 25'b00010001_01001101_01011110_0;
      patterns[4432] = 25'b00010001_01001110_01011111_0;
      patterns[4433] = 25'b00010001_01001111_01100000_0;
      patterns[4434] = 25'b00010001_01010000_01100001_0;
      patterns[4435] = 25'b00010001_01010001_01100010_0;
      patterns[4436] = 25'b00010001_01010010_01100011_0;
      patterns[4437] = 25'b00010001_01010011_01100100_0;
      patterns[4438] = 25'b00010001_01010100_01100101_0;
      patterns[4439] = 25'b00010001_01010101_01100110_0;
      patterns[4440] = 25'b00010001_01010110_01100111_0;
      patterns[4441] = 25'b00010001_01010111_01101000_0;
      patterns[4442] = 25'b00010001_01011000_01101001_0;
      patterns[4443] = 25'b00010001_01011001_01101010_0;
      patterns[4444] = 25'b00010001_01011010_01101011_0;
      patterns[4445] = 25'b00010001_01011011_01101100_0;
      patterns[4446] = 25'b00010001_01011100_01101101_0;
      patterns[4447] = 25'b00010001_01011101_01101110_0;
      patterns[4448] = 25'b00010001_01011110_01101111_0;
      patterns[4449] = 25'b00010001_01011111_01110000_0;
      patterns[4450] = 25'b00010001_01100000_01110001_0;
      patterns[4451] = 25'b00010001_01100001_01110010_0;
      patterns[4452] = 25'b00010001_01100010_01110011_0;
      patterns[4453] = 25'b00010001_01100011_01110100_0;
      patterns[4454] = 25'b00010001_01100100_01110101_0;
      patterns[4455] = 25'b00010001_01100101_01110110_0;
      patterns[4456] = 25'b00010001_01100110_01110111_0;
      patterns[4457] = 25'b00010001_01100111_01111000_0;
      patterns[4458] = 25'b00010001_01101000_01111001_0;
      patterns[4459] = 25'b00010001_01101001_01111010_0;
      patterns[4460] = 25'b00010001_01101010_01111011_0;
      patterns[4461] = 25'b00010001_01101011_01111100_0;
      patterns[4462] = 25'b00010001_01101100_01111101_0;
      patterns[4463] = 25'b00010001_01101101_01111110_0;
      patterns[4464] = 25'b00010001_01101110_01111111_0;
      patterns[4465] = 25'b00010001_01101111_10000000_0;
      patterns[4466] = 25'b00010001_01110000_10000001_0;
      patterns[4467] = 25'b00010001_01110001_10000010_0;
      patterns[4468] = 25'b00010001_01110010_10000011_0;
      patterns[4469] = 25'b00010001_01110011_10000100_0;
      patterns[4470] = 25'b00010001_01110100_10000101_0;
      patterns[4471] = 25'b00010001_01110101_10000110_0;
      patterns[4472] = 25'b00010001_01110110_10000111_0;
      patterns[4473] = 25'b00010001_01110111_10001000_0;
      patterns[4474] = 25'b00010001_01111000_10001001_0;
      patterns[4475] = 25'b00010001_01111001_10001010_0;
      patterns[4476] = 25'b00010001_01111010_10001011_0;
      patterns[4477] = 25'b00010001_01111011_10001100_0;
      patterns[4478] = 25'b00010001_01111100_10001101_0;
      patterns[4479] = 25'b00010001_01111101_10001110_0;
      patterns[4480] = 25'b00010001_01111110_10001111_0;
      patterns[4481] = 25'b00010001_01111111_10010000_0;
      patterns[4482] = 25'b00010001_10000000_10010001_0;
      patterns[4483] = 25'b00010001_10000001_10010010_0;
      patterns[4484] = 25'b00010001_10000010_10010011_0;
      patterns[4485] = 25'b00010001_10000011_10010100_0;
      patterns[4486] = 25'b00010001_10000100_10010101_0;
      patterns[4487] = 25'b00010001_10000101_10010110_0;
      patterns[4488] = 25'b00010001_10000110_10010111_0;
      patterns[4489] = 25'b00010001_10000111_10011000_0;
      patterns[4490] = 25'b00010001_10001000_10011001_0;
      patterns[4491] = 25'b00010001_10001001_10011010_0;
      patterns[4492] = 25'b00010001_10001010_10011011_0;
      patterns[4493] = 25'b00010001_10001011_10011100_0;
      patterns[4494] = 25'b00010001_10001100_10011101_0;
      patterns[4495] = 25'b00010001_10001101_10011110_0;
      patterns[4496] = 25'b00010001_10001110_10011111_0;
      patterns[4497] = 25'b00010001_10001111_10100000_0;
      patterns[4498] = 25'b00010001_10010000_10100001_0;
      patterns[4499] = 25'b00010001_10010001_10100010_0;
      patterns[4500] = 25'b00010001_10010010_10100011_0;
      patterns[4501] = 25'b00010001_10010011_10100100_0;
      patterns[4502] = 25'b00010001_10010100_10100101_0;
      patterns[4503] = 25'b00010001_10010101_10100110_0;
      patterns[4504] = 25'b00010001_10010110_10100111_0;
      patterns[4505] = 25'b00010001_10010111_10101000_0;
      patterns[4506] = 25'b00010001_10011000_10101001_0;
      patterns[4507] = 25'b00010001_10011001_10101010_0;
      patterns[4508] = 25'b00010001_10011010_10101011_0;
      patterns[4509] = 25'b00010001_10011011_10101100_0;
      patterns[4510] = 25'b00010001_10011100_10101101_0;
      patterns[4511] = 25'b00010001_10011101_10101110_0;
      patterns[4512] = 25'b00010001_10011110_10101111_0;
      patterns[4513] = 25'b00010001_10011111_10110000_0;
      patterns[4514] = 25'b00010001_10100000_10110001_0;
      patterns[4515] = 25'b00010001_10100001_10110010_0;
      patterns[4516] = 25'b00010001_10100010_10110011_0;
      patterns[4517] = 25'b00010001_10100011_10110100_0;
      patterns[4518] = 25'b00010001_10100100_10110101_0;
      patterns[4519] = 25'b00010001_10100101_10110110_0;
      patterns[4520] = 25'b00010001_10100110_10110111_0;
      patterns[4521] = 25'b00010001_10100111_10111000_0;
      patterns[4522] = 25'b00010001_10101000_10111001_0;
      patterns[4523] = 25'b00010001_10101001_10111010_0;
      patterns[4524] = 25'b00010001_10101010_10111011_0;
      patterns[4525] = 25'b00010001_10101011_10111100_0;
      patterns[4526] = 25'b00010001_10101100_10111101_0;
      patterns[4527] = 25'b00010001_10101101_10111110_0;
      patterns[4528] = 25'b00010001_10101110_10111111_0;
      patterns[4529] = 25'b00010001_10101111_11000000_0;
      patterns[4530] = 25'b00010001_10110000_11000001_0;
      patterns[4531] = 25'b00010001_10110001_11000010_0;
      patterns[4532] = 25'b00010001_10110010_11000011_0;
      patterns[4533] = 25'b00010001_10110011_11000100_0;
      patterns[4534] = 25'b00010001_10110100_11000101_0;
      patterns[4535] = 25'b00010001_10110101_11000110_0;
      patterns[4536] = 25'b00010001_10110110_11000111_0;
      patterns[4537] = 25'b00010001_10110111_11001000_0;
      patterns[4538] = 25'b00010001_10111000_11001001_0;
      patterns[4539] = 25'b00010001_10111001_11001010_0;
      patterns[4540] = 25'b00010001_10111010_11001011_0;
      patterns[4541] = 25'b00010001_10111011_11001100_0;
      patterns[4542] = 25'b00010001_10111100_11001101_0;
      patterns[4543] = 25'b00010001_10111101_11001110_0;
      patterns[4544] = 25'b00010001_10111110_11001111_0;
      patterns[4545] = 25'b00010001_10111111_11010000_0;
      patterns[4546] = 25'b00010001_11000000_11010001_0;
      patterns[4547] = 25'b00010001_11000001_11010010_0;
      patterns[4548] = 25'b00010001_11000010_11010011_0;
      patterns[4549] = 25'b00010001_11000011_11010100_0;
      patterns[4550] = 25'b00010001_11000100_11010101_0;
      patterns[4551] = 25'b00010001_11000101_11010110_0;
      patterns[4552] = 25'b00010001_11000110_11010111_0;
      patterns[4553] = 25'b00010001_11000111_11011000_0;
      patterns[4554] = 25'b00010001_11001000_11011001_0;
      patterns[4555] = 25'b00010001_11001001_11011010_0;
      patterns[4556] = 25'b00010001_11001010_11011011_0;
      patterns[4557] = 25'b00010001_11001011_11011100_0;
      patterns[4558] = 25'b00010001_11001100_11011101_0;
      patterns[4559] = 25'b00010001_11001101_11011110_0;
      patterns[4560] = 25'b00010001_11001110_11011111_0;
      patterns[4561] = 25'b00010001_11001111_11100000_0;
      patterns[4562] = 25'b00010001_11010000_11100001_0;
      patterns[4563] = 25'b00010001_11010001_11100010_0;
      patterns[4564] = 25'b00010001_11010010_11100011_0;
      patterns[4565] = 25'b00010001_11010011_11100100_0;
      patterns[4566] = 25'b00010001_11010100_11100101_0;
      patterns[4567] = 25'b00010001_11010101_11100110_0;
      patterns[4568] = 25'b00010001_11010110_11100111_0;
      patterns[4569] = 25'b00010001_11010111_11101000_0;
      patterns[4570] = 25'b00010001_11011000_11101001_0;
      patterns[4571] = 25'b00010001_11011001_11101010_0;
      patterns[4572] = 25'b00010001_11011010_11101011_0;
      patterns[4573] = 25'b00010001_11011011_11101100_0;
      patterns[4574] = 25'b00010001_11011100_11101101_0;
      patterns[4575] = 25'b00010001_11011101_11101110_0;
      patterns[4576] = 25'b00010001_11011110_11101111_0;
      patterns[4577] = 25'b00010001_11011111_11110000_0;
      patterns[4578] = 25'b00010001_11100000_11110001_0;
      patterns[4579] = 25'b00010001_11100001_11110010_0;
      patterns[4580] = 25'b00010001_11100010_11110011_0;
      patterns[4581] = 25'b00010001_11100011_11110100_0;
      patterns[4582] = 25'b00010001_11100100_11110101_0;
      patterns[4583] = 25'b00010001_11100101_11110110_0;
      patterns[4584] = 25'b00010001_11100110_11110111_0;
      patterns[4585] = 25'b00010001_11100111_11111000_0;
      patterns[4586] = 25'b00010001_11101000_11111001_0;
      patterns[4587] = 25'b00010001_11101001_11111010_0;
      patterns[4588] = 25'b00010001_11101010_11111011_0;
      patterns[4589] = 25'b00010001_11101011_11111100_0;
      patterns[4590] = 25'b00010001_11101100_11111101_0;
      patterns[4591] = 25'b00010001_11101101_11111110_0;
      patterns[4592] = 25'b00010001_11101110_11111111_0;
      patterns[4593] = 25'b00010001_11101111_00000000_1;
      patterns[4594] = 25'b00010001_11110000_00000001_1;
      patterns[4595] = 25'b00010001_11110001_00000010_1;
      patterns[4596] = 25'b00010001_11110010_00000011_1;
      patterns[4597] = 25'b00010001_11110011_00000100_1;
      patterns[4598] = 25'b00010001_11110100_00000101_1;
      patterns[4599] = 25'b00010001_11110101_00000110_1;
      patterns[4600] = 25'b00010001_11110110_00000111_1;
      patterns[4601] = 25'b00010001_11110111_00001000_1;
      patterns[4602] = 25'b00010001_11111000_00001001_1;
      patterns[4603] = 25'b00010001_11111001_00001010_1;
      patterns[4604] = 25'b00010001_11111010_00001011_1;
      patterns[4605] = 25'b00010001_11111011_00001100_1;
      patterns[4606] = 25'b00010001_11111100_00001101_1;
      patterns[4607] = 25'b00010001_11111101_00001110_1;
      patterns[4608] = 25'b00010001_11111110_00001111_1;
      patterns[4609] = 25'b00010001_11111111_00010000_1;
      patterns[4610] = 25'b00010010_00000000_00010010_0;
      patterns[4611] = 25'b00010010_00000001_00010011_0;
      patterns[4612] = 25'b00010010_00000010_00010100_0;
      patterns[4613] = 25'b00010010_00000011_00010101_0;
      patterns[4614] = 25'b00010010_00000100_00010110_0;
      patterns[4615] = 25'b00010010_00000101_00010111_0;
      patterns[4616] = 25'b00010010_00000110_00011000_0;
      patterns[4617] = 25'b00010010_00000111_00011001_0;
      patterns[4618] = 25'b00010010_00001000_00011010_0;
      patterns[4619] = 25'b00010010_00001001_00011011_0;
      patterns[4620] = 25'b00010010_00001010_00011100_0;
      patterns[4621] = 25'b00010010_00001011_00011101_0;
      patterns[4622] = 25'b00010010_00001100_00011110_0;
      patterns[4623] = 25'b00010010_00001101_00011111_0;
      patterns[4624] = 25'b00010010_00001110_00100000_0;
      patterns[4625] = 25'b00010010_00001111_00100001_0;
      patterns[4626] = 25'b00010010_00010000_00100010_0;
      patterns[4627] = 25'b00010010_00010001_00100011_0;
      patterns[4628] = 25'b00010010_00010010_00100100_0;
      patterns[4629] = 25'b00010010_00010011_00100101_0;
      patterns[4630] = 25'b00010010_00010100_00100110_0;
      patterns[4631] = 25'b00010010_00010101_00100111_0;
      patterns[4632] = 25'b00010010_00010110_00101000_0;
      patterns[4633] = 25'b00010010_00010111_00101001_0;
      patterns[4634] = 25'b00010010_00011000_00101010_0;
      patterns[4635] = 25'b00010010_00011001_00101011_0;
      patterns[4636] = 25'b00010010_00011010_00101100_0;
      patterns[4637] = 25'b00010010_00011011_00101101_0;
      patterns[4638] = 25'b00010010_00011100_00101110_0;
      patterns[4639] = 25'b00010010_00011101_00101111_0;
      patterns[4640] = 25'b00010010_00011110_00110000_0;
      patterns[4641] = 25'b00010010_00011111_00110001_0;
      patterns[4642] = 25'b00010010_00100000_00110010_0;
      patterns[4643] = 25'b00010010_00100001_00110011_0;
      patterns[4644] = 25'b00010010_00100010_00110100_0;
      patterns[4645] = 25'b00010010_00100011_00110101_0;
      patterns[4646] = 25'b00010010_00100100_00110110_0;
      patterns[4647] = 25'b00010010_00100101_00110111_0;
      patterns[4648] = 25'b00010010_00100110_00111000_0;
      patterns[4649] = 25'b00010010_00100111_00111001_0;
      patterns[4650] = 25'b00010010_00101000_00111010_0;
      patterns[4651] = 25'b00010010_00101001_00111011_0;
      patterns[4652] = 25'b00010010_00101010_00111100_0;
      patterns[4653] = 25'b00010010_00101011_00111101_0;
      patterns[4654] = 25'b00010010_00101100_00111110_0;
      patterns[4655] = 25'b00010010_00101101_00111111_0;
      patterns[4656] = 25'b00010010_00101110_01000000_0;
      patterns[4657] = 25'b00010010_00101111_01000001_0;
      patterns[4658] = 25'b00010010_00110000_01000010_0;
      patterns[4659] = 25'b00010010_00110001_01000011_0;
      patterns[4660] = 25'b00010010_00110010_01000100_0;
      patterns[4661] = 25'b00010010_00110011_01000101_0;
      patterns[4662] = 25'b00010010_00110100_01000110_0;
      patterns[4663] = 25'b00010010_00110101_01000111_0;
      patterns[4664] = 25'b00010010_00110110_01001000_0;
      patterns[4665] = 25'b00010010_00110111_01001001_0;
      patterns[4666] = 25'b00010010_00111000_01001010_0;
      patterns[4667] = 25'b00010010_00111001_01001011_0;
      patterns[4668] = 25'b00010010_00111010_01001100_0;
      patterns[4669] = 25'b00010010_00111011_01001101_0;
      patterns[4670] = 25'b00010010_00111100_01001110_0;
      patterns[4671] = 25'b00010010_00111101_01001111_0;
      patterns[4672] = 25'b00010010_00111110_01010000_0;
      patterns[4673] = 25'b00010010_00111111_01010001_0;
      patterns[4674] = 25'b00010010_01000000_01010010_0;
      patterns[4675] = 25'b00010010_01000001_01010011_0;
      patterns[4676] = 25'b00010010_01000010_01010100_0;
      patterns[4677] = 25'b00010010_01000011_01010101_0;
      patterns[4678] = 25'b00010010_01000100_01010110_0;
      patterns[4679] = 25'b00010010_01000101_01010111_0;
      patterns[4680] = 25'b00010010_01000110_01011000_0;
      patterns[4681] = 25'b00010010_01000111_01011001_0;
      patterns[4682] = 25'b00010010_01001000_01011010_0;
      patterns[4683] = 25'b00010010_01001001_01011011_0;
      patterns[4684] = 25'b00010010_01001010_01011100_0;
      patterns[4685] = 25'b00010010_01001011_01011101_0;
      patterns[4686] = 25'b00010010_01001100_01011110_0;
      patterns[4687] = 25'b00010010_01001101_01011111_0;
      patterns[4688] = 25'b00010010_01001110_01100000_0;
      patterns[4689] = 25'b00010010_01001111_01100001_0;
      patterns[4690] = 25'b00010010_01010000_01100010_0;
      patterns[4691] = 25'b00010010_01010001_01100011_0;
      patterns[4692] = 25'b00010010_01010010_01100100_0;
      patterns[4693] = 25'b00010010_01010011_01100101_0;
      patterns[4694] = 25'b00010010_01010100_01100110_0;
      patterns[4695] = 25'b00010010_01010101_01100111_0;
      patterns[4696] = 25'b00010010_01010110_01101000_0;
      patterns[4697] = 25'b00010010_01010111_01101001_0;
      patterns[4698] = 25'b00010010_01011000_01101010_0;
      patterns[4699] = 25'b00010010_01011001_01101011_0;
      patterns[4700] = 25'b00010010_01011010_01101100_0;
      patterns[4701] = 25'b00010010_01011011_01101101_0;
      patterns[4702] = 25'b00010010_01011100_01101110_0;
      patterns[4703] = 25'b00010010_01011101_01101111_0;
      patterns[4704] = 25'b00010010_01011110_01110000_0;
      patterns[4705] = 25'b00010010_01011111_01110001_0;
      patterns[4706] = 25'b00010010_01100000_01110010_0;
      patterns[4707] = 25'b00010010_01100001_01110011_0;
      patterns[4708] = 25'b00010010_01100010_01110100_0;
      patterns[4709] = 25'b00010010_01100011_01110101_0;
      patterns[4710] = 25'b00010010_01100100_01110110_0;
      patterns[4711] = 25'b00010010_01100101_01110111_0;
      patterns[4712] = 25'b00010010_01100110_01111000_0;
      patterns[4713] = 25'b00010010_01100111_01111001_0;
      patterns[4714] = 25'b00010010_01101000_01111010_0;
      patterns[4715] = 25'b00010010_01101001_01111011_0;
      patterns[4716] = 25'b00010010_01101010_01111100_0;
      patterns[4717] = 25'b00010010_01101011_01111101_0;
      patterns[4718] = 25'b00010010_01101100_01111110_0;
      patterns[4719] = 25'b00010010_01101101_01111111_0;
      patterns[4720] = 25'b00010010_01101110_10000000_0;
      patterns[4721] = 25'b00010010_01101111_10000001_0;
      patterns[4722] = 25'b00010010_01110000_10000010_0;
      patterns[4723] = 25'b00010010_01110001_10000011_0;
      patterns[4724] = 25'b00010010_01110010_10000100_0;
      patterns[4725] = 25'b00010010_01110011_10000101_0;
      patterns[4726] = 25'b00010010_01110100_10000110_0;
      patterns[4727] = 25'b00010010_01110101_10000111_0;
      patterns[4728] = 25'b00010010_01110110_10001000_0;
      patterns[4729] = 25'b00010010_01110111_10001001_0;
      patterns[4730] = 25'b00010010_01111000_10001010_0;
      patterns[4731] = 25'b00010010_01111001_10001011_0;
      patterns[4732] = 25'b00010010_01111010_10001100_0;
      patterns[4733] = 25'b00010010_01111011_10001101_0;
      patterns[4734] = 25'b00010010_01111100_10001110_0;
      patterns[4735] = 25'b00010010_01111101_10001111_0;
      patterns[4736] = 25'b00010010_01111110_10010000_0;
      patterns[4737] = 25'b00010010_01111111_10010001_0;
      patterns[4738] = 25'b00010010_10000000_10010010_0;
      patterns[4739] = 25'b00010010_10000001_10010011_0;
      patterns[4740] = 25'b00010010_10000010_10010100_0;
      patterns[4741] = 25'b00010010_10000011_10010101_0;
      patterns[4742] = 25'b00010010_10000100_10010110_0;
      patterns[4743] = 25'b00010010_10000101_10010111_0;
      patterns[4744] = 25'b00010010_10000110_10011000_0;
      patterns[4745] = 25'b00010010_10000111_10011001_0;
      patterns[4746] = 25'b00010010_10001000_10011010_0;
      patterns[4747] = 25'b00010010_10001001_10011011_0;
      patterns[4748] = 25'b00010010_10001010_10011100_0;
      patterns[4749] = 25'b00010010_10001011_10011101_0;
      patterns[4750] = 25'b00010010_10001100_10011110_0;
      patterns[4751] = 25'b00010010_10001101_10011111_0;
      patterns[4752] = 25'b00010010_10001110_10100000_0;
      patterns[4753] = 25'b00010010_10001111_10100001_0;
      patterns[4754] = 25'b00010010_10010000_10100010_0;
      patterns[4755] = 25'b00010010_10010001_10100011_0;
      patterns[4756] = 25'b00010010_10010010_10100100_0;
      patterns[4757] = 25'b00010010_10010011_10100101_0;
      patterns[4758] = 25'b00010010_10010100_10100110_0;
      patterns[4759] = 25'b00010010_10010101_10100111_0;
      patterns[4760] = 25'b00010010_10010110_10101000_0;
      patterns[4761] = 25'b00010010_10010111_10101001_0;
      patterns[4762] = 25'b00010010_10011000_10101010_0;
      patterns[4763] = 25'b00010010_10011001_10101011_0;
      patterns[4764] = 25'b00010010_10011010_10101100_0;
      patterns[4765] = 25'b00010010_10011011_10101101_0;
      patterns[4766] = 25'b00010010_10011100_10101110_0;
      patterns[4767] = 25'b00010010_10011101_10101111_0;
      patterns[4768] = 25'b00010010_10011110_10110000_0;
      patterns[4769] = 25'b00010010_10011111_10110001_0;
      patterns[4770] = 25'b00010010_10100000_10110010_0;
      patterns[4771] = 25'b00010010_10100001_10110011_0;
      patterns[4772] = 25'b00010010_10100010_10110100_0;
      patterns[4773] = 25'b00010010_10100011_10110101_0;
      patterns[4774] = 25'b00010010_10100100_10110110_0;
      patterns[4775] = 25'b00010010_10100101_10110111_0;
      patterns[4776] = 25'b00010010_10100110_10111000_0;
      patterns[4777] = 25'b00010010_10100111_10111001_0;
      patterns[4778] = 25'b00010010_10101000_10111010_0;
      patterns[4779] = 25'b00010010_10101001_10111011_0;
      patterns[4780] = 25'b00010010_10101010_10111100_0;
      patterns[4781] = 25'b00010010_10101011_10111101_0;
      patterns[4782] = 25'b00010010_10101100_10111110_0;
      patterns[4783] = 25'b00010010_10101101_10111111_0;
      patterns[4784] = 25'b00010010_10101110_11000000_0;
      patterns[4785] = 25'b00010010_10101111_11000001_0;
      patterns[4786] = 25'b00010010_10110000_11000010_0;
      patterns[4787] = 25'b00010010_10110001_11000011_0;
      patterns[4788] = 25'b00010010_10110010_11000100_0;
      patterns[4789] = 25'b00010010_10110011_11000101_0;
      patterns[4790] = 25'b00010010_10110100_11000110_0;
      patterns[4791] = 25'b00010010_10110101_11000111_0;
      patterns[4792] = 25'b00010010_10110110_11001000_0;
      patterns[4793] = 25'b00010010_10110111_11001001_0;
      patterns[4794] = 25'b00010010_10111000_11001010_0;
      patterns[4795] = 25'b00010010_10111001_11001011_0;
      patterns[4796] = 25'b00010010_10111010_11001100_0;
      patterns[4797] = 25'b00010010_10111011_11001101_0;
      patterns[4798] = 25'b00010010_10111100_11001110_0;
      patterns[4799] = 25'b00010010_10111101_11001111_0;
      patterns[4800] = 25'b00010010_10111110_11010000_0;
      patterns[4801] = 25'b00010010_10111111_11010001_0;
      patterns[4802] = 25'b00010010_11000000_11010010_0;
      patterns[4803] = 25'b00010010_11000001_11010011_0;
      patterns[4804] = 25'b00010010_11000010_11010100_0;
      patterns[4805] = 25'b00010010_11000011_11010101_0;
      patterns[4806] = 25'b00010010_11000100_11010110_0;
      patterns[4807] = 25'b00010010_11000101_11010111_0;
      patterns[4808] = 25'b00010010_11000110_11011000_0;
      patterns[4809] = 25'b00010010_11000111_11011001_0;
      patterns[4810] = 25'b00010010_11001000_11011010_0;
      patterns[4811] = 25'b00010010_11001001_11011011_0;
      patterns[4812] = 25'b00010010_11001010_11011100_0;
      patterns[4813] = 25'b00010010_11001011_11011101_0;
      patterns[4814] = 25'b00010010_11001100_11011110_0;
      patterns[4815] = 25'b00010010_11001101_11011111_0;
      patterns[4816] = 25'b00010010_11001110_11100000_0;
      patterns[4817] = 25'b00010010_11001111_11100001_0;
      patterns[4818] = 25'b00010010_11010000_11100010_0;
      patterns[4819] = 25'b00010010_11010001_11100011_0;
      patterns[4820] = 25'b00010010_11010010_11100100_0;
      patterns[4821] = 25'b00010010_11010011_11100101_0;
      patterns[4822] = 25'b00010010_11010100_11100110_0;
      patterns[4823] = 25'b00010010_11010101_11100111_0;
      patterns[4824] = 25'b00010010_11010110_11101000_0;
      patterns[4825] = 25'b00010010_11010111_11101001_0;
      patterns[4826] = 25'b00010010_11011000_11101010_0;
      patterns[4827] = 25'b00010010_11011001_11101011_0;
      patterns[4828] = 25'b00010010_11011010_11101100_0;
      patterns[4829] = 25'b00010010_11011011_11101101_0;
      patterns[4830] = 25'b00010010_11011100_11101110_0;
      patterns[4831] = 25'b00010010_11011101_11101111_0;
      patterns[4832] = 25'b00010010_11011110_11110000_0;
      patterns[4833] = 25'b00010010_11011111_11110001_0;
      patterns[4834] = 25'b00010010_11100000_11110010_0;
      patterns[4835] = 25'b00010010_11100001_11110011_0;
      patterns[4836] = 25'b00010010_11100010_11110100_0;
      patterns[4837] = 25'b00010010_11100011_11110101_0;
      patterns[4838] = 25'b00010010_11100100_11110110_0;
      patterns[4839] = 25'b00010010_11100101_11110111_0;
      patterns[4840] = 25'b00010010_11100110_11111000_0;
      patterns[4841] = 25'b00010010_11100111_11111001_0;
      patterns[4842] = 25'b00010010_11101000_11111010_0;
      patterns[4843] = 25'b00010010_11101001_11111011_0;
      patterns[4844] = 25'b00010010_11101010_11111100_0;
      patterns[4845] = 25'b00010010_11101011_11111101_0;
      patterns[4846] = 25'b00010010_11101100_11111110_0;
      patterns[4847] = 25'b00010010_11101101_11111111_0;
      patterns[4848] = 25'b00010010_11101110_00000000_1;
      patterns[4849] = 25'b00010010_11101111_00000001_1;
      patterns[4850] = 25'b00010010_11110000_00000010_1;
      patterns[4851] = 25'b00010010_11110001_00000011_1;
      patterns[4852] = 25'b00010010_11110010_00000100_1;
      patterns[4853] = 25'b00010010_11110011_00000101_1;
      patterns[4854] = 25'b00010010_11110100_00000110_1;
      patterns[4855] = 25'b00010010_11110101_00000111_1;
      patterns[4856] = 25'b00010010_11110110_00001000_1;
      patterns[4857] = 25'b00010010_11110111_00001001_1;
      patterns[4858] = 25'b00010010_11111000_00001010_1;
      patterns[4859] = 25'b00010010_11111001_00001011_1;
      patterns[4860] = 25'b00010010_11111010_00001100_1;
      patterns[4861] = 25'b00010010_11111011_00001101_1;
      patterns[4862] = 25'b00010010_11111100_00001110_1;
      patterns[4863] = 25'b00010010_11111101_00001111_1;
      patterns[4864] = 25'b00010010_11111110_00010000_1;
      patterns[4865] = 25'b00010010_11111111_00010001_1;
      patterns[4866] = 25'b00010011_00000000_00010011_0;
      patterns[4867] = 25'b00010011_00000001_00010100_0;
      patterns[4868] = 25'b00010011_00000010_00010101_0;
      patterns[4869] = 25'b00010011_00000011_00010110_0;
      patterns[4870] = 25'b00010011_00000100_00010111_0;
      patterns[4871] = 25'b00010011_00000101_00011000_0;
      patterns[4872] = 25'b00010011_00000110_00011001_0;
      patterns[4873] = 25'b00010011_00000111_00011010_0;
      patterns[4874] = 25'b00010011_00001000_00011011_0;
      patterns[4875] = 25'b00010011_00001001_00011100_0;
      patterns[4876] = 25'b00010011_00001010_00011101_0;
      patterns[4877] = 25'b00010011_00001011_00011110_0;
      patterns[4878] = 25'b00010011_00001100_00011111_0;
      patterns[4879] = 25'b00010011_00001101_00100000_0;
      patterns[4880] = 25'b00010011_00001110_00100001_0;
      patterns[4881] = 25'b00010011_00001111_00100010_0;
      patterns[4882] = 25'b00010011_00010000_00100011_0;
      patterns[4883] = 25'b00010011_00010001_00100100_0;
      patterns[4884] = 25'b00010011_00010010_00100101_0;
      patterns[4885] = 25'b00010011_00010011_00100110_0;
      patterns[4886] = 25'b00010011_00010100_00100111_0;
      patterns[4887] = 25'b00010011_00010101_00101000_0;
      patterns[4888] = 25'b00010011_00010110_00101001_0;
      patterns[4889] = 25'b00010011_00010111_00101010_0;
      patterns[4890] = 25'b00010011_00011000_00101011_0;
      patterns[4891] = 25'b00010011_00011001_00101100_0;
      patterns[4892] = 25'b00010011_00011010_00101101_0;
      patterns[4893] = 25'b00010011_00011011_00101110_0;
      patterns[4894] = 25'b00010011_00011100_00101111_0;
      patterns[4895] = 25'b00010011_00011101_00110000_0;
      patterns[4896] = 25'b00010011_00011110_00110001_0;
      patterns[4897] = 25'b00010011_00011111_00110010_0;
      patterns[4898] = 25'b00010011_00100000_00110011_0;
      patterns[4899] = 25'b00010011_00100001_00110100_0;
      patterns[4900] = 25'b00010011_00100010_00110101_0;
      patterns[4901] = 25'b00010011_00100011_00110110_0;
      patterns[4902] = 25'b00010011_00100100_00110111_0;
      patterns[4903] = 25'b00010011_00100101_00111000_0;
      patterns[4904] = 25'b00010011_00100110_00111001_0;
      patterns[4905] = 25'b00010011_00100111_00111010_0;
      patterns[4906] = 25'b00010011_00101000_00111011_0;
      patterns[4907] = 25'b00010011_00101001_00111100_0;
      patterns[4908] = 25'b00010011_00101010_00111101_0;
      patterns[4909] = 25'b00010011_00101011_00111110_0;
      patterns[4910] = 25'b00010011_00101100_00111111_0;
      patterns[4911] = 25'b00010011_00101101_01000000_0;
      patterns[4912] = 25'b00010011_00101110_01000001_0;
      patterns[4913] = 25'b00010011_00101111_01000010_0;
      patterns[4914] = 25'b00010011_00110000_01000011_0;
      patterns[4915] = 25'b00010011_00110001_01000100_0;
      patterns[4916] = 25'b00010011_00110010_01000101_0;
      patterns[4917] = 25'b00010011_00110011_01000110_0;
      patterns[4918] = 25'b00010011_00110100_01000111_0;
      patterns[4919] = 25'b00010011_00110101_01001000_0;
      patterns[4920] = 25'b00010011_00110110_01001001_0;
      patterns[4921] = 25'b00010011_00110111_01001010_0;
      patterns[4922] = 25'b00010011_00111000_01001011_0;
      patterns[4923] = 25'b00010011_00111001_01001100_0;
      patterns[4924] = 25'b00010011_00111010_01001101_0;
      patterns[4925] = 25'b00010011_00111011_01001110_0;
      patterns[4926] = 25'b00010011_00111100_01001111_0;
      patterns[4927] = 25'b00010011_00111101_01010000_0;
      patterns[4928] = 25'b00010011_00111110_01010001_0;
      patterns[4929] = 25'b00010011_00111111_01010010_0;
      patterns[4930] = 25'b00010011_01000000_01010011_0;
      patterns[4931] = 25'b00010011_01000001_01010100_0;
      patterns[4932] = 25'b00010011_01000010_01010101_0;
      patterns[4933] = 25'b00010011_01000011_01010110_0;
      patterns[4934] = 25'b00010011_01000100_01010111_0;
      patterns[4935] = 25'b00010011_01000101_01011000_0;
      patterns[4936] = 25'b00010011_01000110_01011001_0;
      patterns[4937] = 25'b00010011_01000111_01011010_0;
      patterns[4938] = 25'b00010011_01001000_01011011_0;
      patterns[4939] = 25'b00010011_01001001_01011100_0;
      patterns[4940] = 25'b00010011_01001010_01011101_0;
      patterns[4941] = 25'b00010011_01001011_01011110_0;
      patterns[4942] = 25'b00010011_01001100_01011111_0;
      patterns[4943] = 25'b00010011_01001101_01100000_0;
      patterns[4944] = 25'b00010011_01001110_01100001_0;
      patterns[4945] = 25'b00010011_01001111_01100010_0;
      patterns[4946] = 25'b00010011_01010000_01100011_0;
      patterns[4947] = 25'b00010011_01010001_01100100_0;
      patterns[4948] = 25'b00010011_01010010_01100101_0;
      patterns[4949] = 25'b00010011_01010011_01100110_0;
      patterns[4950] = 25'b00010011_01010100_01100111_0;
      patterns[4951] = 25'b00010011_01010101_01101000_0;
      patterns[4952] = 25'b00010011_01010110_01101001_0;
      patterns[4953] = 25'b00010011_01010111_01101010_0;
      patterns[4954] = 25'b00010011_01011000_01101011_0;
      patterns[4955] = 25'b00010011_01011001_01101100_0;
      patterns[4956] = 25'b00010011_01011010_01101101_0;
      patterns[4957] = 25'b00010011_01011011_01101110_0;
      patterns[4958] = 25'b00010011_01011100_01101111_0;
      patterns[4959] = 25'b00010011_01011101_01110000_0;
      patterns[4960] = 25'b00010011_01011110_01110001_0;
      patterns[4961] = 25'b00010011_01011111_01110010_0;
      patterns[4962] = 25'b00010011_01100000_01110011_0;
      patterns[4963] = 25'b00010011_01100001_01110100_0;
      patterns[4964] = 25'b00010011_01100010_01110101_0;
      patterns[4965] = 25'b00010011_01100011_01110110_0;
      patterns[4966] = 25'b00010011_01100100_01110111_0;
      patterns[4967] = 25'b00010011_01100101_01111000_0;
      patterns[4968] = 25'b00010011_01100110_01111001_0;
      patterns[4969] = 25'b00010011_01100111_01111010_0;
      patterns[4970] = 25'b00010011_01101000_01111011_0;
      patterns[4971] = 25'b00010011_01101001_01111100_0;
      patterns[4972] = 25'b00010011_01101010_01111101_0;
      patterns[4973] = 25'b00010011_01101011_01111110_0;
      patterns[4974] = 25'b00010011_01101100_01111111_0;
      patterns[4975] = 25'b00010011_01101101_10000000_0;
      patterns[4976] = 25'b00010011_01101110_10000001_0;
      patterns[4977] = 25'b00010011_01101111_10000010_0;
      patterns[4978] = 25'b00010011_01110000_10000011_0;
      patterns[4979] = 25'b00010011_01110001_10000100_0;
      patterns[4980] = 25'b00010011_01110010_10000101_0;
      patterns[4981] = 25'b00010011_01110011_10000110_0;
      patterns[4982] = 25'b00010011_01110100_10000111_0;
      patterns[4983] = 25'b00010011_01110101_10001000_0;
      patterns[4984] = 25'b00010011_01110110_10001001_0;
      patterns[4985] = 25'b00010011_01110111_10001010_0;
      patterns[4986] = 25'b00010011_01111000_10001011_0;
      patterns[4987] = 25'b00010011_01111001_10001100_0;
      patterns[4988] = 25'b00010011_01111010_10001101_0;
      patterns[4989] = 25'b00010011_01111011_10001110_0;
      patterns[4990] = 25'b00010011_01111100_10001111_0;
      patterns[4991] = 25'b00010011_01111101_10010000_0;
      patterns[4992] = 25'b00010011_01111110_10010001_0;
      patterns[4993] = 25'b00010011_01111111_10010010_0;
      patterns[4994] = 25'b00010011_10000000_10010011_0;
      patterns[4995] = 25'b00010011_10000001_10010100_0;
      patterns[4996] = 25'b00010011_10000010_10010101_0;
      patterns[4997] = 25'b00010011_10000011_10010110_0;
      patterns[4998] = 25'b00010011_10000100_10010111_0;
      patterns[4999] = 25'b00010011_10000101_10011000_0;
      patterns[5000] = 25'b00010011_10000110_10011001_0;
      patterns[5001] = 25'b00010011_10000111_10011010_0;
      patterns[5002] = 25'b00010011_10001000_10011011_0;
      patterns[5003] = 25'b00010011_10001001_10011100_0;
      patterns[5004] = 25'b00010011_10001010_10011101_0;
      patterns[5005] = 25'b00010011_10001011_10011110_0;
      patterns[5006] = 25'b00010011_10001100_10011111_0;
      patterns[5007] = 25'b00010011_10001101_10100000_0;
      patterns[5008] = 25'b00010011_10001110_10100001_0;
      patterns[5009] = 25'b00010011_10001111_10100010_0;
      patterns[5010] = 25'b00010011_10010000_10100011_0;
      patterns[5011] = 25'b00010011_10010001_10100100_0;
      patterns[5012] = 25'b00010011_10010010_10100101_0;
      patterns[5013] = 25'b00010011_10010011_10100110_0;
      patterns[5014] = 25'b00010011_10010100_10100111_0;
      patterns[5015] = 25'b00010011_10010101_10101000_0;
      patterns[5016] = 25'b00010011_10010110_10101001_0;
      patterns[5017] = 25'b00010011_10010111_10101010_0;
      patterns[5018] = 25'b00010011_10011000_10101011_0;
      patterns[5019] = 25'b00010011_10011001_10101100_0;
      patterns[5020] = 25'b00010011_10011010_10101101_0;
      patterns[5021] = 25'b00010011_10011011_10101110_0;
      patterns[5022] = 25'b00010011_10011100_10101111_0;
      patterns[5023] = 25'b00010011_10011101_10110000_0;
      patterns[5024] = 25'b00010011_10011110_10110001_0;
      patterns[5025] = 25'b00010011_10011111_10110010_0;
      patterns[5026] = 25'b00010011_10100000_10110011_0;
      patterns[5027] = 25'b00010011_10100001_10110100_0;
      patterns[5028] = 25'b00010011_10100010_10110101_0;
      patterns[5029] = 25'b00010011_10100011_10110110_0;
      patterns[5030] = 25'b00010011_10100100_10110111_0;
      patterns[5031] = 25'b00010011_10100101_10111000_0;
      patterns[5032] = 25'b00010011_10100110_10111001_0;
      patterns[5033] = 25'b00010011_10100111_10111010_0;
      patterns[5034] = 25'b00010011_10101000_10111011_0;
      patterns[5035] = 25'b00010011_10101001_10111100_0;
      patterns[5036] = 25'b00010011_10101010_10111101_0;
      patterns[5037] = 25'b00010011_10101011_10111110_0;
      patterns[5038] = 25'b00010011_10101100_10111111_0;
      patterns[5039] = 25'b00010011_10101101_11000000_0;
      patterns[5040] = 25'b00010011_10101110_11000001_0;
      patterns[5041] = 25'b00010011_10101111_11000010_0;
      patterns[5042] = 25'b00010011_10110000_11000011_0;
      patterns[5043] = 25'b00010011_10110001_11000100_0;
      patterns[5044] = 25'b00010011_10110010_11000101_0;
      patterns[5045] = 25'b00010011_10110011_11000110_0;
      patterns[5046] = 25'b00010011_10110100_11000111_0;
      patterns[5047] = 25'b00010011_10110101_11001000_0;
      patterns[5048] = 25'b00010011_10110110_11001001_0;
      patterns[5049] = 25'b00010011_10110111_11001010_0;
      patterns[5050] = 25'b00010011_10111000_11001011_0;
      patterns[5051] = 25'b00010011_10111001_11001100_0;
      patterns[5052] = 25'b00010011_10111010_11001101_0;
      patterns[5053] = 25'b00010011_10111011_11001110_0;
      patterns[5054] = 25'b00010011_10111100_11001111_0;
      patterns[5055] = 25'b00010011_10111101_11010000_0;
      patterns[5056] = 25'b00010011_10111110_11010001_0;
      patterns[5057] = 25'b00010011_10111111_11010010_0;
      patterns[5058] = 25'b00010011_11000000_11010011_0;
      patterns[5059] = 25'b00010011_11000001_11010100_0;
      patterns[5060] = 25'b00010011_11000010_11010101_0;
      patterns[5061] = 25'b00010011_11000011_11010110_0;
      patterns[5062] = 25'b00010011_11000100_11010111_0;
      patterns[5063] = 25'b00010011_11000101_11011000_0;
      patterns[5064] = 25'b00010011_11000110_11011001_0;
      patterns[5065] = 25'b00010011_11000111_11011010_0;
      patterns[5066] = 25'b00010011_11001000_11011011_0;
      patterns[5067] = 25'b00010011_11001001_11011100_0;
      patterns[5068] = 25'b00010011_11001010_11011101_0;
      patterns[5069] = 25'b00010011_11001011_11011110_0;
      patterns[5070] = 25'b00010011_11001100_11011111_0;
      patterns[5071] = 25'b00010011_11001101_11100000_0;
      patterns[5072] = 25'b00010011_11001110_11100001_0;
      patterns[5073] = 25'b00010011_11001111_11100010_0;
      patterns[5074] = 25'b00010011_11010000_11100011_0;
      patterns[5075] = 25'b00010011_11010001_11100100_0;
      patterns[5076] = 25'b00010011_11010010_11100101_0;
      patterns[5077] = 25'b00010011_11010011_11100110_0;
      patterns[5078] = 25'b00010011_11010100_11100111_0;
      patterns[5079] = 25'b00010011_11010101_11101000_0;
      patterns[5080] = 25'b00010011_11010110_11101001_0;
      patterns[5081] = 25'b00010011_11010111_11101010_0;
      patterns[5082] = 25'b00010011_11011000_11101011_0;
      patterns[5083] = 25'b00010011_11011001_11101100_0;
      patterns[5084] = 25'b00010011_11011010_11101101_0;
      patterns[5085] = 25'b00010011_11011011_11101110_0;
      patterns[5086] = 25'b00010011_11011100_11101111_0;
      patterns[5087] = 25'b00010011_11011101_11110000_0;
      patterns[5088] = 25'b00010011_11011110_11110001_0;
      patterns[5089] = 25'b00010011_11011111_11110010_0;
      patterns[5090] = 25'b00010011_11100000_11110011_0;
      patterns[5091] = 25'b00010011_11100001_11110100_0;
      patterns[5092] = 25'b00010011_11100010_11110101_0;
      patterns[5093] = 25'b00010011_11100011_11110110_0;
      patterns[5094] = 25'b00010011_11100100_11110111_0;
      patterns[5095] = 25'b00010011_11100101_11111000_0;
      patterns[5096] = 25'b00010011_11100110_11111001_0;
      patterns[5097] = 25'b00010011_11100111_11111010_0;
      patterns[5098] = 25'b00010011_11101000_11111011_0;
      patterns[5099] = 25'b00010011_11101001_11111100_0;
      patterns[5100] = 25'b00010011_11101010_11111101_0;
      patterns[5101] = 25'b00010011_11101011_11111110_0;
      patterns[5102] = 25'b00010011_11101100_11111111_0;
      patterns[5103] = 25'b00010011_11101101_00000000_1;
      patterns[5104] = 25'b00010011_11101110_00000001_1;
      patterns[5105] = 25'b00010011_11101111_00000010_1;
      patterns[5106] = 25'b00010011_11110000_00000011_1;
      patterns[5107] = 25'b00010011_11110001_00000100_1;
      patterns[5108] = 25'b00010011_11110010_00000101_1;
      patterns[5109] = 25'b00010011_11110011_00000110_1;
      patterns[5110] = 25'b00010011_11110100_00000111_1;
      patterns[5111] = 25'b00010011_11110101_00001000_1;
      patterns[5112] = 25'b00010011_11110110_00001001_1;
      patterns[5113] = 25'b00010011_11110111_00001010_1;
      patterns[5114] = 25'b00010011_11111000_00001011_1;
      patterns[5115] = 25'b00010011_11111001_00001100_1;
      patterns[5116] = 25'b00010011_11111010_00001101_1;
      patterns[5117] = 25'b00010011_11111011_00001110_1;
      patterns[5118] = 25'b00010011_11111100_00001111_1;
      patterns[5119] = 25'b00010011_11111101_00010000_1;
      patterns[5120] = 25'b00010011_11111110_00010001_1;
      patterns[5121] = 25'b00010011_11111111_00010010_1;
      patterns[5122] = 25'b00010100_00000000_00010100_0;
      patterns[5123] = 25'b00010100_00000001_00010101_0;
      patterns[5124] = 25'b00010100_00000010_00010110_0;
      patterns[5125] = 25'b00010100_00000011_00010111_0;
      patterns[5126] = 25'b00010100_00000100_00011000_0;
      patterns[5127] = 25'b00010100_00000101_00011001_0;
      patterns[5128] = 25'b00010100_00000110_00011010_0;
      patterns[5129] = 25'b00010100_00000111_00011011_0;
      patterns[5130] = 25'b00010100_00001000_00011100_0;
      patterns[5131] = 25'b00010100_00001001_00011101_0;
      patterns[5132] = 25'b00010100_00001010_00011110_0;
      patterns[5133] = 25'b00010100_00001011_00011111_0;
      patterns[5134] = 25'b00010100_00001100_00100000_0;
      patterns[5135] = 25'b00010100_00001101_00100001_0;
      patterns[5136] = 25'b00010100_00001110_00100010_0;
      patterns[5137] = 25'b00010100_00001111_00100011_0;
      patterns[5138] = 25'b00010100_00010000_00100100_0;
      patterns[5139] = 25'b00010100_00010001_00100101_0;
      patterns[5140] = 25'b00010100_00010010_00100110_0;
      patterns[5141] = 25'b00010100_00010011_00100111_0;
      patterns[5142] = 25'b00010100_00010100_00101000_0;
      patterns[5143] = 25'b00010100_00010101_00101001_0;
      patterns[5144] = 25'b00010100_00010110_00101010_0;
      patterns[5145] = 25'b00010100_00010111_00101011_0;
      patterns[5146] = 25'b00010100_00011000_00101100_0;
      patterns[5147] = 25'b00010100_00011001_00101101_0;
      patterns[5148] = 25'b00010100_00011010_00101110_0;
      patterns[5149] = 25'b00010100_00011011_00101111_0;
      patterns[5150] = 25'b00010100_00011100_00110000_0;
      patterns[5151] = 25'b00010100_00011101_00110001_0;
      patterns[5152] = 25'b00010100_00011110_00110010_0;
      patterns[5153] = 25'b00010100_00011111_00110011_0;
      patterns[5154] = 25'b00010100_00100000_00110100_0;
      patterns[5155] = 25'b00010100_00100001_00110101_0;
      patterns[5156] = 25'b00010100_00100010_00110110_0;
      patterns[5157] = 25'b00010100_00100011_00110111_0;
      patterns[5158] = 25'b00010100_00100100_00111000_0;
      patterns[5159] = 25'b00010100_00100101_00111001_0;
      patterns[5160] = 25'b00010100_00100110_00111010_0;
      patterns[5161] = 25'b00010100_00100111_00111011_0;
      patterns[5162] = 25'b00010100_00101000_00111100_0;
      patterns[5163] = 25'b00010100_00101001_00111101_0;
      patterns[5164] = 25'b00010100_00101010_00111110_0;
      patterns[5165] = 25'b00010100_00101011_00111111_0;
      patterns[5166] = 25'b00010100_00101100_01000000_0;
      patterns[5167] = 25'b00010100_00101101_01000001_0;
      patterns[5168] = 25'b00010100_00101110_01000010_0;
      patterns[5169] = 25'b00010100_00101111_01000011_0;
      patterns[5170] = 25'b00010100_00110000_01000100_0;
      patterns[5171] = 25'b00010100_00110001_01000101_0;
      patterns[5172] = 25'b00010100_00110010_01000110_0;
      patterns[5173] = 25'b00010100_00110011_01000111_0;
      patterns[5174] = 25'b00010100_00110100_01001000_0;
      patterns[5175] = 25'b00010100_00110101_01001001_0;
      patterns[5176] = 25'b00010100_00110110_01001010_0;
      patterns[5177] = 25'b00010100_00110111_01001011_0;
      patterns[5178] = 25'b00010100_00111000_01001100_0;
      patterns[5179] = 25'b00010100_00111001_01001101_0;
      patterns[5180] = 25'b00010100_00111010_01001110_0;
      patterns[5181] = 25'b00010100_00111011_01001111_0;
      patterns[5182] = 25'b00010100_00111100_01010000_0;
      patterns[5183] = 25'b00010100_00111101_01010001_0;
      patterns[5184] = 25'b00010100_00111110_01010010_0;
      patterns[5185] = 25'b00010100_00111111_01010011_0;
      patterns[5186] = 25'b00010100_01000000_01010100_0;
      patterns[5187] = 25'b00010100_01000001_01010101_0;
      patterns[5188] = 25'b00010100_01000010_01010110_0;
      patterns[5189] = 25'b00010100_01000011_01010111_0;
      patterns[5190] = 25'b00010100_01000100_01011000_0;
      patterns[5191] = 25'b00010100_01000101_01011001_0;
      patterns[5192] = 25'b00010100_01000110_01011010_0;
      patterns[5193] = 25'b00010100_01000111_01011011_0;
      patterns[5194] = 25'b00010100_01001000_01011100_0;
      patterns[5195] = 25'b00010100_01001001_01011101_0;
      patterns[5196] = 25'b00010100_01001010_01011110_0;
      patterns[5197] = 25'b00010100_01001011_01011111_0;
      patterns[5198] = 25'b00010100_01001100_01100000_0;
      patterns[5199] = 25'b00010100_01001101_01100001_0;
      patterns[5200] = 25'b00010100_01001110_01100010_0;
      patterns[5201] = 25'b00010100_01001111_01100011_0;
      patterns[5202] = 25'b00010100_01010000_01100100_0;
      patterns[5203] = 25'b00010100_01010001_01100101_0;
      patterns[5204] = 25'b00010100_01010010_01100110_0;
      patterns[5205] = 25'b00010100_01010011_01100111_0;
      patterns[5206] = 25'b00010100_01010100_01101000_0;
      patterns[5207] = 25'b00010100_01010101_01101001_0;
      patterns[5208] = 25'b00010100_01010110_01101010_0;
      patterns[5209] = 25'b00010100_01010111_01101011_0;
      patterns[5210] = 25'b00010100_01011000_01101100_0;
      patterns[5211] = 25'b00010100_01011001_01101101_0;
      patterns[5212] = 25'b00010100_01011010_01101110_0;
      patterns[5213] = 25'b00010100_01011011_01101111_0;
      patterns[5214] = 25'b00010100_01011100_01110000_0;
      patterns[5215] = 25'b00010100_01011101_01110001_0;
      patterns[5216] = 25'b00010100_01011110_01110010_0;
      patterns[5217] = 25'b00010100_01011111_01110011_0;
      patterns[5218] = 25'b00010100_01100000_01110100_0;
      patterns[5219] = 25'b00010100_01100001_01110101_0;
      patterns[5220] = 25'b00010100_01100010_01110110_0;
      patterns[5221] = 25'b00010100_01100011_01110111_0;
      patterns[5222] = 25'b00010100_01100100_01111000_0;
      patterns[5223] = 25'b00010100_01100101_01111001_0;
      patterns[5224] = 25'b00010100_01100110_01111010_0;
      patterns[5225] = 25'b00010100_01100111_01111011_0;
      patterns[5226] = 25'b00010100_01101000_01111100_0;
      patterns[5227] = 25'b00010100_01101001_01111101_0;
      patterns[5228] = 25'b00010100_01101010_01111110_0;
      patterns[5229] = 25'b00010100_01101011_01111111_0;
      patterns[5230] = 25'b00010100_01101100_10000000_0;
      patterns[5231] = 25'b00010100_01101101_10000001_0;
      patterns[5232] = 25'b00010100_01101110_10000010_0;
      patterns[5233] = 25'b00010100_01101111_10000011_0;
      patterns[5234] = 25'b00010100_01110000_10000100_0;
      patterns[5235] = 25'b00010100_01110001_10000101_0;
      patterns[5236] = 25'b00010100_01110010_10000110_0;
      patterns[5237] = 25'b00010100_01110011_10000111_0;
      patterns[5238] = 25'b00010100_01110100_10001000_0;
      patterns[5239] = 25'b00010100_01110101_10001001_0;
      patterns[5240] = 25'b00010100_01110110_10001010_0;
      patterns[5241] = 25'b00010100_01110111_10001011_0;
      patterns[5242] = 25'b00010100_01111000_10001100_0;
      patterns[5243] = 25'b00010100_01111001_10001101_0;
      patterns[5244] = 25'b00010100_01111010_10001110_0;
      patterns[5245] = 25'b00010100_01111011_10001111_0;
      patterns[5246] = 25'b00010100_01111100_10010000_0;
      patterns[5247] = 25'b00010100_01111101_10010001_0;
      patterns[5248] = 25'b00010100_01111110_10010010_0;
      patterns[5249] = 25'b00010100_01111111_10010011_0;
      patterns[5250] = 25'b00010100_10000000_10010100_0;
      patterns[5251] = 25'b00010100_10000001_10010101_0;
      patterns[5252] = 25'b00010100_10000010_10010110_0;
      patterns[5253] = 25'b00010100_10000011_10010111_0;
      patterns[5254] = 25'b00010100_10000100_10011000_0;
      patterns[5255] = 25'b00010100_10000101_10011001_0;
      patterns[5256] = 25'b00010100_10000110_10011010_0;
      patterns[5257] = 25'b00010100_10000111_10011011_0;
      patterns[5258] = 25'b00010100_10001000_10011100_0;
      patterns[5259] = 25'b00010100_10001001_10011101_0;
      patterns[5260] = 25'b00010100_10001010_10011110_0;
      patterns[5261] = 25'b00010100_10001011_10011111_0;
      patterns[5262] = 25'b00010100_10001100_10100000_0;
      patterns[5263] = 25'b00010100_10001101_10100001_0;
      patterns[5264] = 25'b00010100_10001110_10100010_0;
      patterns[5265] = 25'b00010100_10001111_10100011_0;
      patterns[5266] = 25'b00010100_10010000_10100100_0;
      patterns[5267] = 25'b00010100_10010001_10100101_0;
      patterns[5268] = 25'b00010100_10010010_10100110_0;
      patterns[5269] = 25'b00010100_10010011_10100111_0;
      patterns[5270] = 25'b00010100_10010100_10101000_0;
      patterns[5271] = 25'b00010100_10010101_10101001_0;
      patterns[5272] = 25'b00010100_10010110_10101010_0;
      patterns[5273] = 25'b00010100_10010111_10101011_0;
      patterns[5274] = 25'b00010100_10011000_10101100_0;
      patterns[5275] = 25'b00010100_10011001_10101101_0;
      patterns[5276] = 25'b00010100_10011010_10101110_0;
      patterns[5277] = 25'b00010100_10011011_10101111_0;
      patterns[5278] = 25'b00010100_10011100_10110000_0;
      patterns[5279] = 25'b00010100_10011101_10110001_0;
      patterns[5280] = 25'b00010100_10011110_10110010_0;
      patterns[5281] = 25'b00010100_10011111_10110011_0;
      patterns[5282] = 25'b00010100_10100000_10110100_0;
      patterns[5283] = 25'b00010100_10100001_10110101_0;
      patterns[5284] = 25'b00010100_10100010_10110110_0;
      patterns[5285] = 25'b00010100_10100011_10110111_0;
      patterns[5286] = 25'b00010100_10100100_10111000_0;
      patterns[5287] = 25'b00010100_10100101_10111001_0;
      patterns[5288] = 25'b00010100_10100110_10111010_0;
      patterns[5289] = 25'b00010100_10100111_10111011_0;
      patterns[5290] = 25'b00010100_10101000_10111100_0;
      patterns[5291] = 25'b00010100_10101001_10111101_0;
      patterns[5292] = 25'b00010100_10101010_10111110_0;
      patterns[5293] = 25'b00010100_10101011_10111111_0;
      patterns[5294] = 25'b00010100_10101100_11000000_0;
      patterns[5295] = 25'b00010100_10101101_11000001_0;
      patterns[5296] = 25'b00010100_10101110_11000010_0;
      patterns[5297] = 25'b00010100_10101111_11000011_0;
      patterns[5298] = 25'b00010100_10110000_11000100_0;
      patterns[5299] = 25'b00010100_10110001_11000101_0;
      patterns[5300] = 25'b00010100_10110010_11000110_0;
      patterns[5301] = 25'b00010100_10110011_11000111_0;
      patterns[5302] = 25'b00010100_10110100_11001000_0;
      patterns[5303] = 25'b00010100_10110101_11001001_0;
      patterns[5304] = 25'b00010100_10110110_11001010_0;
      patterns[5305] = 25'b00010100_10110111_11001011_0;
      patterns[5306] = 25'b00010100_10111000_11001100_0;
      patterns[5307] = 25'b00010100_10111001_11001101_0;
      patterns[5308] = 25'b00010100_10111010_11001110_0;
      patterns[5309] = 25'b00010100_10111011_11001111_0;
      patterns[5310] = 25'b00010100_10111100_11010000_0;
      patterns[5311] = 25'b00010100_10111101_11010001_0;
      patterns[5312] = 25'b00010100_10111110_11010010_0;
      patterns[5313] = 25'b00010100_10111111_11010011_0;
      patterns[5314] = 25'b00010100_11000000_11010100_0;
      patterns[5315] = 25'b00010100_11000001_11010101_0;
      patterns[5316] = 25'b00010100_11000010_11010110_0;
      patterns[5317] = 25'b00010100_11000011_11010111_0;
      patterns[5318] = 25'b00010100_11000100_11011000_0;
      patterns[5319] = 25'b00010100_11000101_11011001_0;
      patterns[5320] = 25'b00010100_11000110_11011010_0;
      patterns[5321] = 25'b00010100_11000111_11011011_0;
      patterns[5322] = 25'b00010100_11001000_11011100_0;
      patterns[5323] = 25'b00010100_11001001_11011101_0;
      patterns[5324] = 25'b00010100_11001010_11011110_0;
      patterns[5325] = 25'b00010100_11001011_11011111_0;
      patterns[5326] = 25'b00010100_11001100_11100000_0;
      patterns[5327] = 25'b00010100_11001101_11100001_0;
      patterns[5328] = 25'b00010100_11001110_11100010_0;
      patterns[5329] = 25'b00010100_11001111_11100011_0;
      patterns[5330] = 25'b00010100_11010000_11100100_0;
      patterns[5331] = 25'b00010100_11010001_11100101_0;
      patterns[5332] = 25'b00010100_11010010_11100110_0;
      patterns[5333] = 25'b00010100_11010011_11100111_0;
      patterns[5334] = 25'b00010100_11010100_11101000_0;
      patterns[5335] = 25'b00010100_11010101_11101001_0;
      patterns[5336] = 25'b00010100_11010110_11101010_0;
      patterns[5337] = 25'b00010100_11010111_11101011_0;
      patterns[5338] = 25'b00010100_11011000_11101100_0;
      patterns[5339] = 25'b00010100_11011001_11101101_0;
      patterns[5340] = 25'b00010100_11011010_11101110_0;
      patterns[5341] = 25'b00010100_11011011_11101111_0;
      patterns[5342] = 25'b00010100_11011100_11110000_0;
      patterns[5343] = 25'b00010100_11011101_11110001_0;
      patterns[5344] = 25'b00010100_11011110_11110010_0;
      patterns[5345] = 25'b00010100_11011111_11110011_0;
      patterns[5346] = 25'b00010100_11100000_11110100_0;
      patterns[5347] = 25'b00010100_11100001_11110101_0;
      patterns[5348] = 25'b00010100_11100010_11110110_0;
      patterns[5349] = 25'b00010100_11100011_11110111_0;
      patterns[5350] = 25'b00010100_11100100_11111000_0;
      patterns[5351] = 25'b00010100_11100101_11111001_0;
      patterns[5352] = 25'b00010100_11100110_11111010_0;
      patterns[5353] = 25'b00010100_11100111_11111011_0;
      patterns[5354] = 25'b00010100_11101000_11111100_0;
      patterns[5355] = 25'b00010100_11101001_11111101_0;
      patterns[5356] = 25'b00010100_11101010_11111110_0;
      patterns[5357] = 25'b00010100_11101011_11111111_0;
      patterns[5358] = 25'b00010100_11101100_00000000_1;
      patterns[5359] = 25'b00010100_11101101_00000001_1;
      patterns[5360] = 25'b00010100_11101110_00000010_1;
      patterns[5361] = 25'b00010100_11101111_00000011_1;
      patterns[5362] = 25'b00010100_11110000_00000100_1;
      patterns[5363] = 25'b00010100_11110001_00000101_1;
      patterns[5364] = 25'b00010100_11110010_00000110_1;
      patterns[5365] = 25'b00010100_11110011_00000111_1;
      patterns[5366] = 25'b00010100_11110100_00001000_1;
      patterns[5367] = 25'b00010100_11110101_00001001_1;
      patterns[5368] = 25'b00010100_11110110_00001010_1;
      patterns[5369] = 25'b00010100_11110111_00001011_1;
      patterns[5370] = 25'b00010100_11111000_00001100_1;
      patterns[5371] = 25'b00010100_11111001_00001101_1;
      patterns[5372] = 25'b00010100_11111010_00001110_1;
      patterns[5373] = 25'b00010100_11111011_00001111_1;
      patterns[5374] = 25'b00010100_11111100_00010000_1;
      patterns[5375] = 25'b00010100_11111101_00010001_1;
      patterns[5376] = 25'b00010100_11111110_00010010_1;
      patterns[5377] = 25'b00010100_11111111_00010011_1;
      patterns[5378] = 25'b00010101_00000000_00010101_0;
      patterns[5379] = 25'b00010101_00000001_00010110_0;
      patterns[5380] = 25'b00010101_00000010_00010111_0;
      patterns[5381] = 25'b00010101_00000011_00011000_0;
      patterns[5382] = 25'b00010101_00000100_00011001_0;
      patterns[5383] = 25'b00010101_00000101_00011010_0;
      patterns[5384] = 25'b00010101_00000110_00011011_0;
      patterns[5385] = 25'b00010101_00000111_00011100_0;
      patterns[5386] = 25'b00010101_00001000_00011101_0;
      patterns[5387] = 25'b00010101_00001001_00011110_0;
      patterns[5388] = 25'b00010101_00001010_00011111_0;
      patterns[5389] = 25'b00010101_00001011_00100000_0;
      patterns[5390] = 25'b00010101_00001100_00100001_0;
      patterns[5391] = 25'b00010101_00001101_00100010_0;
      patterns[5392] = 25'b00010101_00001110_00100011_0;
      patterns[5393] = 25'b00010101_00001111_00100100_0;
      patterns[5394] = 25'b00010101_00010000_00100101_0;
      patterns[5395] = 25'b00010101_00010001_00100110_0;
      patterns[5396] = 25'b00010101_00010010_00100111_0;
      patterns[5397] = 25'b00010101_00010011_00101000_0;
      patterns[5398] = 25'b00010101_00010100_00101001_0;
      patterns[5399] = 25'b00010101_00010101_00101010_0;
      patterns[5400] = 25'b00010101_00010110_00101011_0;
      patterns[5401] = 25'b00010101_00010111_00101100_0;
      patterns[5402] = 25'b00010101_00011000_00101101_0;
      patterns[5403] = 25'b00010101_00011001_00101110_0;
      patterns[5404] = 25'b00010101_00011010_00101111_0;
      patterns[5405] = 25'b00010101_00011011_00110000_0;
      patterns[5406] = 25'b00010101_00011100_00110001_0;
      patterns[5407] = 25'b00010101_00011101_00110010_0;
      patterns[5408] = 25'b00010101_00011110_00110011_0;
      patterns[5409] = 25'b00010101_00011111_00110100_0;
      patterns[5410] = 25'b00010101_00100000_00110101_0;
      patterns[5411] = 25'b00010101_00100001_00110110_0;
      patterns[5412] = 25'b00010101_00100010_00110111_0;
      patterns[5413] = 25'b00010101_00100011_00111000_0;
      patterns[5414] = 25'b00010101_00100100_00111001_0;
      patterns[5415] = 25'b00010101_00100101_00111010_0;
      patterns[5416] = 25'b00010101_00100110_00111011_0;
      patterns[5417] = 25'b00010101_00100111_00111100_0;
      patterns[5418] = 25'b00010101_00101000_00111101_0;
      patterns[5419] = 25'b00010101_00101001_00111110_0;
      patterns[5420] = 25'b00010101_00101010_00111111_0;
      patterns[5421] = 25'b00010101_00101011_01000000_0;
      patterns[5422] = 25'b00010101_00101100_01000001_0;
      patterns[5423] = 25'b00010101_00101101_01000010_0;
      patterns[5424] = 25'b00010101_00101110_01000011_0;
      patterns[5425] = 25'b00010101_00101111_01000100_0;
      patterns[5426] = 25'b00010101_00110000_01000101_0;
      patterns[5427] = 25'b00010101_00110001_01000110_0;
      patterns[5428] = 25'b00010101_00110010_01000111_0;
      patterns[5429] = 25'b00010101_00110011_01001000_0;
      patterns[5430] = 25'b00010101_00110100_01001001_0;
      patterns[5431] = 25'b00010101_00110101_01001010_0;
      patterns[5432] = 25'b00010101_00110110_01001011_0;
      patterns[5433] = 25'b00010101_00110111_01001100_0;
      patterns[5434] = 25'b00010101_00111000_01001101_0;
      patterns[5435] = 25'b00010101_00111001_01001110_0;
      patterns[5436] = 25'b00010101_00111010_01001111_0;
      patterns[5437] = 25'b00010101_00111011_01010000_0;
      patterns[5438] = 25'b00010101_00111100_01010001_0;
      patterns[5439] = 25'b00010101_00111101_01010010_0;
      patterns[5440] = 25'b00010101_00111110_01010011_0;
      patterns[5441] = 25'b00010101_00111111_01010100_0;
      patterns[5442] = 25'b00010101_01000000_01010101_0;
      patterns[5443] = 25'b00010101_01000001_01010110_0;
      patterns[5444] = 25'b00010101_01000010_01010111_0;
      patterns[5445] = 25'b00010101_01000011_01011000_0;
      patterns[5446] = 25'b00010101_01000100_01011001_0;
      patterns[5447] = 25'b00010101_01000101_01011010_0;
      patterns[5448] = 25'b00010101_01000110_01011011_0;
      patterns[5449] = 25'b00010101_01000111_01011100_0;
      patterns[5450] = 25'b00010101_01001000_01011101_0;
      patterns[5451] = 25'b00010101_01001001_01011110_0;
      patterns[5452] = 25'b00010101_01001010_01011111_0;
      patterns[5453] = 25'b00010101_01001011_01100000_0;
      patterns[5454] = 25'b00010101_01001100_01100001_0;
      patterns[5455] = 25'b00010101_01001101_01100010_0;
      patterns[5456] = 25'b00010101_01001110_01100011_0;
      patterns[5457] = 25'b00010101_01001111_01100100_0;
      patterns[5458] = 25'b00010101_01010000_01100101_0;
      patterns[5459] = 25'b00010101_01010001_01100110_0;
      patterns[5460] = 25'b00010101_01010010_01100111_0;
      patterns[5461] = 25'b00010101_01010011_01101000_0;
      patterns[5462] = 25'b00010101_01010100_01101001_0;
      patterns[5463] = 25'b00010101_01010101_01101010_0;
      patterns[5464] = 25'b00010101_01010110_01101011_0;
      patterns[5465] = 25'b00010101_01010111_01101100_0;
      patterns[5466] = 25'b00010101_01011000_01101101_0;
      patterns[5467] = 25'b00010101_01011001_01101110_0;
      patterns[5468] = 25'b00010101_01011010_01101111_0;
      patterns[5469] = 25'b00010101_01011011_01110000_0;
      patterns[5470] = 25'b00010101_01011100_01110001_0;
      patterns[5471] = 25'b00010101_01011101_01110010_0;
      patterns[5472] = 25'b00010101_01011110_01110011_0;
      patterns[5473] = 25'b00010101_01011111_01110100_0;
      patterns[5474] = 25'b00010101_01100000_01110101_0;
      patterns[5475] = 25'b00010101_01100001_01110110_0;
      patterns[5476] = 25'b00010101_01100010_01110111_0;
      patterns[5477] = 25'b00010101_01100011_01111000_0;
      patterns[5478] = 25'b00010101_01100100_01111001_0;
      patterns[5479] = 25'b00010101_01100101_01111010_0;
      patterns[5480] = 25'b00010101_01100110_01111011_0;
      patterns[5481] = 25'b00010101_01100111_01111100_0;
      patterns[5482] = 25'b00010101_01101000_01111101_0;
      patterns[5483] = 25'b00010101_01101001_01111110_0;
      patterns[5484] = 25'b00010101_01101010_01111111_0;
      patterns[5485] = 25'b00010101_01101011_10000000_0;
      patterns[5486] = 25'b00010101_01101100_10000001_0;
      patterns[5487] = 25'b00010101_01101101_10000010_0;
      patterns[5488] = 25'b00010101_01101110_10000011_0;
      patterns[5489] = 25'b00010101_01101111_10000100_0;
      patterns[5490] = 25'b00010101_01110000_10000101_0;
      patterns[5491] = 25'b00010101_01110001_10000110_0;
      patterns[5492] = 25'b00010101_01110010_10000111_0;
      patterns[5493] = 25'b00010101_01110011_10001000_0;
      patterns[5494] = 25'b00010101_01110100_10001001_0;
      patterns[5495] = 25'b00010101_01110101_10001010_0;
      patterns[5496] = 25'b00010101_01110110_10001011_0;
      patterns[5497] = 25'b00010101_01110111_10001100_0;
      patterns[5498] = 25'b00010101_01111000_10001101_0;
      patterns[5499] = 25'b00010101_01111001_10001110_0;
      patterns[5500] = 25'b00010101_01111010_10001111_0;
      patterns[5501] = 25'b00010101_01111011_10010000_0;
      patterns[5502] = 25'b00010101_01111100_10010001_0;
      patterns[5503] = 25'b00010101_01111101_10010010_0;
      patterns[5504] = 25'b00010101_01111110_10010011_0;
      patterns[5505] = 25'b00010101_01111111_10010100_0;
      patterns[5506] = 25'b00010101_10000000_10010101_0;
      patterns[5507] = 25'b00010101_10000001_10010110_0;
      patterns[5508] = 25'b00010101_10000010_10010111_0;
      patterns[5509] = 25'b00010101_10000011_10011000_0;
      patterns[5510] = 25'b00010101_10000100_10011001_0;
      patterns[5511] = 25'b00010101_10000101_10011010_0;
      patterns[5512] = 25'b00010101_10000110_10011011_0;
      patterns[5513] = 25'b00010101_10000111_10011100_0;
      patterns[5514] = 25'b00010101_10001000_10011101_0;
      patterns[5515] = 25'b00010101_10001001_10011110_0;
      patterns[5516] = 25'b00010101_10001010_10011111_0;
      patterns[5517] = 25'b00010101_10001011_10100000_0;
      patterns[5518] = 25'b00010101_10001100_10100001_0;
      patterns[5519] = 25'b00010101_10001101_10100010_0;
      patterns[5520] = 25'b00010101_10001110_10100011_0;
      patterns[5521] = 25'b00010101_10001111_10100100_0;
      patterns[5522] = 25'b00010101_10010000_10100101_0;
      patterns[5523] = 25'b00010101_10010001_10100110_0;
      patterns[5524] = 25'b00010101_10010010_10100111_0;
      patterns[5525] = 25'b00010101_10010011_10101000_0;
      patterns[5526] = 25'b00010101_10010100_10101001_0;
      patterns[5527] = 25'b00010101_10010101_10101010_0;
      patterns[5528] = 25'b00010101_10010110_10101011_0;
      patterns[5529] = 25'b00010101_10010111_10101100_0;
      patterns[5530] = 25'b00010101_10011000_10101101_0;
      patterns[5531] = 25'b00010101_10011001_10101110_0;
      patterns[5532] = 25'b00010101_10011010_10101111_0;
      patterns[5533] = 25'b00010101_10011011_10110000_0;
      patterns[5534] = 25'b00010101_10011100_10110001_0;
      patterns[5535] = 25'b00010101_10011101_10110010_0;
      patterns[5536] = 25'b00010101_10011110_10110011_0;
      patterns[5537] = 25'b00010101_10011111_10110100_0;
      patterns[5538] = 25'b00010101_10100000_10110101_0;
      patterns[5539] = 25'b00010101_10100001_10110110_0;
      patterns[5540] = 25'b00010101_10100010_10110111_0;
      patterns[5541] = 25'b00010101_10100011_10111000_0;
      patterns[5542] = 25'b00010101_10100100_10111001_0;
      patterns[5543] = 25'b00010101_10100101_10111010_0;
      patterns[5544] = 25'b00010101_10100110_10111011_0;
      patterns[5545] = 25'b00010101_10100111_10111100_0;
      patterns[5546] = 25'b00010101_10101000_10111101_0;
      patterns[5547] = 25'b00010101_10101001_10111110_0;
      patterns[5548] = 25'b00010101_10101010_10111111_0;
      patterns[5549] = 25'b00010101_10101011_11000000_0;
      patterns[5550] = 25'b00010101_10101100_11000001_0;
      patterns[5551] = 25'b00010101_10101101_11000010_0;
      patterns[5552] = 25'b00010101_10101110_11000011_0;
      patterns[5553] = 25'b00010101_10101111_11000100_0;
      patterns[5554] = 25'b00010101_10110000_11000101_0;
      patterns[5555] = 25'b00010101_10110001_11000110_0;
      patterns[5556] = 25'b00010101_10110010_11000111_0;
      patterns[5557] = 25'b00010101_10110011_11001000_0;
      patterns[5558] = 25'b00010101_10110100_11001001_0;
      patterns[5559] = 25'b00010101_10110101_11001010_0;
      patterns[5560] = 25'b00010101_10110110_11001011_0;
      patterns[5561] = 25'b00010101_10110111_11001100_0;
      patterns[5562] = 25'b00010101_10111000_11001101_0;
      patterns[5563] = 25'b00010101_10111001_11001110_0;
      patterns[5564] = 25'b00010101_10111010_11001111_0;
      patterns[5565] = 25'b00010101_10111011_11010000_0;
      patterns[5566] = 25'b00010101_10111100_11010001_0;
      patterns[5567] = 25'b00010101_10111101_11010010_0;
      patterns[5568] = 25'b00010101_10111110_11010011_0;
      patterns[5569] = 25'b00010101_10111111_11010100_0;
      patterns[5570] = 25'b00010101_11000000_11010101_0;
      patterns[5571] = 25'b00010101_11000001_11010110_0;
      patterns[5572] = 25'b00010101_11000010_11010111_0;
      patterns[5573] = 25'b00010101_11000011_11011000_0;
      patterns[5574] = 25'b00010101_11000100_11011001_0;
      patterns[5575] = 25'b00010101_11000101_11011010_0;
      patterns[5576] = 25'b00010101_11000110_11011011_0;
      patterns[5577] = 25'b00010101_11000111_11011100_0;
      patterns[5578] = 25'b00010101_11001000_11011101_0;
      patterns[5579] = 25'b00010101_11001001_11011110_0;
      patterns[5580] = 25'b00010101_11001010_11011111_0;
      patterns[5581] = 25'b00010101_11001011_11100000_0;
      patterns[5582] = 25'b00010101_11001100_11100001_0;
      patterns[5583] = 25'b00010101_11001101_11100010_0;
      patterns[5584] = 25'b00010101_11001110_11100011_0;
      patterns[5585] = 25'b00010101_11001111_11100100_0;
      patterns[5586] = 25'b00010101_11010000_11100101_0;
      patterns[5587] = 25'b00010101_11010001_11100110_0;
      patterns[5588] = 25'b00010101_11010010_11100111_0;
      patterns[5589] = 25'b00010101_11010011_11101000_0;
      patterns[5590] = 25'b00010101_11010100_11101001_0;
      patterns[5591] = 25'b00010101_11010101_11101010_0;
      patterns[5592] = 25'b00010101_11010110_11101011_0;
      patterns[5593] = 25'b00010101_11010111_11101100_0;
      patterns[5594] = 25'b00010101_11011000_11101101_0;
      patterns[5595] = 25'b00010101_11011001_11101110_0;
      patterns[5596] = 25'b00010101_11011010_11101111_0;
      patterns[5597] = 25'b00010101_11011011_11110000_0;
      patterns[5598] = 25'b00010101_11011100_11110001_0;
      patterns[5599] = 25'b00010101_11011101_11110010_0;
      patterns[5600] = 25'b00010101_11011110_11110011_0;
      patterns[5601] = 25'b00010101_11011111_11110100_0;
      patterns[5602] = 25'b00010101_11100000_11110101_0;
      patterns[5603] = 25'b00010101_11100001_11110110_0;
      patterns[5604] = 25'b00010101_11100010_11110111_0;
      patterns[5605] = 25'b00010101_11100011_11111000_0;
      patterns[5606] = 25'b00010101_11100100_11111001_0;
      patterns[5607] = 25'b00010101_11100101_11111010_0;
      patterns[5608] = 25'b00010101_11100110_11111011_0;
      patterns[5609] = 25'b00010101_11100111_11111100_0;
      patterns[5610] = 25'b00010101_11101000_11111101_0;
      patterns[5611] = 25'b00010101_11101001_11111110_0;
      patterns[5612] = 25'b00010101_11101010_11111111_0;
      patterns[5613] = 25'b00010101_11101011_00000000_1;
      patterns[5614] = 25'b00010101_11101100_00000001_1;
      patterns[5615] = 25'b00010101_11101101_00000010_1;
      patterns[5616] = 25'b00010101_11101110_00000011_1;
      patterns[5617] = 25'b00010101_11101111_00000100_1;
      patterns[5618] = 25'b00010101_11110000_00000101_1;
      patterns[5619] = 25'b00010101_11110001_00000110_1;
      patterns[5620] = 25'b00010101_11110010_00000111_1;
      patterns[5621] = 25'b00010101_11110011_00001000_1;
      patterns[5622] = 25'b00010101_11110100_00001001_1;
      patterns[5623] = 25'b00010101_11110101_00001010_1;
      patterns[5624] = 25'b00010101_11110110_00001011_1;
      patterns[5625] = 25'b00010101_11110111_00001100_1;
      patterns[5626] = 25'b00010101_11111000_00001101_1;
      patterns[5627] = 25'b00010101_11111001_00001110_1;
      patterns[5628] = 25'b00010101_11111010_00001111_1;
      patterns[5629] = 25'b00010101_11111011_00010000_1;
      patterns[5630] = 25'b00010101_11111100_00010001_1;
      patterns[5631] = 25'b00010101_11111101_00010010_1;
      patterns[5632] = 25'b00010101_11111110_00010011_1;
      patterns[5633] = 25'b00010101_11111111_00010100_1;
      patterns[5634] = 25'b00010110_00000000_00010110_0;
      patterns[5635] = 25'b00010110_00000001_00010111_0;
      patterns[5636] = 25'b00010110_00000010_00011000_0;
      patterns[5637] = 25'b00010110_00000011_00011001_0;
      patterns[5638] = 25'b00010110_00000100_00011010_0;
      patterns[5639] = 25'b00010110_00000101_00011011_0;
      patterns[5640] = 25'b00010110_00000110_00011100_0;
      patterns[5641] = 25'b00010110_00000111_00011101_0;
      patterns[5642] = 25'b00010110_00001000_00011110_0;
      patterns[5643] = 25'b00010110_00001001_00011111_0;
      patterns[5644] = 25'b00010110_00001010_00100000_0;
      patterns[5645] = 25'b00010110_00001011_00100001_0;
      patterns[5646] = 25'b00010110_00001100_00100010_0;
      patterns[5647] = 25'b00010110_00001101_00100011_0;
      patterns[5648] = 25'b00010110_00001110_00100100_0;
      patterns[5649] = 25'b00010110_00001111_00100101_0;
      patterns[5650] = 25'b00010110_00010000_00100110_0;
      patterns[5651] = 25'b00010110_00010001_00100111_0;
      patterns[5652] = 25'b00010110_00010010_00101000_0;
      patterns[5653] = 25'b00010110_00010011_00101001_0;
      patterns[5654] = 25'b00010110_00010100_00101010_0;
      patterns[5655] = 25'b00010110_00010101_00101011_0;
      patterns[5656] = 25'b00010110_00010110_00101100_0;
      patterns[5657] = 25'b00010110_00010111_00101101_0;
      patterns[5658] = 25'b00010110_00011000_00101110_0;
      patterns[5659] = 25'b00010110_00011001_00101111_0;
      patterns[5660] = 25'b00010110_00011010_00110000_0;
      patterns[5661] = 25'b00010110_00011011_00110001_0;
      patterns[5662] = 25'b00010110_00011100_00110010_0;
      patterns[5663] = 25'b00010110_00011101_00110011_0;
      patterns[5664] = 25'b00010110_00011110_00110100_0;
      patterns[5665] = 25'b00010110_00011111_00110101_0;
      patterns[5666] = 25'b00010110_00100000_00110110_0;
      patterns[5667] = 25'b00010110_00100001_00110111_0;
      patterns[5668] = 25'b00010110_00100010_00111000_0;
      patterns[5669] = 25'b00010110_00100011_00111001_0;
      patterns[5670] = 25'b00010110_00100100_00111010_0;
      patterns[5671] = 25'b00010110_00100101_00111011_0;
      patterns[5672] = 25'b00010110_00100110_00111100_0;
      patterns[5673] = 25'b00010110_00100111_00111101_0;
      patterns[5674] = 25'b00010110_00101000_00111110_0;
      patterns[5675] = 25'b00010110_00101001_00111111_0;
      patterns[5676] = 25'b00010110_00101010_01000000_0;
      patterns[5677] = 25'b00010110_00101011_01000001_0;
      patterns[5678] = 25'b00010110_00101100_01000010_0;
      patterns[5679] = 25'b00010110_00101101_01000011_0;
      patterns[5680] = 25'b00010110_00101110_01000100_0;
      patterns[5681] = 25'b00010110_00101111_01000101_0;
      patterns[5682] = 25'b00010110_00110000_01000110_0;
      patterns[5683] = 25'b00010110_00110001_01000111_0;
      patterns[5684] = 25'b00010110_00110010_01001000_0;
      patterns[5685] = 25'b00010110_00110011_01001001_0;
      patterns[5686] = 25'b00010110_00110100_01001010_0;
      patterns[5687] = 25'b00010110_00110101_01001011_0;
      patterns[5688] = 25'b00010110_00110110_01001100_0;
      patterns[5689] = 25'b00010110_00110111_01001101_0;
      patterns[5690] = 25'b00010110_00111000_01001110_0;
      patterns[5691] = 25'b00010110_00111001_01001111_0;
      patterns[5692] = 25'b00010110_00111010_01010000_0;
      patterns[5693] = 25'b00010110_00111011_01010001_0;
      patterns[5694] = 25'b00010110_00111100_01010010_0;
      patterns[5695] = 25'b00010110_00111101_01010011_0;
      patterns[5696] = 25'b00010110_00111110_01010100_0;
      patterns[5697] = 25'b00010110_00111111_01010101_0;
      patterns[5698] = 25'b00010110_01000000_01010110_0;
      patterns[5699] = 25'b00010110_01000001_01010111_0;
      patterns[5700] = 25'b00010110_01000010_01011000_0;
      patterns[5701] = 25'b00010110_01000011_01011001_0;
      patterns[5702] = 25'b00010110_01000100_01011010_0;
      patterns[5703] = 25'b00010110_01000101_01011011_0;
      patterns[5704] = 25'b00010110_01000110_01011100_0;
      patterns[5705] = 25'b00010110_01000111_01011101_0;
      patterns[5706] = 25'b00010110_01001000_01011110_0;
      patterns[5707] = 25'b00010110_01001001_01011111_0;
      patterns[5708] = 25'b00010110_01001010_01100000_0;
      patterns[5709] = 25'b00010110_01001011_01100001_0;
      patterns[5710] = 25'b00010110_01001100_01100010_0;
      patterns[5711] = 25'b00010110_01001101_01100011_0;
      patterns[5712] = 25'b00010110_01001110_01100100_0;
      patterns[5713] = 25'b00010110_01001111_01100101_0;
      patterns[5714] = 25'b00010110_01010000_01100110_0;
      patterns[5715] = 25'b00010110_01010001_01100111_0;
      patterns[5716] = 25'b00010110_01010010_01101000_0;
      patterns[5717] = 25'b00010110_01010011_01101001_0;
      patterns[5718] = 25'b00010110_01010100_01101010_0;
      patterns[5719] = 25'b00010110_01010101_01101011_0;
      patterns[5720] = 25'b00010110_01010110_01101100_0;
      patterns[5721] = 25'b00010110_01010111_01101101_0;
      patterns[5722] = 25'b00010110_01011000_01101110_0;
      patterns[5723] = 25'b00010110_01011001_01101111_0;
      patterns[5724] = 25'b00010110_01011010_01110000_0;
      patterns[5725] = 25'b00010110_01011011_01110001_0;
      patterns[5726] = 25'b00010110_01011100_01110010_0;
      patterns[5727] = 25'b00010110_01011101_01110011_0;
      patterns[5728] = 25'b00010110_01011110_01110100_0;
      patterns[5729] = 25'b00010110_01011111_01110101_0;
      patterns[5730] = 25'b00010110_01100000_01110110_0;
      patterns[5731] = 25'b00010110_01100001_01110111_0;
      patterns[5732] = 25'b00010110_01100010_01111000_0;
      patterns[5733] = 25'b00010110_01100011_01111001_0;
      patterns[5734] = 25'b00010110_01100100_01111010_0;
      patterns[5735] = 25'b00010110_01100101_01111011_0;
      patterns[5736] = 25'b00010110_01100110_01111100_0;
      patterns[5737] = 25'b00010110_01100111_01111101_0;
      patterns[5738] = 25'b00010110_01101000_01111110_0;
      patterns[5739] = 25'b00010110_01101001_01111111_0;
      patterns[5740] = 25'b00010110_01101010_10000000_0;
      patterns[5741] = 25'b00010110_01101011_10000001_0;
      patterns[5742] = 25'b00010110_01101100_10000010_0;
      patterns[5743] = 25'b00010110_01101101_10000011_0;
      patterns[5744] = 25'b00010110_01101110_10000100_0;
      patterns[5745] = 25'b00010110_01101111_10000101_0;
      patterns[5746] = 25'b00010110_01110000_10000110_0;
      patterns[5747] = 25'b00010110_01110001_10000111_0;
      patterns[5748] = 25'b00010110_01110010_10001000_0;
      patterns[5749] = 25'b00010110_01110011_10001001_0;
      patterns[5750] = 25'b00010110_01110100_10001010_0;
      patterns[5751] = 25'b00010110_01110101_10001011_0;
      patterns[5752] = 25'b00010110_01110110_10001100_0;
      patterns[5753] = 25'b00010110_01110111_10001101_0;
      patterns[5754] = 25'b00010110_01111000_10001110_0;
      patterns[5755] = 25'b00010110_01111001_10001111_0;
      patterns[5756] = 25'b00010110_01111010_10010000_0;
      patterns[5757] = 25'b00010110_01111011_10010001_0;
      patterns[5758] = 25'b00010110_01111100_10010010_0;
      patterns[5759] = 25'b00010110_01111101_10010011_0;
      patterns[5760] = 25'b00010110_01111110_10010100_0;
      patterns[5761] = 25'b00010110_01111111_10010101_0;
      patterns[5762] = 25'b00010110_10000000_10010110_0;
      patterns[5763] = 25'b00010110_10000001_10010111_0;
      patterns[5764] = 25'b00010110_10000010_10011000_0;
      patterns[5765] = 25'b00010110_10000011_10011001_0;
      patterns[5766] = 25'b00010110_10000100_10011010_0;
      patterns[5767] = 25'b00010110_10000101_10011011_0;
      patterns[5768] = 25'b00010110_10000110_10011100_0;
      patterns[5769] = 25'b00010110_10000111_10011101_0;
      patterns[5770] = 25'b00010110_10001000_10011110_0;
      patterns[5771] = 25'b00010110_10001001_10011111_0;
      patterns[5772] = 25'b00010110_10001010_10100000_0;
      patterns[5773] = 25'b00010110_10001011_10100001_0;
      patterns[5774] = 25'b00010110_10001100_10100010_0;
      patterns[5775] = 25'b00010110_10001101_10100011_0;
      patterns[5776] = 25'b00010110_10001110_10100100_0;
      patterns[5777] = 25'b00010110_10001111_10100101_0;
      patterns[5778] = 25'b00010110_10010000_10100110_0;
      patterns[5779] = 25'b00010110_10010001_10100111_0;
      patterns[5780] = 25'b00010110_10010010_10101000_0;
      patterns[5781] = 25'b00010110_10010011_10101001_0;
      patterns[5782] = 25'b00010110_10010100_10101010_0;
      patterns[5783] = 25'b00010110_10010101_10101011_0;
      patterns[5784] = 25'b00010110_10010110_10101100_0;
      patterns[5785] = 25'b00010110_10010111_10101101_0;
      patterns[5786] = 25'b00010110_10011000_10101110_0;
      patterns[5787] = 25'b00010110_10011001_10101111_0;
      patterns[5788] = 25'b00010110_10011010_10110000_0;
      patterns[5789] = 25'b00010110_10011011_10110001_0;
      patterns[5790] = 25'b00010110_10011100_10110010_0;
      patterns[5791] = 25'b00010110_10011101_10110011_0;
      patterns[5792] = 25'b00010110_10011110_10110100_0;
      patterns[5793] = 25'b00010110_10011111_10110101_0;
      patterns[5794] = 25'b00010110_10100000_10110110_0;
      patterns[5795] = 25'b00010110_10100001_10110111_0;
      patterns[5796] = 25'b00010110_10100010_10111000_0;
      patterns[5797] = 25'b00010110_10100011_10111001_0;
      patterns[5798] = 25'b00010110_10100100_10111010_0;
      patterns[5799] = 25'b00010110_10100101_10111011_0;
      patterns[5800] = 25'b00010110_10100110_10111100_0;
      patterns[5801] = 25'b00010110_10100111_10111101_0;
      patterns[5802] = 25'b00010110_10101000_10111110_0;
      patterns[5803] = 25'b00010110_10101001_10111111_0;
      patterns[5804] = 25'b00010110_10101010_11000000_0;
      patterns[5805] = 25'b00010110_10101011_11000001_0;
      patterns[5806] = 25'b00010110_10101100_11000010_0;
      patterns[5807] = 25'b00010110_10101101_11000011_0;
      patterns[5808] = 25'b00010110_10101110_11000100_0;
      patterns[5809] = 25'b00010110_10101111_11000101_0;
      patterns[5810] = 25'b00010110_10110000_11000110_0;
      patterns[5811] = 25'b00010110_10110001_11000111_0;
      patterns[5812] = 25'b00010110_10110010_11001000_0;
      patterns[5813] = 25'b00010110_10110011_11001001_0;
      patterns[5814] = 25'b00010110_10110100_11001010_0;
      patterns[5815] = 25'b00010110_10110101_11001011_0;
      patterns[5816] = 25'b00010110_10110110_11001100_0;
      patterns[5817] = 25'b00010110_10110111_11001101_0;
      patterns[5818] = 25'b00010110_10111000_11001110_0;
      patterns[5819] = 25'b00010110_10111001_11001111_0;
      patterns[5820] = 25'b00010110_10111010_11010000_0;
      patterns[5821] = 25'b00010110_10111011_11010001_0;
      patterns[5822] = 25'b00010110_10111100_11010010_0;
      patterns[5823] = 25'b00010110_10111101_11010011_0;
      patterns[5824] = 25'b00010110_10111110_11010100_0;
      patterns[5825] = 25'b00010110_10111111_11010101_0;
      patterns[5826] = 25'b00010110_11000000_11010110_0;
      patterns[5827] = 25'b00010110_11000001_11010111_0;
      patterns[5828] = 25'b00010110_11000010_11011000_0;
      patterns[5829] = 25'b00010110_11000011_11011001_0;
      patterns[5830] = 25'b00010110_11000100_11011010_0;
      patterns[5831] = 25'b00010110_11000101_11011011_0;
      patterns[5832] = 25'b00010110_11000110_11011100_0;
      patterns[5833] = 25'b00010110_11000111_11011101_0;
      patterns[5834] = 25'b00010110_11001000_11011110_0;
      patterns[5835] = 25'b00010110_11001001_11011111_0;
      patterns[5836] = 25'b00010110_11001010_11100000_0;
      patterns[5837] = 25'b00010110_11001011_11100001_0;
      patterns[5838] = 25'b00010110_11001100_11100010_0;
      patterns[5839] = 25'b00010110_11001101_11100011_0;
      patterns[5840] = 25'b00010110_11001110_11100100_0;
      patterns[5841] = 25'b00010110_11001111_11100101_0;
      patterns[5842] = 25'b00010110_11010000_11100110_0;
      patterns[5843] = 25'b00010110_11010001_11100111_0;
      patterns[5844] = 25'b00010110_11010010_11101000_0;
      patterns[5845] = 25'b00010110_11010011_11101001_0;
      patterns[5846] = 25'b00010110_11010100_11101010_0;
      patterns[5847] = 25'b00010110_11010101_11101011_0;
      patterns[5848] = 25'b00010110_11010110_11101100_0;
      patterns[5849] = 25'b00010110_11010111_11101101_0;
      patterns[5850] = 25'b00010110_11011000_11101110_0;
      patterns[5851] = 25'b00010110_11011001_11101111_0;
      patterns[5852] = 25'b00010110_11011010_11110000_0;
      patterns[5853] = 25'b00010110_11011011_11110001_0;
      patterns[5854] = 25'b00010110_11011100_11110010_0;
      patterns[5855] = 25'b00010110_11011101_11110011_0;
      patterns[5856] = 25'b00010110_11011110_11110100_0;
      patterns[5857] = 25'b00010110_11011111_11110101_0;
      patterns[5858] = 25'b00010110_11100000_11110110_0;
      patterns[5859] = 25'b00010110_11100001_11110111_0;
      patterns[5860] = 25'b00010110_11100010_11111000_0;
      patterns[5861] = 25'b00010110_11100011_11111001_0;
      patterns[5862] = 25'b00010110_11100100_11111010_0;
      patterns[5863] = 25'b00010110_11100101_11111011_0;
      patterns[5864] = 25'b00010110_11100110_11111100_0;
      patterns[5865] = 25'b00010110_11100111_11111101_0;
      patterns[5866] = 25'b00010110_11101000_11111110_0;
      patterns[5867] = 25'b00010110_11101001_11111111_0;
      patterns[5868] = 25'b00010110_11101010_00000000_1;
      patterns[5869] = 25'b00010110_11101011_00000001_1;
      patterns[5870] = 25'b00010110_11101100_00000010_1;
      patterns[5871] = 25'b00010110_11101101_00000011_1;
      patterns[5872] = 25'b00010110_11101110_00000100_1;
      patterns[5873] = 25'b00010110_11101111_00000101_1;
      patterns[5874] = 25'b00010110_11110000_00000110_1;
      patterns[5875] = 25'b00010110_11110001_00000111_1;
      patterns[5876] = 25'b00010110_11110010_00001000_1;
      patterns[5877] = 25'b00010110_11110011_00001001_1;
      patterns[5878] = 25'b00010110_11110100_00001010_1;
      patterns[5879] = 25'b00010110_11110101_00001011_1;
      patterns[5880] = 25'b00010110_11110110_00001100_1;
      patterns[5881] = 25'b00010110_11110111_00001101_1;
      patterns[5882] = 25'b00010110_11111000_00001110_1;
      patterns[5883] = 25'b00010110_11111001_00001111_1;
      patterns[5884] = 25'b00010110_11111010_00010000_1;
      patterns[5885] = 25'b00010110_11111011_00010001_1;
      patterns[5886] = 25'b00010110_11111100_00010010_1;
      patterns[5887] = 25'b00010110_11111101_00010011_1;
      patterns[5888] = 25'b00010110_11111110_00010100_1;
      patterns[5889] = 25'b00010110_11111111_00010101_1;
      patterns[5890] = 25'b00010111_00000000_00010111_0;
      patterns[5891] = 25'b00010111_00000001_00011000_0;
      patterns[5892] = 25'b00010111_00000010_00011001_0;
      patterns[5893] = 25'b00010111_00000011_00011010_0;
      patterns[5894] = 25'b00010111_00000100_00011011_0;
      patterns[5895] = 25'b00010111_00000101_00011100_0;
      patterns[5896] = 25'b00010111_00000110_00011101_0;
      patterns[5897] = 25'b00010111_00000111_00011110_0;
      patterns[5898] = 25'b00010111_00001000_00011111_0;
      patterns[5899] = 25'b00010111_00001001_00100000_0;
      patterns[5900] = 25'b00010111_00001010_00100001_0;
      patterns[5901] = 25'b00010111_00001011_00100010_0;
      patterns[5902] = 25'b00010111_00001100_00100011_0;
      patterns[5903] = 25'b00010111_00001101_00100100_0;
      patterns[5904] = 25'b00010111_00001110_00100101_0;
      patterns[5905] = 25'b00010111_00001111_00100110_0;
      patterns[5906] = 25'b00010111_00010000_00100111_0;
      patterns[5907] = 25'b00010111_00010001_00101000_0;
      patterns[5908] = 25'b00010111_00010010_00101001_0;
      patterns[5909] = 25'b00010111_00010011_00101010_0;
      patterns[5910] = 25'b00010111_00010100_00101011_0;
      patterns[5911] = 25'b00010111_00010101_00101100_0;
      patterns[5912] = 25'b00010111_00010110_00101101_0;
      patterns[5913] = 25'b00010111_00010111_00101110_0;
      patterns[5914] = 25'b00010111_00011000_00101111_0;
      patterns[5915] = 25'b00010111_00011001_00110000_0;
      patterns[5916] = 25'b00010111_00011010_00110001_0;
      patterns[5917] = 25'b00010111_00011011_00110010_0;
      patterns[5918] = 25'b00010111_00011100_00110011_0;
      patterns[5919] = 25'b00010111_00011101_00110100_0;
      patterns[5920] = 25'b00010111_00011110_00110101_0;
      patterns[5921] = 25'b00010111_00011111_00110110_0;
      patterns[5922] = 25'b00010111_00100000_00110111_0;
      patterns[5923] = 25'b00010111_00100001_00111000_0;
      patterns[5924] = 25'b00010111_00100010_00111001_0;
      patterns[5925] = 25'b00010111_00100011_00111010_0;
      patterns[5926] = 25'b00010111_00100100_00111011_0;
      patterns[5927] = 25'b00010111_00100101_00111100_0;
      patterns[5928] = 25'b00010111_00100110_00111101_0;
      patterns[5929] = 25'b00010111_00100111_00111110_0;
      patterns[5930] = 25'b00010111_00101000_00111111_0;
      patterns[5931] = 25'b00010111_00101001_01000000_0;
      patterns[5932] = 25'b00010111_00101010_01000001_0;
      patterns[5933] = 25'b00010111_00101011_01000010_0;
      patterns[5934] = 25'b00010111_00101100_01000011_0;
      patterns[5935] = 25'b00010111_00101101_01000100_0;
      patterns[5936] = 25'b00010111_00101110_01000101_0;
      patterns[5937] = 25'b00010111_00101111_01000110_0;
      patterns[5938] = 25'b00010111_00110000_01000111_0;
      patterns[5939] = 25'b00010111_00110001_01001000_0;
      patterns[5940] = 25'b00010111_00110010_01001001_0;
      patterns[5941] = 25'b00010111_00110011_01001010_0;
      patterns[5942] = 25'b00010111_00110100_01001011_0;
      patterns[5943] = 25'b00010111_00110101_01001100_0;
      patterns[5944] = 25'b00010111_00110110_01001101_0;
      patterns[5945] = 25'b00010111_00110111_01001110_0;
      patterns[5946] = 25'b00010111_00111000_01001111_0;
      patterns[5947] = 25'b00010111_00111001_01010000_0;
      patterns[5948] = 25'b00010111_00111010_01010001_0;
      patterns[5949] = 25'b00010111_00111011_01010010_0;
      patterns[5950] = 25'b00010111_00111100_01010011_0;
      patterns[5951] = 25'b00010111_00111101_01010100_0;
      patterns[5952] = 25'b00010111_00111110_01010101_0;
      patterns[5953] = 25'b00010111_00111111_01010110_0;
      patterns[5954] = 25'b00010111_01000000_01010111_0;
      patterns[5955] = 25'b00010111_01000001_01011000_0;
      patterns[5956] = 25'b00010111_01000010_01011001_0;
      patterns[5957] = 25'b00010111_01000011_01011010_0;
      patterns[5958] = 25'b00010111_01000100_01011011_0;
      patterns[5959] = 25'b00010111_01000101_01011100_0;
      patterns[5960] = 25'b00010111_01000110_01011101_0;
      patterns[5961] = 25'b00010111_01000111_01011110_0;
      patterns[5962] = 25'b00010111_01001000_01011111_0;
      patterns[5963] = 25'b00010111_01001001_01100000_0;
      patterns[5964] = 25'b00010111_01001010_01100001_0;
      patterns[5965] = 25'b00010111_01001011_01100010_0;
      patterns[5966] = 25'b00010111_01001100_01100011_0;
      patterns[5967] = 25'b00010111_01001101_01100100_0;
      patterns[5968] = 25'b00010111_01001110_01100101_0;
      patterns[5969] = 25'b00010111_01001111_01100110_0;
      patterns[5970] = 25'b00010111_01010000_01100111_0;
      patterns[5971] = 25'b00010111_01010001_01101000_0;
      patterns[5972] = 25'b00010111_01010010_01101001_0;
      patterns[5973] = 25'b00010111_01010011_01101010_0;
      patterns[5974] = 25'b00010111_01010100_01101011_0;
      patterns[5975] = 25'b00010111_01010101_01101100_0;
      patterns[5976] = 25'b00010111_01010110_01101101_0;
      patterns[5977] = 25'b00010111_01010111_01101110_0;
      patterns[5978] = 25'b00010111_01011000_01101111_0;
      patterns[5979] = 25'b00010111_01011001_01110000_0;
      patterns[5980] = 25'b00010111_01011010_01110001_0;
      patterns[5981] = 25'b00010111_01011011_01110010_0;
      patterns[5982] = 25'b00010111_01011100_01110011_0;
      patterns[5983] = 25'b00010111_01011101_01110100_0;
      patterns[5984] = 25'b00010111_01011110_01110101_0;
      patterns[5985] = 25'b00010111_01011111_01110110_0;
      patterns[5986] = 25'b00010111_01100000_01110111_0;
      patterns[5987] = 25'b00010111_01100001_01111000_0;
      patterns[5988] = 25'b00010111_01100010_01111001_0;
      patterns[5989] = 25'b00010111_01100011_01111010_0;
      patterns[5990] = 25'b00010111_01100100_01111011_0;
      patterns[5991] = 25'b00010111_01100101_01111100_0;
      patterns[5992] = 25'b00010111_01100110_01111101_0;
      patterns[5993] = 25'b00010111_01100111_01111110_0;
      patterns[5994] = 25'b00010111_01101000_01111111_0;
      patterns[5995] = 25'b00010111_01101001_10000000_0;
      patterns[5996] = 25'b00010111_01101010_10000001_0;
      patterns[5997] = 25'b00010111_01101011_10000010_0;
      patterns[5998] = 25'b00010111_01101100_10000011_0;
      patterns[5999] = 25'b00010111_01101101_10000100_0;
      patterns[6000] = 25'b00010111_01101110_10000101_0;
      patterns[6001] = 25'b00010111_01101111_10000110_0;
      patterns[6002] = 25'b00010111_01110000_10000111_0;
      patterns[6003] = 25'b00010111_01110001_10001000_0;
      patterns[6004] = 25'b00010111_01110010_10001001_0;
      patterns[6005] = 25'b00010111_01110011_10001010_0;
      patterns[6006] = 25'b00010111_01110100_10001011_0;
      patterns[6007] = 25'b00010111_01110101_10001100_0;
      patterns[6008] = 25'b00010111_01110110_10001101_0;
      patterns[6009] = 25'b00010111_01110111_10001110_0;
      patterns[6010] = 25'b00010111_01111000_10001111_0;
      patterns[6011] = 25'b00010111_01111001_10010000_0;
      patterns[6012] = 25'b00010111_01111010_10010001_0;
      patterns[6013] = 25'b00010111_01111011_10010010_0;
      patterns[6014] = 25'b00010111_01111100_10010011_0;
      patterns[6015] = 25'b00010111_01111101_10010100_0;
      patterns[6016] = 25'b00010111_01111110_10010101_0;
      patterns[6017] = 25'b00010111_01111111_10010110_0;
      patterns[6018] = 25'b00010111_10000000_10010111_0;
      patterns[6019] = 25'b00010111_10000001_10011000_0;
      patterns[6020] = 25'b00010111_10000010_10011001_0;
      patterns[6021] = 25'b00010111_10000011_10011010_0;
      patterns[6022] = 25'b00010111_10000100_10011011_0;
      patterns[6023] = 25'b00010111_10000101_10011100_0;
      patterns[6024] = 25'b00010111_10000110_10011101_0;
      patterns[6025] = 25'b00010111_10000111_10011110_0;
      patterns[6026] = 25'b00010111_10001000_10011111_0;
      patterns[6027] = 25'b00010111_10001001_10100000_0;
      patterns[6028] = 25'b00010111_10001010_10100001_0;
      patterns[6029] = 25'b00010111_10001011_10100010_0;
      patterns[6030] = 25'b00010111_10001100_10100011_0;
      patterns[6031] = 25'b00010111_10001101_10100100_0;
      patterns[6032] = 25'b00010111_10001110_10100101_0;
      patterns[6033] = 25'b00010111_10001111_10100110_0;
      patterns[6034] = 25'b00010111_10010000_10100111_0;
      patterns[6035] = 25'b00010111_10010001_10101000_0;
      patterns[6036] = 25'b00010111_10010010_10101001_0;
      patterns[6037] = 25'b00010111_10010011_10101010_0;
      patterns[6038] = 25'b00010111_10010100_10101011_0;
      patterns[6039] = 25'b00010111_10010101_10101100_0;
      patterns[6040] = 25'b00010111_10010110_10101101_0;
      patterns[6041] = 25'b00010111_10010111_10101110_0;
      patterns[6042] = 25'b00010111_10011000_10101111_0;
      patterns[6043] = 25'b00010111_10011001_10110000_0;
      patterns[6044] = 25'b00010111_10011010_10110001_0;
      patterns[6045] = 25'b00010111_10011011_10110010_0;
      patterns[6046] = 25'b00010111_10011100_10110011_0;
      patterns[6047] = 25'b00010111_10011101_10110100_0;
      patterns[6048] = 25'b00010111_10011110_10110101_0;
      patterns[6049] = 25'b00010111_10011111_10110110_0;
      patterns[6050] = 25'b00010111_10100000_10110111_0;
      patterns[6051] = 25'b00010111_10100001_10111000_0;
      patterns[6052] = 25'b00010111_10100010_10111001_0;
      patterns[6053] = 25'b00010111_10100011_10111010_0;
      patterns[6054] = 25'b00010111_10100100_10111011_0;
      patterns[6055] = 25'b00010111_10100101_10111100_0;
      patterns[6056] = 25'b00010111_10100110_10111101_0;
      patterns[6057] = 25'b00010111_10100111_10111110_0;
      patterns[6058] = 25'b00010111_10101000_10111111_0;
      patterns[6059] = 25'b00010111_10101001_11000000_0;
      patterns[6060] = 25'b00010111_10101010_11000001_0;
      patterns[6061] = 25'b00010111_10101011_11000010_0;
      patterns[6062] = 25'b00010111_10101100_11000011_0;
      patterns[6063] = 25'b00010111_10101101_11000100_0;
      patterns[6064] = 25'b00010111_10101110_11000101_0;
      patterns[6065] = 25'b00010111_10101111_11000110_0;
      patterns[6066] = 25'b00010111_10110000_11000111_0;
      patterns[6067] = 25'b00010111_10110001_11001000_0;
      patterns[6068] = 25'b00010111_10110010_11001001_0;
      patterns[6069] = 25'b00010111_10110011_11001010_0;
      patterns[6070] = 25'b00010111_10110100_11001011_0;
      patterns[6071] = 25'b00010111_10110101_11001100_0;
      patterns[6072] = 25'b00010111_10110110_11001101_0;
      patterns[6073] = 25'b00010111_10110111_11001110_0;
      patterns[6074] = 25'b00010111_10111000_11001111_0;
      patterns[6075] = 25'b00010111_10111001_11010000_0;
      patterns[6076] = 25'b00010111_10111010_11010001_0;
      patterns[6077] = 25'b00010111_10111011_11010010_0;
      patterns[6078] = 25'b00010111_10111100_11010011_0;
      patterns[6079] = 25'b00010111_10111101_11010100_0;
      patterns[6080] = 25'b00010111_10111110_11010101_0;
      patterns[6081] = 25'b00010111_10111111_11010110_0;
      patterns[6082] = 25'b00010111_11000000_11010111_0;
      patterns[6083] = 25'b00010111_11000001_11011000_0;
      patterns[6084] = 25'b00010111_11000010_11011001_0;
      patterns[6085] = 25'b00010111_11000011_11011010_0;
      patterns[6086] = 25'b00010111_11000100_11011011_0;
      patterns[6087] = 25'b00010111_11000101_11011100_0;
      patterns[6088] = 25'b00010111_11000110_11011101_0;
      patterns[6089] = 25'b00010111_11000111_11011110_0;
      patterns[6090] = 25'b00010111_11001000_11011111_0;
      patterns[6091] = 25'b00010111_11001001_11100000_0;
      patterns[6092] = 25'b00010111_11001010_11100001_0;
      patterns[6093] = 25'b00010111_11001011_11100010_0;
      patterns[6094] = 25'b00010111_11001100_11100011_0;
      patterns[6095] = 25'b00010111_11001101_11100100_0;
      patterns[6096] = 25'b00010111_11001110_11100101_0;
      patterns[6097] = 25'b00010111_11001111_11100110_0;
      patterns[6098] = 25'b00010111_11010000_11100111_0;
      patterns[6099] = 25'b00010111_11010001_11101000_0;
      patterns[6100] = 25'b00010111_11010010_11101001_0;
      patterns[6101] = 25'b00010111_11010011_11101010_0;
      patterns[6102] = 25'b00010111_11010100_11101011_0;
      patterns[6103] = 25'b00010111_11010101_11101100_0;
      patterns[6104] = 25'b00010111_11010110_11101101_0;
      patterns[6105] = 25'b00010111_11010111_11101110_0;
      patterns[6106] = 25'b00010111_11011000_11101111_0;
      patterns[6107] = 25'b00010111_11011001_11110000_0;
      patterns[6108] = 25'b00010111_11011010_11110001_0;
      patterns[6109] = 25'b00010111_11011011_11110010_0;
      patterns[6110] = 25'b00010111_11011100_11110011_0;
      patterns[6111] = 25'b00010111_11011101_11110100_0;
      patterns[6112] = 25'b00010111_11011110_11110101_0;
      patterns[6113] = 25'b00010111_11011111_11110110_0;
      patterns[6114] = 25'b00010111_11100000_11110111_0;
      patterns[6115] = 25'b00010111_11100001_11111000_0;
      patterns[6116] = 25'b00010111_11100010_11111001_0;
      patterns[6117] = 25'b00010111_11100011_11111010_0;
      patterns[6118] = 25'b00010111_11100100_11111011_0;
      patterns[6119] = 25'b00010111_11100101_11111100_0;
      patterns[6120] = 25'b00010111_11100110_11111101_0;
      patterns[6121] = 25'b00010111_11100111_11111110_0;
      patterns[6122] = 25'b00010111_11101000_11111111_0;
      patterns[6123] = 25'b00010111_11101001_00000000_1;
      patterns[6124] = 25'b00010111_11101010_00000001_1;
      patterns[6125] = 25'b00010111_11101011_00000010_1;
      patterns[6126] = 25'b00010111_11101100_00000011_1;
      patterns[6127] = 25'b00010111_11101101_00000100_1;
      patterns[6128] = 25'b00010111_11101110_00000101_1;
      patterns[6129] = 25'b00010111_11101111_00000110_1;
      patterns[6130] = 25'b00010111_11110000_00000111_1;
      patterns[6131] = 25'b00010111_11110001_00001000_1;
      patterns[6132] = 25'b00010111_11110010_00001001_1;
      patterns[6133] = 25'b00010111_11110011_00001010_1;
      patterns[6134] = 25'b00010111_11110100_00001011_1;
      patterns[6135] = 25'b00010111_11110101_00001100_1;
      patterns[6136] = 25'b00010111_11110110_00001101_1;
      patterns[6137] = 25'b00010111_11110111_00001110_1;
      patterns[6138] = 25'b00010111_11111000_00001111_1;
      patterns[6139] = 25'b00010111_11111001_00010000_1;
      patterns[6140] = 25'b00010111_11111010_00010001_1;
      patterns[6141] = 25'b00010111_11111011_00010010_1;
      patterns[6142] = 25'b00010111_11111100_00010011_1;
      patterns[6143] = 25'b00010111_11111101_00010100_1;
      patterns[6144] = 25'b00010111_11111110_00010101_1;
      patterns[6145] = 25'b00010111_11111111_00010110_1;
      patterns[6146] = 25'b00011000_00000000_00011000_0;
      patterns[6147] = 25'b00011000_00000001_00011001_0;
      patterns[6148] = 25'b00011000_00000010_00011010_0;
      patterns[6149] = 25'b00011000_00000011_00011011_0;
      patterns[6150] = 25'b00011000_00000100_00011100_0;
      patterns[6151] = 25'b00011000_00000101_00011101_0;
      patterns[6152] = 25'b00011000_00000110_00011110_0;
      patterns[6153] = 25'b00011000_00000111_00011111_0;
      patterns[6154] = 25'b00011000_00001000_00100000_0;
      patterns[6155] = 25'b00011000_00001001_00100001_0;
      patterns[6156] = 25'b00011000_00001010_00100010_0;
      patterns[6157] = 25'b00011000_00001011_00100011_0;
      patterns[6158] = 25'b00011000_00001100_00100100_0;
      patterns[6159] = 25'b00011000_00001101_00100101_0;
      patterns[6160] = 25'b00011000_00001110_00100110_0;
      patterns[6161] = 25'b00011000_00001111_00100111_0;
      patterns[6162] = 25'b00011000_00010000_00101000_0;
      patterns[6163] = 25'b00011000_00010001_00101001_0;
      patterns[6164] = 25'b00011000_00010010_00101010_0;
      patterns[6165] = 25'b00011000_00010011_00101011_0;
      patterns[6166] = 25'b00011000_00010100_00101100_0;
      patterns[6167] = 25'b00011000_00010101_00101101_0;
      patterns[6168] = 25'b00011000_00010110_00101110_0;
      patterns[6169] = 25'b00011000_00010111_00101111_0;
      patterns[6170] = 25'b00011000_00011000_00110000_0;
      patterns[6171] = 25'b00011000_00011001_00110001_0;
      patterns[6172] = 25'b00011000_00011010_00110010_0;
      patterns[6173] = 25'b00011000_00011011_00110011_0;
      patterns[6174] = 25'b00011000_00011100_00110100_0;
      patterns[6175] = 25'b00011000_00011101_00110101_0;
      patterns[6176] = 25'b00011000_00011110_00110110_0;
      patterns[6177] = 25'b00011000_00011111_00110111_0;
      patterns[6178] = 25'b00011000_00100000_00111000_0;
      patterns[6179] = 25'b00011000_00100001_00111001_0;
      patterns[6180] = 25'b00011000_00100010_00111010_0;
      patterns[6181] = 25'b00011000_00100011_00111011_0;
      patterns[6182] = 25'b00011000_00100100_00111100_0;
      patterns[6183] = 25'b00011000_00100101_00111101_0;
      patterns[6184] = 25'b00011000_00100110_00111110_0;
      patterns[6185] = 25'b00011000_00100111_00111111_0;
      patterns[6186] = 25'b00011000_00101000_01000000_0;
      patterns[6187] = 25'b00011000_00101001_01000001_0;
      patterns[6188] = 25'b00011000_00101010_01000010_0;
      patterns[6189] = 25'b00011000_00101011_01000011_0;
      patterns[6190] = 25'b00011000_00101100_01000100_0;
      patterns[6191] = 25'b00011000_00101101_01000101_0;
      patterns[6192] = 25'b00011000_00101110_01000110_0;
      patterns[6193] = 25'b00011000_00101111_01000111_0;
      patterns[6194] = 25'b00011000_00110000_01001000_0;
      patterns[6195] = 25'b00011000_00110001_01001001_0;
      patterns[6196] = 25'b00011000_00110010_01001010_0;
      patterns[6197] = 25'b00011000_00110011_01001011_0;
      patterns[6198] = 25'b00011000_00110100_01001100_0;
      patterns[6199] = 25'b00011000_00110101_01001101_0;
      patterns[6200] = 25'b00011000_00110110_01001110_0;
      patterns[6201] = 25'b00011000_00110111_01001111_0;
      patterns[6202] = 25'b00011000_00111000_01010000_0;
      patterns[6203] = 25'b00011000_00111001_01010001_0;
      patterns[6204] = 25'b00011000_00111010_01010010_0;
      patterns[6205] = 25'b00011000_00111011_01010011_0;
      patterns[6206] = 25'b00011000_00111100_01010100_0;
      patterns[6207] = 25'b00011000_00111101_01010101_0;
      patterns[6208] = 25'b00011000_00111110_01010110_0;
      patterns[6209] = 25'b00011000_00111111_01010111_0;
      patterns[6210] = 25'b00011000_01000000_01011000_0;
      patterns[6211] = 25'b00011000_01000001_01011001_0;
      patterns[6212] = 25'b00011000_01000010_01011010_0;
      patterns[6213] = 25'b00011000_01000011_01011011_0;
      patterns[6214] = 25'b00011000_01000100_01011100_0;
      patterns[6215] = 25'b00011000_01000101_01011101_0;
      patterns[6216] = 25'b00011000_01000110_01011110_0;
      patterns[6217] = 25'b00011000_01000111_01011111_0;
      patterns[6218] = 25'b00011000_01001000_01100000_0;
      patterns[6219] = 25'b00011000_01001001_01100001_0;
      patterns[6220] = 25'b00011000_01001010_01100010_0;
      patterns[6221] = 25'b00011000_01001011_01100011_0;
      patterns[6222] = 25'b00011000_01001100_01100100_0;
      patterns[6223] = 25'b00011000_01001101_01100101_0;
      patterns[6224] = 25'b00011000_01001110_01100110_0;
      patterns[6225] = 25'b00011000_01001111_01100111_0;
      patterns[6226] = 25'b00011000_01010000_01101000_0;
      patterns[6227] = 25'b00011000_01010001_01101001_0;
      patterns[6228] = 25'b00011000_01010010_01101010_0;
      patterns[6229] = 25'b00011000_01010011_01101011_0;
      patterns[6230] = 25'b00011000_01010100_01101100_0;
      patterns[6231] = 25'b00011000_01010101_01101101_0;
      patterns[6232] = 25'b00011000_01010110_01101110_0;
      patterns[6233] = 25'b00011000_01010111_01101111_0;
      patterns[6234] = 25'b00011000_01011000_01110000_0;
      patterns[6235] = 25'b00011000_01011001_01110001_0;
      patterns[6236] = 25'b00011000_01011010_01110010_0;
      patterns[6237] = 25'b00011000_01011011_01110011_0;
      patterns[6238] = 25'b00011000_01011100_01110100_0;
      patterns[6239] = 25'b00011000_01011101_01110101_0;
      patterns[6240] = 25'b00011000_01011110_01110110_0;
      patterns[6241] = 25'b00011000_01011111_01110111_0;
      patterns[6242] = 25'b00011000_01100000_01111000_0;
      patterns[6243] = 25'b00011000_01100001_01111001_0;
      patterns[6244] = 25'b00011000_01100010_01111010_0;
      patterns[6245] = 25'b00011000_01100011_01111011_0;
      patterns[6246] = 25'b00011000_01100100_01111100_0;
      patterns[6247] = 25'b00011000_01100101_01111101_0;
      patterns[6248] = 25'b00011000_01100110_01111110_0;
      patterns[6249] = 25'b00011000_01100111_01111111_0;
      patterns[6250] = 25'b00011000_01101000_10000000_0;
      patterns[6251] = 25'b00011000_01101001_10000001_0;
      patterns[6252] = 25'b00011000_01101010_10000010_0;
      patterns[6253] = 25'b00011000_01101011_10000011_0;
      patterns[6254] = 25'b00011000_01101100_10000100_0;
      patterns[6255] = 25'b00011000_01101101_10000101_0;
      patterns[6256] = 25'b00011000_01101110_10000110_0;
      patterns[6257] = 25'b00011000_01101111_10000111_0;
      patterns[6258] = 25'b00011000_01110000_10001000_0;
      patterns[6259] = 25'b00011000_01110001_10001001_0;
      patterns[6260] = 25'b00011000_01110010_10001010_0;
      patterns[6261] = 25'b00011000_01110011_10001011_0;
      patterns[6262] = 25'b00011000_01110100_10001100_0;
      patterns[6263] = 25'b00011000_01110101_10001101_0;
      patterns[6264] = 25'b00011000_01110110_10001110_0;
      patterns[6265] = 25'b00011000_01110111_10001111_0;
      patterns[6266] = 25'b00011000_01111000_10010000_0;
      patterns[6267] = 25'b00011000_01111001_10010001_0;
      patterns[6268] = 25'b00011000_01111010_10010010_0;
      patterns[6269] = 25'b00011000_01111011_10010011_0;
      patterns[6270] = 25'b00011000_01111100_10010100_0;
      patterns[6271] = 25'b00011000_01111101_10010101_0;
      patterns[6272] = 25'b00011000_01111110_10010110_0;
      patterns[6273] = 25'b00011000_01111111_10010111_0;
      patterns[6274] = 25'b00011000_10000000_10011000_0;
      patterns[6275] = 25'b00011000_10000001_10011001_0;
      patterns[6276] = 25'b00011000_10000010_10011010_0;
      patterns[6277] = 25'b00011000_10000011_10011011_0;
      patterns[6278] = 25'b00011000_10000100_10011100_0;
      patterns[6279] = 25'b00011000_10000101_10011101_0;
      patterns[6280] = 25'b00011000_10000110_10011110_0;
      patterns[6281] = 25'b00011000_10000111_10011111_0;
      patterns[6282] = 25'b00011000_10001000_10100000_0;
      patterns[6283] = 25'b00011000_10001001_10100001_0;
      patterns[6284] = 25'b00011000_10001010_10100010_0;
      patterns[6285] = 25'b00011000_10001011_10100011_0;
      patterns[6286] = 25'b00011000_10001100_10100100_0;
      patterns[6287] = 25'b00011000_10001101_10100101_0;
      patterns[6288] = 25'b00011000_10001110_10100110_0;
      patterns[6289] = 25'b00011000_10001111_10100111_0;
      patterns[6290] = 25'b00011000_10010000_10101000_0;
      patterns[6291] = 25'b00011000_10010001_10101001_0;
      patterns[6292] = 25'b00011000_10010010_10101010_0;
      patterns[6293] = 25'b00011000_10010011_10101011_0;
      patterns[6294] = 25'b00011000_10010100_10101100_0;
      patterns[6295] = 25'b00011000_10010101_10101101_0;
      patterns[6296] = 25'b00011000_10010110_10101110_0;
      patterns[6297] = 25'b00011000_10010111_10101111_0;
      patterns[6298] = 25'b00011000_10011000_10110000_0;
      patterns[6299] = 25'b00011000_10011001_10110001_0;
      patterns[6300] = 25'b00011000_10011010_10110010_0;
      patterns[6301] = 25'b00011000_10011011_10110011_0;
      patterns[6302] = 25'b00011000_10011100_10110100_0;
      patterns[6303] = 25'b00011000_10011101_10110101_0;
      patterns[6304] = 25'b00011000_10011110_10110110_0;
      patterns[6305] = 25'b00011000_10011111_10110111_0;
      patterns[6306] = 25'b00011000_10100000_10111000_0;
      patterns[6307] = 25'b00011000_10100001_10111001_0;
      patterns[6308] = 25'b00011000_10100010_10111010_0;
      patterns[6309] = 25'b00011000_10100011_10111011_0;
      patterns[6310] = 25'b00011000_10100100_10111100_0;
      patterns[6311] = 25'b00011000_10100101_10111101_0;
      patterns[6312] = 25'b00011000_10100110_10111110_0;
      patterns[6313] = 25'b00011000_10100111_10111111_0;
      patterns[6314] = 25'b00011000_10101000_11000000_0;
      patterns[6315] = 25'b00011000_10101001_11000001_0;
      patterns[6316] = 25'b00011000_10101010_11000010_0;
      patterns[6317] = 25'b00011000_10101011_11000011_0;
      patterns[6318] = 25'b00011000_10101100_11000100_0;
      patterns[6319] = 25'b00011000_10101101_11000101_0;
      patterns[6320] = 25'b00011000_10101110_11000110_0;
      patterns[6321] = 25'b00011000_10101111_11000111_0;
      patterns[6322] = 25'b00011000_10110000_11001000_0;
      patterns[6323] = 25'b00011000_10110001_11001001_0;
      patterns[6324] = 25'b00011000_10110010_11001010_0;
      patterns[6325] = 25'b00011000_10110011_11001011_0;
      patterns[6326] = 25'b00011000_10110100_11001100_0;
      patterns[6327] = 25'b00011000_10110101_11001101_0;
      patterns[6328] = 25'b00011000_10110110_11001110_0;
      patterns[6329] = 25'b00011000_10110111_11001111_0;
      patterns[6330] = 25'b00011000_10111000_11010000_0;
      patterns[6331] = 25'b00011000_10111001_11010001_0;
      patterns[6332] = 25'b00011000_10111010_11010010_0;
      patterns[6333] = 25'b00011000_10111011_11010011_0;
      patterns[6334] = 25'b00011000_10111100_11010100_0;
      patterns[6335] = 25'b00011000_10111101_11010101_0;
      patterns[6336] = 25'b00011000_10111110_11010110_0;
      patterns[6337] = 25'b00011000_10111111_11010111_0;
      patterns[6338] = 25'b00011000_11000000_11011000_0;
      patterns[6339] = 25'b00011000_11000001_11011001_0;
      patterns[6340] = 25'b00011000_11000010_11011010_0;
      patterns[6341] = 25'b00011000_11000011_11011011_0;
      patterns[6342] = 25'b00011000_11000100_11011100_0;
      patterns[6343] = 25'b00011000_11000101_11011101_0;
      patterns[6344] = 25'b00011000_11000110_11011110_0;
      patterns[6345] = 25'b00011000_11000111_11011111_0;
      patterns[6346] = 25'b00011000_11001000_11100000_0;
      patterns[6347] = 25'b00011000_11001001_11100001_0;
      patterns[6348] = 25'b00011000_11001010_11100010_0;
      patterns[6349] = 25'b00011000_11001011_11100011_0;
      patterns[6350] = 25'b00011000_11001100_11100100_0;
      patterns[6351] = 25'b00011000_11001101_11100101_0;
      patterns[6352] = 25'b00011000_11001110_11100110_0;
      patterns[6353] = 25'b00011000_11001111_11100111_0;
      patterns[6354] = 25'b00011000_11010000_11101000_0;
      patterns[6355] = 25'b00011000_11010001_11101001_0;
      patterns[6356] = 25'b00011000_11010010_11101010_0;
      patterns[6357] = 25'b00011000_11010011_11101011_0;
      patterns[6358] = 25'b00011000_11010100_11101100_0;
      patterns[6359] = 25'b00011000_11010101_11101101_0;
      patterns[6360] = 25'b00011000_11010110_11101110_0;
      patterns[6361] = 25'b00011000_11010111_11101111_0;
      patterns[6362] = 25'b00011000_11011000_11110000_0;
      patterns[6363] = 25'b00011000_11011001_11110001_0;
      patterns[6364] = 25'b00011000_11011010_11110010_0;
      patterns[6365] = 25'b00011000_11011011_11110011_0;
      patterns[6366] = 25'b00011000_11011100_11110100_0;
      patterns[6367] = 25'b00011000_11011101_11110101_0;
      patterns[6368] = 25'b00011000_11011110_11110110_0;
      patterns[6369] = 25'b00011000_11011111_11110111_0;
      patterns[6370] = 25'b00011000_11100000_11111000_0;
      patterns[6371] = 25'b00011000_11100001_11111001_0;
      patterns[6372] = 25'b00011000_11100010_11111010_0;
      patterns[6373] = 25'b00011000_11100011_11111011_0;
      patterns[6374] = 25'b00011000_11100100_11111100_0;
      patterns[6375] = 25'b00011000_11100101_11111101_0;
      patterns[6376] = 25'b00011000_11100110_11111110_0;
      patterns[6377] = 25'b00011000_11100111_11111111_0;
      patterns[6378] = 25'b00011000_11101000_00000000_1;
      patterns[6379] = 25'b00011000_11101001_00000001_1;
      patterns[6380] = 25'b00011000_11101010_00000010_1;
      patterns[6381] = 25'b00011000_11101011_00000011_1;
      patterns[6382] = 25'b00011000_11101100_00000100_1;
      patterns[6383] = 25'b00011000_11101101_00000101_1;
      patterns[6384] = 25'b00011000_11101110_00000110_1;
      patterns[6385] = 25'b00011000_11101111_00000111_1;
      patterns[6386] = 25'b00011000_11110000_00001000_1;
      patterns[6387] = 25'b00011000_11110001_00001001_1;
      patterns[6388] = 25'b00011000_11110010_00001010_1;
      patterns[6389] = 25'b00011000_11110011_00001011_1;
      patterns[6390] = 25'b00011000_11110100_00001100_1;
      patterns[6391] = 25'b00011000_11110101_00001101_1;
      patterns[6392] = 25'b00011000_11110110_00001110_1;
      patterns[6393] = 25'b00011000_11110111_00001111_1;
      patterns[6394] = 25'b00011000_11111000_00010000_1;
      patterns[6395] = 25'b00011000_11111001_00010001_1;
      patterns[6396] = 25'b00011000_11111010_00010010_1;
      patterns[6397] = 25'b00011000_11111011_00010011_1;
      patterns[6398] = 25'b00011000_11111100_00010100_1;
      patterns[6399] = 25'b00011000_11111101_00010101_1;
      patterns[6400] = 25'b00011000_11111110_00010110_1;
      patterns[6401] = 25'b00011000_11111111_00010111_1;
      patterns[6402] = 25'b00011001_00000000_00011001_0;
      patterns[6403] = 25'b00011001_00000001_00011010_0;
      patterns[6404] = 25'b00011001_00000010_00011011_0;
      patterns[6405] = 25'b00011001_00000011_00011100_0;
      patterns[6406] = 25'b00011001_00000100_00011101_0;
      patterns[6407] = 25'b00011001_00000101_00011110_0;
      patterns[6408] = 25'b00011001_00000110_00011111_0;
      patterns[6409] = 25'b00011001_00000111_00100000_0;
      patterns[6410] = 25'b00011001_00001000_00100001_0;
      patterns[6411] = 25'b00011001_00001001_00100010_0;
      patterns[6412] = 25'b00011001_00001010_00100011_0;
      patterns[6413] = 25'b00011001_00001011_00100100_0;
      patterns[6414] = 25'b00011001_00001100_00100101_0;
      patterns[6415] = 25'b00011001_00001101_00100110_0;
      patterns[6416] = 25'b00011001_00001110_00100111_0;
      patterns[6417] = 25'b00011001_00001111_00101000_0;
      patterns[6418] = 25'b00011001_00010000_00101001_0;
      patterns[6419] = 25'b00011001_00010001_00101010_0;
      patterns[6420] = 25'b00011001_00010010_00101011_0;
      patterns[6421] = 25'b00011001_00010011_00101100_0;
      patterns[6422] = 25'b00011001_00010100_00101101_0;
      patterns[6423] = 25'b00011001_00010101_00101110_0;
      patterns[6424] = 25'b00011001_00010110_00101111_0;
      patterns[6425] = 25'b00011001_00010111_00110000_0;
      patterns[6426] = 25'b00011001_00011000_00110001_0;
      patterns[6427] = 25'b00011001_00011001_00110010_0;
      patterns[6428] = 25'b00011001_00011010_00110011_0;
      patterns[6429] = 25'b00011001_00011011_00110100_0;
      patterns[6430] = 25'b00011001_00011100_00110101_0;
      patterns[6431] = 25'b00011001_00011101_00110110_0;
      patterns[6432] = 25'b00011001_00011110_00110111_0;
      patterns[6433] = 25'b00011001_00011111_00111000_0;
      patterns[6434] = 25'b00011001_00100000_00111001_0;
      patterns[6435] = 25'b00011001_00100001_00111010_0;
      patterns[6436] = 25'b00011001_00100010_00111011_0;
      patterns[6437] = 25'b00011001_00100011_00111100_0;
      patterns[6438] = 25'b00011001_00100100_00111101_0;
      patterns[6439] = 25'b00011001_00100101_00111110_0;
      patterns[6440] = 25'b00011001_00100110_00111111_0;
      patterns[6441] = 25'b00011001_00100111_01000000_0;
      patterns[6442] = 25'b00011001_00101000_01000001_0;
      patterns[6443] = 25'b00011001_00101001_01000010_0;
      patterns[6444] = 25'b00011001_00101010_01000011_0;
      patterns[6445] = 25'b00011001_00101011_01000100_0;
      patterns[6446] = 25'b00011001_00101100_01000101_0;
      patterns[6447] = 25'b00011001_00101101_01000110_0;
      patterns[6448] = 25'b00011001_00101110_01000111_0;
      patterns[6449] = 25'b00011001_00101111_01001000_0;
      patterns[6450] = 25'b00011001_00110000_01001001_0;
      patterns[6451] = 25'b00011001_00110001_01001010_0;
      patterns[6452] = 25'b00011001_00110010_01001011_0;
      patterns[6453] = 25'b00011001_00110011_01001100_0;
      patterns[6454] = 25'b00011001_00110100_01001101_0;
      patterns[6455] = 25'b00011001_00110101_01001110_0;
      patterns[6456] = 25'b00011001_00110110_01001111_0;
      patterns[6457] = 25'b00011001_00110111_01010000_0;
      patterns[6458] = 25'b00011001_00111000_01010001_0;
      patterns[6459] = 25'b00011001_00111001_01010010_0;
      patterns[6460] = 25'b00011001_00111010_01010011_0;
      patterns[6461] = 25'b00011001_00111011_01010100_0;
      patterns[6462] = 25'b00011001_00111100_01010101_0;
      patterns[6463] = 25'b00011001_00111101_01010110_0;
      patterns[6464] = 25'b00011001_00111110_01010111_0;
      patterns[6465] = 25'b00011001_00111111_01011000_0;
      patterns[6466] = 25'b00011001_01000000_01011001_0;
      patterns[6467] = 25'b00011001_01000001_01011010_0;
      patterns[6468] = 25'b00011001_01000010_01011011_0;
      patterns[6469] = 25'b00011001_01000011_01011100_0;
      patterns[6470] = 25'b00011001_01000100_01011101_0;
      patterns[6471] = 25'b00011001_01000101_01011110_0;
      patterns[6472] = 25'b00011001_01000110_01011111_0;
      patterns[6473] = 25'b00011001_01000111_01100000_0;
      patterns[6474] = 25'b00011001_01001000_01100001_0;
      patterns[6475] = 25'b00011001_01001001_01100010_0;
      patterns[6476] = 25'b00011001_01001010_01100011_0;
      patterns[6477] = 25'b00011001_01001011_01100100_0;
      patterns[6478] = 25'b00011001_01001100_01100101_0;
      patterns[6479] = 25'b00011001_01001101_01100110_0;
      patterns[6480] = 25'b00011001_01001110_01100111_0;
      patterns[6481] = 25'b00011001_01001111_01101000_0;
      patterns[6482] = 25'b00011001_01010000_01101001_0;
      patterns[6483] = 25'b00011001_01010001_01101010_0;
      patterns[6484] = 25'b00011001_01010010_01101011_0;
      patterns[6485] = 25'b00011001_01010011_01101100_0;
      patterns[6486] = 25'b00011001_01010100_01101101_0;
      patterns[6487] = 25'b00011001_01010101_01101110_0;
      patterns[6488] = 25'b00011001_01010110_01101111_0;
      patterns[6489] = 25'b00011001_01010111_01110000_0;
      patterns[6490] = 25'b00011001_01011000_01110001_0;
      patterns[6491] = 25'b00011001_01011001_01110010_0;
      patterns[6492] = 25'b00011001_01011010_01110011_0;
      patterns[6493] = 25'b00011001_01011011_01110100_0;
      patterns[6494] = 25'b00011001_01011100_01110101_0;
      patterns[6495] = 25'b00011001_01011101_01110110_0;
      patterns[6496] = 25'b00011001_01011110_01110111_0;
      patterns[6497] = 25'b00011001_01011111_01111000_0;
      patterns[6498] = 25'b00011001_01100000_01111001_0;
      patterns[6499] = 25'b00011001_01100001_01111010_0;
      patterns[6500] = 25'b00011001_01100010_01111011_0;
      patterns[6501] = 25'b00011001_01100011_01111100_0;
      patterns[6502] = 25'b00011001_01100100_01111101_0;
      patterns[6503] = 25'b00011001_01100101_01111110_0;
      patterns[6504] = 25'b00011001_01100110_01111111_0;
      patterns[6505] = 25'b00011001_01100111_10000000_0;
      patterns[6506] = 25'b00011001_01101000_10000001_0;
      patterns[6507] = 25'b00011001_01101001_10000010_0;
      patterns[6508] = 25'b00011001_01101010_10000011_0;
      patterns[6509] = 25'b00011001_01101011_10000100_0;
      patterns[6510] = 25'b00011001_01101100_10000101_0;
      patterns[6511] = 25'b00011001_01101101_10000110_0;
      patterns[6512] = 25'b00011001_01101110_10000111_0;
      patterns[6513] = 25'b00011001_01101111_10001000_0;
      patterns[6514] = 25'b00011001_01110000_10001001_0;
      patterns[6515] = 25'b00011001_01110001_10001010_0;
      patterns[6516] = 25'b00011001_01110010_10001011_0;
      patterns[6517] = 25'b00011001_01110011_10001100_0;
      patterns[6518] = 25'b00011001_01110100_10001101_0;
      patterns[6519] = 25'b00011001_01110101_10001110_0;
      patterns[6520] = 25'b00011001_01110110_10001111_0;
      patterns[6521] = 25'b00011001_01110111_10010000_0;
      patterns[6522] = 25'b00011001_01111000_10010001_0;
      patterns[6523] = 25'b00011001_01111001_10010010_0;
      patterns[6524] = 25'b00011001_01111010_10010011_0;
      patterns[6525] = 25'b00011001_01111011_10010100_0;
      patterns[6526] = 25'b00011001_01111100_10010101_0;
      patterns[6527] = 25'b00011001_01111101_10010110_0;
      patterns[6528] = 25'b00011001_01111110_10010111_0;
      patterns[6529] = 25'b00011001_01111111_10011000_0;
      patterns[6530] = 25'b00011001_10000000_10011001_0;
      patterns[6531] = 25'b00011001_10000001_10011010_0;
      patterns[6532] = 25'b00011001_10000010_10011011_0;
      patterns[6533] = 25'b00011001_10000011_10011100_0;
      patterns[6534] = 25'b00011001_10000100_10011101_0;
      patterns[6535] = 25'b00011001_10000101_10011110_0;
      patterns[6536] = 25'b00011001_10000110_10011111_0;
      patterns[6537] = 25'b00011001_10000111_10100000_0;
      patterns[6538] = 25'b00011001_10001000_10100001_0;
      patterns[6539] = 25'b00011001_10001001_10100010_0;
      patterns[6540] = 25'b00011001_10001010_10100011_0;
      patterns[6541] = 25'b00011001_10001011_10100100_0;
      patterns[6542] = 25'b00011001_10001100_10100101_0;
      patterns[6543] = 25'b00011001_10001101_10100110_0;
      patterns[6544] = 25'b00011001_10001110_10100111_0;
      patterns[6545] = 25'b00011001_10001111_10101000_0;
      patterns[6546] = 25'b00011001_10010000_10101001_0;
      patterns[6547] = 25'b00011001_10010001_10101010_0;
      patterns[6548] = 25'b00011001_10010010_10101011_0;
      patterns[6549] = 25'b00011001_10010011_10101100_0;
      patterns[6550] = 25'b00011001_10010100_10101101_0;
      patterns[6551] = 25'b00011001_10010101_10101110_0;
      patterns[6552] = 25'b00011001_10010110_10101111_0;
      patterns[6553] = 25'b00011001_10010111_10110000_0;
      patterns[6554] = 25'b00011001_10011000_10110001_0;
      patterns[6555] = 25'b00011001_10011001_10110010_0;
      patterns[6556] = 25'b00011001_10011010_10110011_0;
      patterns[6557] = 25'b00011001_10011011_10110100_0;
      patterns[6558] = 25'b00011001_10011100_10110101_0;
      patterns[6559] = 25'b00011001_10011101_10110110_0;
      patterns[6560] = 25'b00011001_10011110_10110111_0;
      patterns[6561] = 25'b00011001_10011111_10111000_0;
      patterns[6562] = 25'b00011001_10100000_10111001_0;
      patterns[6563] = 25'b00011001_10100001_10111010_0;
      patterns[6564] = 25'b00011001_10100010_10111011_0;
      patterns[6565] = 25'b00011001_10100011_10111100_0;
      patterns[6566] = 25'b00011001_10100100_10111101_0;
      patterns[6567] = 25'b00011001_10100101_10111110_0;
      patterns[6568] = 25'b00011001_10100110_10111111_0;
      patterns[6569] = 25'b00011001_10100111_11000000_0;
      patterns[6570] = 25'b00011001_10101000_11000001_0;
      patterns[6571] = 25'b00011001_10101001_11000010_0;
      patterns[6572] = 25'b00011001_10101010_11000011_0;
      patterns[6573] = 25'b00011001_10101011_11000100_0;
      patterns[6574] = 25'b00011001_10101100_11000101_0;
      patterns[6575] = 25'b00011001_10101101_11000110_0;
      patterns[6576] = 25'b00011001_10101110_11000111_0;
      patterns[6577] = 25'b00011001_10101111_11001000_0;
      patterns[6578] = 25'b00011001_10110000_11001001_0;
      patterns[6579] = 25'b00011001_10110001_11001010_0;
      patterns[6580] = 25'b00011001_10110010_11001011_0;
      patterns[6581] = 25'b00011001_10110011_11001100_0;
      patterns[6582] = 25'b00011001_10110100_11001101_0;
      patterns[6583] = 25'b00011001_10110101_11001110_0;
      patterns[6584] = 25'b00011001_10110110_11001111_0;
      patterns[6585] = 25'b00011001_10110111_11010000_0;
      patterns[6586] = 25'b00011001_10111000_11010001_0;
      patterns[6587] = 25'b00011001_10111001_11010010_0;
      patterns[6588] = 25'b00011001_10111010_11010011_0;
      patterns[6589] = 25'b00011001_10111011_11010100_0;
      patterns[6590] = 25'b00011001_10111100_11010101_0;
      patterns[6591] = 25'b00011001_10111101_11010110_0;
      patterns[6592] = 25'b00011001_10111110_11010111_0;
      patterns[6593] = 25'b00011001_10111111_11011000_0;
      patterns[6594] = 25'b00011001_11000000_11011001_0;
      patterns[6595] = 25'b00011001_11000001_11011010_0;
      patterns[6596] = 25'b00011001_11000010_11011011_0;
      patterns[6597] = 25'b00011001_11000011_11011100_0;
      patterns[6598] = 25'b00011001_11000100_11011101_0;
      patterns[6599] = 25'b00011001_11000101_11011110_0;
      patterns[6600] = 25'b00011001_11000110_11011111_0;
      patterns[6601] = 25'b00011001_11000111_11100000_0;
      patterns[6602] = 25'b00011001_11001000_11100001_0;
      patterns[6603] = 25'b00011001_11001001_11100010_0;
      patterns[6604] = 25'b00011001_11001010_11100011_0;
      patterns[6605] = 25'b00011001_11001011_11100100_0;
      patterns[6606] = 25'b00011001_11001100_11100101_0;
      patterns[6607] = 25'b00011001_11001101_11100110_0;
      patterns[6608] = 25'b00011001_11001110_11100111_0;
      patterns[6609] = 25'b00011001_11001111_11101000_0;
      patterns[6610] = 25'b00011001_11010000_11101001_0;
      patterns[6611] = 25'b00011001_11010001_11101010_0;
      patterns[6612] = 25'b00011001_11010010_11101011_0;
      patterns[6613] = 25'b00011001_11010011_11101100_0;
      patterns[6614] = 25'b00011001_11010100_11101101_0;
      patterns[6615] = 25'b00011001_11010101_11101110_0;
      patterns[6616] = 25'b00011001_11010110_11101111_0;
      patterns[6617] = 25'b00011001_11010111_11110000_0;
      patterns[6618] = 25'b00011001_11011000_11110001_0;
      patterns[6619] = 25'b00011001_11011001_11110010_0;
      patterns[6620] = 25'b00011001_11011010_11110011_0;
      patterns[6621] = 25'b00011001_11011011_11110100_0;
      patterns[6622] = 25'b00011001_11011100_11110101_0;
      patterns[6623] = 25'b00011001_11011101_11110110_0;
      patterns[6624] = 25'b00011001_11011110_11110111_0;
      patterns[6625] = 25'b00011001_11011111_11111000_0;
      patterns[6626] = 25'b00011001_11100000_11111001_0;
      patterns[6627] = 25'b00011001_11100001_11111010_0;
      patterns[6628] = 25'b00011001_11100010_11111011_0;
      patterns[6629] = 25'b00011001_11100011_11111100_0;
      patterns[6630] = 25'b00011001_11100100_11111101_0;
      patterns[6631] = 25'b00011001_11100101_11111110_0;
      patterns[6632] = 25'b00011001_11100110_11111111_0;
      patterns[6633] = 25'b00011001_11100111_00000000_1;
      patterns[6634] = 25'b00011001_11101000_00000001_1;
      patterns[6635] = 25'b00011001_11101001_00000010_1;
      patterns[6636] = 25'b00011001_11101010_00000011_1;
      patterns[6637] = 25'b00011001_11101011_00000100_1;
      patterns[6638] = 25'b00011001_11101100_00000101_1;
      patterns[6639] = 25'b00011001_11101101_00000110_1;
      patterns[6640] = 25'b00011001_11101110_00000111_1;
      patterns[6641] = 25'b00011001_11101111_00001000_1;
      patterns[6642] = 25'b00011001_11110000_00001001_1;
      patterns[6643] = 25'b00011001_11110001_00001010_1;
      patterns[6644] = 25'b00011001_11110010_00001011_1;
      patterns[6645] = 25'b00011001_11110011_00001100_1;
      patterns[6646] = 25'b00011001_11110100_00001101_1;
      patterns[6647] = 25'b00011001_11110101_00001110_1;
      patterns[6648] = 25'b00011001_11110110_00001111_1;
      patterns[6649] = 25'b00011001_11110111_00010000_1;
      patterns[6650] = 25'b00011001_11111000_00010001_1;
      patterns[6651] = 25'b00011001_11111001_00010010_1;
      patterns[6652] = 25'b00011001_11111010_00010011_1;
      patterns[6653] = 25'b00011001_11111011_00010100_1;
      patterns[6654] = 25'b00011001_11111100_00010101_1;
      patterns[6655] = 25'b00011001_11111101_00010110_1;
      patterns[6656] = 25'b00011001_11111110_00010111_1;
      patterns[6657] = 25'b00011001_11111111_00011000_1;
      patterns[6658] = 25'b00011010_00000000_00011010_0;
      patterns[6659] = 25'b00011010_00000001_00011011_0;
      patterns[6660] = 25'b00011010_00000010_00011100_0;
      patterns[6661] = 25'b00011010_00000011_00011101_0;
      patterns[6662] = 25'b00011010_00000100_00011110_0;
      patterns[6663] = 25'b00011010_00000101_00011111_0;
      patterns[6664] = 25'b00011010_00000110_00100000_0;
      patterns[6665] = 25'b00011010_00000111_00100001_0;
      patterns[6666] = 25'b00011010_00001000_00100010_0;
      patterns[6667] = 25'b00011010_00001001_00100011_0;
      patterns[6668] = 25'b00011010_00001010_00100100_0;
      patterns[6669] = 25'b00011010_00001011_00100101_0;
      patterns[6670] = 25'b00011010_00001100_00100110_0;
      patterns[6671] = 25'b00011010_00001101_00100111_0;
      patterns[6672] = 25'b00011010_00001110_00101000_0;
      patterns[6673] = 25'b00011010_00001111_00101001_0;
      patterns[6674] = 25'b00011010_00010000_00101010_0;
      patterns[6675] = 25'b00011010_00010001_00101011_0;
      patterns[6676] = 25'b00011010_00010010_00101100_0;
      patterns[6677] = 25'b00011010_00010011_00101101_0;
      patterns[6678] = 25'b00011010_00010100_00101110_0;
      patterns[6679] = 25'b00011010_00010101_00101111_0;
      patterns[6680] = 25'b00011010_00010110_00110000_0;
      patterns[6681] = 25'b00011010_00010111_00110001_0;
      patterns[6682] = 25'b00011010_00011000_00110010_0;
      patterns[6683] = 25'b00011010_00011001_00110011_0;
      patterns[6684] = 25'b00011010_00011010_00110100_0;
      patterns[6685] = 25'b00011010_00011011_00110101_0;
      patterns[6686] = 25'b00011010_00011100_00110110_0;
      patterns[6687] = 25'b00011010_00011101_00110111_0;
      patterns[6688] = 25'b00011010_00011110_00111000_0;
      patterns[6689] = 25'b00011010_00011111_00111001_0;
      patterns[6690] = 25'b00011010_00100000_00111010_0;
      patterns[6691] = 25'b00011010_00100001_00111011_0;
      patterns[6692] = 25'b00011010_00100010_00111100_0;
      patterns[6693] = 25'b00011010_00100011_00111101_0;
      patterns[6694] = 25'b00011010_00100100_00111110_0;
      patterns[6695] = 25'b00011010_00100101_00111111_0;
      patterns[6696] = 25'b00011010_00100110_01000000_0;
      patterns[6697] = 25'b00011010_00100111_01000001_0;
      patterns[6698] = 25'b00011010_00101000_01000010_0;
      patterns[6699] = 25'b00011010_00101001_01000011_0;
      patterns[6700] = 25'b00011010_00101010_01000100_0;
      patterns[6701] = 25'b00011010_00101011_01000101_0;
      patterns[6702] = 25'b00011010_00101100_01000110_0;
      patterns[6703] = 25'b00011010_00101101_01000111_0;
      patterns[6704] = 25'b00011010_00101110_01001000_0;
      patterns[6705] = 25'b00011010_00101111_01001001_0;
      patterns[6706] = 25'b00011010_00110000_01001010_0;
      patterns[6707] = 25'b00011010_00110001_01001011_0;
      patterns[6708] = 25'b00011010_00110010_01001100_0;
      patterns[6709] = 25'b00011010_00110011_01001101_0;
      patterns[6710] = 25'b00011010_00110100_01001110_0;
      patterns[6711] = 25'b00011010_00110101_01001111_0;
      patterns[6712] = 25'b00011010_00110110_01010000_0;
      patterns[6713] = 25'b00011010_00110111_01010001_0;
      patterns[6714] = 25'b00011010_00111000_01010010_0;
      patterns[6715] = 25'b00011010_00111001_01010011_0;
      patterns[6716] = 25'b00011010_00111010_01010100_0;
      patterns[6717] = 25'b00011010_00111011_01010101_0;
      patterns[6718] = 25'b00011010_00111100_01010110_0;
      patterns[6719] = 25'b00011010_00111101_01010111_0;
      patterns[6720] = 25'b00011010_00111110_01011000_0;
      patterns[6721] = 25'b00011010_00111111_01011001_0;
      patterns[6722] = 25'b00011010_01000000_01011010_0;
      patterns[6723] = 25'b00011010_01000001_01011011_0;
      patterns[6724] = 25'b00011010_01000010_01011100_0;
      patterns[6725] = 25'b00011010_01000011_01011101_0;
      patterns[6726] = 25'b00011010_01000100_01011110_0;
      patterns[6727] = 25'b00011010_01000101_01011111_0;
      patterns[6728] = 25'b00011010_01000110_01100000_0;
      patterns[6729] = 25'b00011010_01000111_01100001_0;
      patterns[6730] = 25'b00011010_01001000_01100010_0;
      patterns[6731] = 25'b00011010_01001001_01100011_0;
      patterns[6732] = 25'b00011010_01001010_01100100_0;
      patterns[6733] = 25'b00011010_01001011_01100101_0;
      patterns[6734] = 25'b00011010_01001100_01100110_0;
      patterns[6735] = 25'b00011010_01001101_01100111_0;
      patterns[6736] = 25'b00011010_01001110_01101000_0;
      patterns[6737] = 25'b00011010_01001111_01101001_0;
      patterns[6738] = 25'b00011010_01010000_01101010_0;
      patterns[6739] = 25'b00011010_01010001_01101011_0;
      patterns[6740] = 25'b00011010_01010010_01101100_0;
      patterns[6741] = 25'b00011010_01010011_01101101_0;
      patterns[6742] = 25'b00011010_01010100_01101110_0;
      patterns[6743] = 25'b00011010_01010101_01101111_0;
      patterns[6744] = 25'b00011010_01010110_01110000_0;
      patterns[6745] = 25'b00011010_01010111_01110001_0;
      patterns[6746] = 25'b00011010_01011000_01110010_0;
      patterns[6747] = 25'b00011010_01011001_01110011_0;
      patterns[6748] = 25'b00011010_01011010_01110100_0;
      patterns[6749] = 25'b00011010_01011011_01110101_0;
      patterns[6750] = 25'b00011010_01011100_01110110_0;
      patterns[6751] = 25'b00011010_01011101_01110111_0;
      patterns[6752] = 25'b00011010_01011110_01111000_0;
      patterns[6753] = 25'b00011010_01011111_01111001_0;
      patterns[6754] = 25'b00011010_01100000_01111010_0;
      patterns[6755] = 25'b00011010_01100001_01111011_0;
      patterns[6756] = 25'b00011010_01100010_01111100_0;
      patterns[6757] = 25'b00011010_01100011_01111101_0;
      patterns[6758] = 25'b00011010_01100100_01111110_0;
      patterns[6759] = 25'b00011010_01100101_01111111_0;
      patterns[6760] = 25'b00011010_01100110_10000000_0;
      patterns[6761] = 25'b00011010_01100111_10000001_0;
      patterns[6762] = 25'b00011010_01101000_10000010_0;
      patterns[6763] = 25'b00011010_01101001_10000011_0;
      patterns[6764] = 25'b00011010_01101010_10000100_0;
      patterns[6765] = 25'b00011010_01101011_10000101_0;
      patterns[6766] = 25'b00011010_01101100_10000110_0;
      patterns[6767] = 25'b00011010_01101101_10000111_0;
      patterns[6768] = 25'b00011010_01101110_10001000_0;
      patterns[6769] = 25'b00011010_01101111_10001001_0;
      patterns[6770] = 25'b00011010_01110000_10001010_0;
      patterns[6771] = 25'b00011010_01110001_10001011_0;
      patterns[6772] = 25'b00011010_01110010_10001100_0;
      patterns[6773] = 25'b00011010_01110011_10001101_0;
      patterns[6774] = 25'b00011010_01110100_10001110_0;
      patterns[6775] = 25'b00011010_01110101_10001111_0;
      patterns[6776] = 25'b00011010_01110110_10010000_0;
      patterns[6777] = 25'b00011010_01110111_10010001_0;
      patterns[6778] = 25'b00011010_01111000_10010010_0;
      patterns[6779] = 25'b00011010_01111001_10010011_0;
      patterns[6780] = 25'b00011010_01111010_10010100_0;
      patterns[6781] = 25'b00011010_01111011_10010101_0;
      patterns[6782] = 25'b00011010_01111100_10010110_0;
      patterns[6783] = 25'b00011010_01111101_10010111_0;
      patterns[6784] = 25'b00011010_01111110_10011000_0;
      patterns[6785] = 25'b00011010_01111111_10011001_0;
      patterns[6786] = 25'b00011010_10000000_10011010_0;
      patterns[6787] = 25'b00011010_10000001_10011011_0;
      patterns[6788] = 25'b00011010_10000010_10011100_0;
      patterns[6789] = 25'b00011010_10000011_10011101_0;
      patterns[6790] = 25'b00011010_10000100_10011110_0;
      patterns[6791] = 25'b00011010_10000101_10011111_0;
      patterns[6792] = 25'b00011010_10000110_10100000_0;
      patterns[6793] = 25'b00011010_10000111_10100001_0;
      patterns[6794] = 25'b00011010_10001000_10100010_0;
      patterns[6795] = 25'b00011010_10001001_10100011_0;
      patterns[6796] = 25'b00011010_10001010_10100100_0;
      patterns[6797] = 25'b00011010_10001011_10100101_0;
      patterns[6798] = 25'b00011010_10001100_10100110_0;
      patterns[6799] = 25'b00011010_10001101_10100111_0;
      patterns[6800] = 25'b00011010_10001110_10101000_0;
      patterns[6801] = 25'b00011010_10001111_10101001_0;
      patterns[6802] = 25'b00011010_10010000_10101010_0;
      patterns[6803] = 25'b00011010_10010001_10101011_0;
      patterns[6804] = 25'b00011010_10010010_10101100_0;
      patterns[6805] = 25'b00011010_10010011_10101101_0;
      patterns[6806] = 25'b00011010_10010100_10101110_0;
      patterns[6807] = 25'b00011010_10010101_10101111_0;
      patterns[6808] = 25'b00011010_10010110_10110000_0;
      patterns[6809] = 25'b00011010_10010111_10110001_0;
      patterns[6810] = 25'b00011010_10011000_10110010_0;
      patterns[6811] = 25'b00011010_10011001_10110011_0;
      patterns[6812] = 25'b00011010_10011010_10110100_0;
      patterns[6813] = 25'b00011010_10011011_10110101_0;
      patterns[6814] = 25'b00011010_10011100_10110110_0;
      patterns[6815] = 25'b00011010_10011101_10110111_0;
      patterns[6816] = 25'b00011010_10011110_10111000_0;
      patterns[6817] = 25'b00011010_10011111_10111001_0;
      patterns[6818] = 25'b00011010_10100000_10111010_0;
      patterns[6819] = 25'b00011010_10100001_10111011_0;
      patterns[6820] = 25'b00011010_10100010_10111100_0;
      patterns[6821] = 25'b00011010_10100011_10111101_0;
      patterns[6822] = 25'b00011010_10100100_10111110_0;
      patterns[6823] = 25'b00011010_10100101_10111111_0;
      patterns[6824] = 25'b00011010_10100110_11000000_0;
      patterns[6825] = 25'b00011010_10100111_11000001_0;
      patterns[6826] = 25'b00011010_10101000_11000010_0;
      patterns[6827] = 25'b00011010_10101001_11000011_0;
      patterns[6828] = 25'b00011010_10101010_11000100_0;
      patterns[6829] = 25'b00011010_10101011_11000101_0;
      patterns[6830] = 25'b00011010_10101100_11000110_0;
      patterns[6831] = 25'b00011010_10101101_11000111_0;
      patterns[6832] = 25'b00011010_10101110_11001000_0;
      patterns[6833] = 25'b00011010_10101111_11001001_0;
      patterns[6834] = 25'b00011010_10110000_11001010_0;
      patterns[6835] = 25'b00011010_10110001_11001011_0;
      patterns[6836] = 25'b00011010_10110010_11001100_0;
      patterns[6837] = 25'b00011010_10110011_11001101_0;
      patterns[6838] = 25'b00011010_10110100_11001110_0;
      patterns[6839] = 25'b00011010_10110101_11001111_0;
      patterns[6840] = 25'b00011010_10110110_11010000_0;
      patterns[6841] = 25'b00011010_10110111_11010001_0;
      patterns[6842] = 25'b00011010_10111000_11010010_0;
      patterns[6843] = 25'b00011010_10111001_11010011_0;
      patterns[6844] = 25'b00011010_10111010_11010100_0;
      patterns[6845] = 25'b00011010_10111011_11010101_0;
      patterns[6846] = 25'b00011010_10111100_11010110_0;
      patterns[6847] = 25'b00011010_10111101_11010111_0;
      patterns[6848] = 25'b00011010_10111110_11011000_0;
      patterns[6849] = 25'b00011010_10111111_11011001_0;
      patterns[6850] = 25'b00011010_11000000_11011010_0;
      patterns[6851] = 25'b00011010_11000001_11011011_0;
      patterns[6852] = 25'b00011010_11000010_11011100_0;
      patterns[6853] = 25'b00011010_11000011_11011101_0;
      patterns[6854] = 25'b00011010_11000100_11011110_0;
      patterns[6855] = 25'b00011010_11000101_11011111_0;
      patterns[6856] = 25'b00011010_11000110_11100000_0;
      patterns[6857] = 25'b00011010_11000111_11100001_0;
      patterns[6858] = 25'b00011010_11001000_11100010_0;
      patterns[6859] = 25'b00011010_11001001_11100011_0;
      patterns[6860] = 25'b00011010_11001010_11100100_0;
      patterns[6861] = 25'b00011010_11001011_11100101_0;
      patterns[6862] = 25'b00011010_11001100_11100110_0;
      patterns[6863] = 25'b00011010_11001101_11100111_0;
      patterns[6864] = 25'b00011010_11001110_11101000_0;
      patterns[6865] = 25'b00011010_11001111_11101001_0;
      patterns[6866] = 25'b00011010_11010000_11101010_0;
      patterns[6867] = 25'b00011010_11010001_11101011_0;
      patterns[6868] = 25'b00011010_11010010_11101100_0;
      patterns[6869] = 25'b00011010_11010011_11101101_0;
      patterns[6870] = 25'b00011010_11010100_11101110_0;
      patterns[6871] = 25'b00011010_11010101_11101111_0;
      patterns[6872] = 25'b00011010_11010110_11110000_0;
      patterns[6873] = 25'b00011010_11010111_11110001_0;
      patterns[6874] = 25'b00011010_11011000_11110010_0;
      patterns[6875] = 25'b00011010_11011001_11110011_0;
      patterns[6876] = 25'b00011010_11011010_11110100_0;
      patterns[6877] = 25'b00011010_11011011_11110101_0;
      patterns[6878] = 25'b00011010_11011100_11110110_0;
      patterns[6879] = 25'b00011010_11011101_11110111_0;
      patterns[6880] = 25'b00011010_11011110_11111000_0;
      patterns[6881] = 25'b00011010_11011111_11111001_0;
      patterns[6882] = 25'b00011010_11100000_11111010_0;
      patterns[6883] = 25'b00011010_11100001_11111011_0;
      patterns[6884] = 25'b00011010_11100010_11111100_0;
      patterns[6885] = 25'b00011010_11100011_11111101_0;
      patterns[6886] = 25'b00011010_11100100_11111110_0;
      patterns[6887] = 25'b00011010_11100101_11111111_0;
      patterns[6888] = 25'b00011010_11100110_00000000_1;
      patterns[6889] = 25'b00011010_11100111_00000001_1;
      patterns[6890] = 25'b00011010_11101000_00000010_1;
      patterns[6891] = 25'b00011010_11101001_00000011_1;
      patterns[6892] = 25'b00011010_11101010_00000100_1;
      patterns[6893] = 25'b00011010_11101011_00000101_1;
      patterns[6894] = 25'b00011010_11101100_00000110_1;
      patterns[6895] = 25'b00011010_11101101_00000111_1;
      patterns[6896] = 25'b00011010_11101110_00001000_1;
      patterns[6897] = 25'b00011010_11101111_00001001_1;
      patterns[6898] = 25'b00011010_11110000_00001010_1;
      patterns[6899] = 25'b00011010_11110001_00001011_1;
      patterns[6900] = 25'b00011010_11110010_00001100_1;
      patterns[6901] = 25'b00011010_11110011_00001101_1;
      patterns[6902] = 25'b00011010_11110100_00001110_1;
      patterns[6903] = 25'b00011010_11110101_00001111_1;
      patterns[6904] = 25'b00011010_11110110_00010000_1;
      patterns[6905] = 25'b00011010_11110111_00010001_1;
      patterns[6906] = 25'b00011010_11111000_00010010_1;
      patterns[6907] = 25'b00011010_11111001_00010011_1;
      patterns[6908] = 25'b00011010_11111010_00010100_1;
      patterns[6909] = 25'b00011010_11111011_00010101_1;
      patterns[6910] = 25'b00011010_11111100_00010110_1;
      patterns[6911] = 25'b00011010_11111101_00010111_1;
      patterns[6912] = 25'b00011010_11111110_00011000_1;
      patterns[6913] = 25'b00011010_11111111_00011001_1;
      patterns[6914] = 25'b00011011_00000000_00011011_0;
      patterns[6915] = 25'b00011011_00000001_00011100_0;
      patterns[6916] = 25'b00011011_00000010_00011101_0;
      patterns[6917] = 25'b00011011_00000011_00011110_0;
      patterns[6918] = 25'b00011011_00000100_00011111_0;
      patterns[6919] = 25'b00011011_00000101_00100000_0;
      patterns[6920] = 25'b00011011_00000110_00100001_0;
      patterns[6921] = 25'b00011011_00000111_00100010_0;
      patterns[6922] = 25'b00011011_00001000_00100011_0;
      patterns[6923] = 25'b00011011_00001001_00100100_0;
      patterns[6924] = 25'b00011011_00001010_00100101_0;
      patterns[6925] = 25'b00011011_00001011_00100110_0;
      patterns[6926] = 25'b00011011_00001100_00100111_0;
      patterns[6927] = 25'b00011011_00001101_00101000_0;
      patterns[6928] = 25'b00011011_00001110_00101001_0;
      patterns[6929] = 25'b00011011_00001111_00101010_0;
      patterns[6930] = 25'b00011011_00010000_00101011_0;
      patterns[6931] = 25'b00011011_00010001_00101100_0;
      patterns[6932] = 25'b00011011_00010010_00101101_0;
      patterns[6933] = 25'b00011011_00010011_00101110_0;
      patterns[6934] = 25'b00011011_00010100_00101111_0;
      patterns[6935] = 25'b00011011_00010101_00110000_0;
      patterns[6936] = 25'b00011011_00010110_00110001_0;
      patterns[6937] = 25'b00011011_00010111_00110010_0;
      patterns[6938] = 25'b00011011_00011000_00110011_0;
      patterns[6939] = 25'b00011011_00011001_00110100_0;
      patterns[6940] = 25'b00011011_00011010_00110101_0;
      patterns[6941] = 25'b00011011_00011011_00110110_0;
      patterns[6942] = 25'b00011011_00011100_00110111_0;
      patterns[6943] = 25'b00011011_00011101_00111000_0;
      patterns[6944] = 25'b00011011_00011110_00111001_0;
      patterns[6945] = 25'b00011011_00011111_00111010_0;
      patterns[6946] = 25'b00011011_00100000_00111011_0;
      patterns[6947] = 25'b00011011_00100001_00111100_0;
      patterns[6948] = 25'b00011011_00100010_00111101_0;
      patterns[6949] = 25'b00011011_00100011_00111110_0;
      patterns[6950] = 25'b00011011_00100100_00111111_0;
      patterns[6951] = 25'b00011011_00100101_01000000_0;
      patterns[6952] = 25'b00011011_00100110_01000001_0;
      patterns[6953] = 25'b00011011_00100111_01000010_0;
      patterns[6954] = 25'b00011011_00101000_01000011_0;
      patterns[6955] = 25'b00011011_00101001_01000100_0;
      patterns[6956] = 25'b00011011_00101010_01000101_0;
      patterns[6957] = 25'b00011011_00101011_01000110_0;
      patterns[6958] = 25'b00011011_00101100_01000111_0;
      patterns[6959] = 25'b00011011_00101101_01001000_0;
      patterns[6960] = 25'b00011011_00101110_01001001_0;
      patterns[6961] = 25'b00011011_00101111_01001010_0;
      patterns[6962] = 25'b00011011_00110000_01001011_0;
      patterns[6963] = 25'b00011011_00110001_01001100_0;
      patterns[6964] = 25'b00011011_00110010_01001101_0;
      patterns[6965] = 25'b00011011_00110011_01001110_0;
      patterns[6966] = 25'b00011011_00110100_01001111_0;
      patterns[6967] = 25'b00011011_00110101_01010000_0;
      patterns[6968] = 25'b00011011_00110110_01010001_0;
      patterns[6969] = 25'b00011011_00110111_01010010_0;
      patterns[6970] = 25'b00011011_00111000_01010011_0;
      patterns[6971] = 25'b00011011_00111001_01010100_0;
      patterns[6972] = 25'b00011011_00111010_01010101_0;
      patterns[6973] = 25'b00011011_00111011_01010110_0;
      patterns[6974] = 25'b00011011_00111100_01010111_0;
      patterns[6975] = 25'b00011011_00111101_01011000_0;
      patterns[6976] = 25'b00011011_00111110_01011001_0;
      patterns[6977] = 25'b00011011_00111111_01011010_0;
      patterns[6978] = 25'b00011011_01000000_01011011_0;
      patterns[6979] = 25'b00011011_01000001_01011100_0;
      patterns[6980] = 25'b00011011_01000010_01011101_0;
      patterns[6981] = 25'b00011011_01000011_01011110_0;
      patterns[6982] = 25'b00011011_01000100_01011111_0;
      patterns[6983] = 25'b00011011_01000101_01100000_0;
      patterns[6984] = 25'b00011011_01000110_01100001_0;
      patterns[6985] = 25'b00011011_01000111_01100010_0;
      patterns[6986] = 25'b00011011_01001000_01100011_0;
      patterns[6987] = 25'b00011011_01001001_01100100_0;
      patterns[6988] = 25'b00011011_01001010_01100101_0;
      patterns[6989] = 25'b00011011_01001011_01100110_0;
      patterns[6990] = 25'b00011011_01001100_01100111_0;
      patterns[6991] = 25'b00011011_01001101_01101000_0;
      patterns[6992] = 25'b00011011_01001110_01101001_0;
      patterns[6993] = 25'b00011011_01001111_01101010_0;
      patterns[6994] = 25'b00011011_01010000_01101011_0;
      patterns[6995] = 25'b00011011_01010001_01101100_0;
      patterns[6996] = 25'b00011011_01010010_01101101_0;
      patterns[6997] = 25'b00011011_01010011_01101110_0;
      patterns[6998] = 25'b00011011_01010100_01101111_0;
      patterns[6999] = 25'b00011011_01010101_01110000_0;
      patterns[7000] = 25'b00011011_01010110_01110001_0;
      patterns[7001] = 25'b00011011_01010111_01110010_0;
      patterns[7002] = 25'b00011011_01011000_01110011_0;
      patterns[7003] = 25'b00011011_01011001_01110100_0;
      patterns[7004] = 25'b00011011_01011010_01110101_0;
      patterns[7005] = 25'b00011011_01011011_01110110_0;
      patterns[7006] = 25'b00011011_01011100_01110111_0;
      patterns[7007] = 25'b00011011_01011101_01111000_0;
      patterns[7008] = 25'b00011011_01011110_01111001_0;
      patterns[7009] = 25'b00011011_01011111_01111010_0;
      patterns[7010] = 25'b00011011_01100000_01111011_0;
      patterns[7011] = 25'b00011011_01100001_01111100_0;
      patterns[7012] = 25'b00011011_01100010_01111101_0;
      patterns[7013] = 25'b00011011_01100011_01111110_0;
      patterns[7014] = 25'b00011011_01100100_01111111_0;
      patterns[7015] = 25'b00011011_01100101_10000000_0;
      patterns[7016] = 25'b00011011_01100110_10000001_0;
      patterns[7017] = 25'b00011011_01100111_10000010_0;
      patterns[7018] = 25'b00011011_01101000_10000011_0;
      patterns[7019] = 25'b00011011_01101001_10000100_0;
      patterns[7020] = 25'b00011011_01101010_10000101_0;
      patterns[7021] = 25'b00011011_01101011_10000110_0;
      patterns[7022] = 25'b00011011_01101100_10000111_0;
      patterns[7023] = 25'b00011011_01101101_10001000_0;
      patterns[7024] = 25'b00011011_01101110_10001001_0;
      patterns[7025] = 25'b00011011_01101111_10001010_0;
      patterns[7026] = 25'b00011011_01110000_10001011_0;
      patterns[7027] = 25'b00011011_01110001_10001100_0;
      patterns[7028] = 25'b00011011_01110010_10001101_0;
      patterns[7029] = 25'b00011011_01110011_10001110_0;
      patterns[7030] = 25'b00011011_01110100_10001111_0;
      patterns[7031] = 25'b00011011_01110101_10010000_0;
      patterns[7032] = 25'b00011011_01110110_10010001_0;
      patterns[7033] = 25'b00011011_01110111_10010010_0;
      patterns[7034] = 25'b00011011_01111000_10010011_0;
      patterns[7035] = 25'b00011011_01111001_10010100_0;
      patterns[7036] = 25'b00011011_01111010_10010101_0;
      patterns[7037] = 25'b00011011_01111011_10010110_0;
      patterns[7038] = 25'b00011011_01111100_10010111_0;
      patterns[7039] = 25'b00011011_01111101_10011000_0;
      patterns[7040] = 25'b00011011_01111110_10011001_0;
      patterns[7041] = 25'b00011011_01111111_10011010_0;
      patterns[7042] = 25'b00011011_10000000_10011011_0;
      patterns[7043] = 25'b00011011_10000001_10011100_0;
      patterns[7044] = 25'b00011011_10000010_10011101_0;
      patterns[7045] = 25'b00011011_10000011_10011110_0;
      patterns[7046] = 25'b00011011_10000100_10011111_0;
      patterns[7047] = 25'b00011011_10000101_10100000_0;
      patterns[7048] = 25'b00011011_10000110_10100001_0;
      patterns[7049] = 25'b00011011_10000111_10100010_0;
      patterns[7050] = 25'b00011011_10001000_10100011_0;
      patterns[7051] = 25'b00011011_10001001_10100100_0;
      patterns[7052] = 25'b00011011_10001010_10100101_0;
      patterns[7053] = 25'b00011011_10001011_10100110_0;
      patterns[7054] = 25'b00011011_10001100_10100111_0;
      patterns[7055] = 25'b00011011_10001101_10101000_0;
      patterns[7056] = 25'b00011011_10001110_10101001_0;
      patterns[7057] = 25'b00011011_10001111_10101010_0;
      patterns[7058] = 25'b00011011_10010000_10101011_0;
      patterns[7059] = 25'b00011011_10010001_10101100_0;
      patterns[7060] = 25'b00011011_10010010_10101101_0;
      patterns[7061] = 25'b00011011_10010011_10101110_0;
      patterns[7062] = 25'b00011011_10010100_10101111_0;
      patterns[7063] = 25'b00011011_10010101_10110000_0;
      patterns[7064] = 25'b00011011_10010110_10110001_0;
      patterns[7065] = 25'b00011011_10010111_10110010_0;
      patterns[7066] = 25'b00011011_10011000_10110011_0;
      patterns[7067] = 25'b00011011_10011001_10110100_0;
      patterns[7068] = 25'b00011011_10011010_10110101_0;
      patterns[7069] = 25'b00011011_10011011_10110110_0;
      patterns[7070] = 25'b00011011_10011100_10110111_0;
      patterns[7071] = 25'b00011011_10011101_10111000_0;
      patterns[7072] = 25'b00011011_10011110_10111001_0;
      patterns[7073] = 25'b00011011_10011111_10111010_0;
      patterns[7074] = 25'b00011011_10100000_10111011_0;
      patterns[7075] = 25'b00011011_10100001_10111100_0;
      patterns[7076] = 25'b00011011_10100010_10111101_0;
      patterns[7077] = 25'b00011011_10100011_10111110_0;
      patterns[7078] = 25'b00011011_10100100_10111111_0;
      patterns[7079] = 25'b00011011_10100101_11000000_0;
      patterns[7080] = 25'b00011011_10100110_11000001_0;
      patterns[7081] = 25'b00011011_10100111_11000010_0;
      patterns[7082] = 25'b00011011_10101000_11000011_0;
      patterns[7083] = 25'b00011011_10101001_11000100_0;
      patterns[7084] = 25'b00011011_10101010_11000101_0;
      patterns[7085] = 25'b00011011_10101011_11000110_0;
      patterns[7086] = 25'b00011011_10101100_11000111_0;
      patterns[7087] = 25'b00011011_10101101_11001000_0;
      patterns[7088] = 25'b00011011_10101110_11001001_0;
      patterns[7089] = 25'b00011011_10101111_11001010_0;
      patterns[7090] = 25'b00011011_10110000_11001011_0;
      patterns[7091] = 25'b00011011_10110001_11001100_0;
      patterns[7092] = 25'b00011011_10110010_11001101_0;
      patterns[7093] = 25'b00011011_10110011_11001110_0;
      patterns[7094] = 25'b00011011_10110100_11001111_0;
      patterns[7095] = 25'b00011011_10110101_11010000_0;
      patterns[7096] = 25'b00011011_10110110_11010001_0;
      patterns[7097] = 25'b00011011_10110111_11010010_0;
      patterns[7098] = 25'b00011011_10111000_11010011_0;
      patterns[7099] = 25'b00011011_10111001_11010100_0;
      patterns[7100] = 25'b00011011_10111010_11010101_0;
      patterns[7101] = 25'b00011011_10111011_11010110_0;
      patterns[7102] = 25'b00011011_10111100_11010111_0;
      patterns[7103] = 25'b00011011_10111101_11011000_0;
      patterns[7104] = 25'b00011011_10111110_11011001_0;
      patterns[7105] = 25'b00011011_10111111_11011010_0;
      patterns[7106] = 25'b00011011_11000000_11011011_0;
      patterns[7107] = 25'b00011011_11000001_11011100_0;
      patterns[7108] = 25'b00011011_11000010_11011101_0;
      patterns[7109] = 25'b00011011_11000011_11011110_0;
      patterns[7110] = 25'b00011011_11000100_11011111_0;
      patterns[7111] = 25'b00011011_11000101_11100000_0;
      patterns[7112] = 25'b00011011_11000110_11100001_0;
      patterns[7113] = 25'b00011011_11000111_11100010_0;
      patterns[7114] = 25'b00011011_11001000_11100011_0;
      patterns[7115] = 25'b00011011_11001001_11100100_0;
      patterns[7116] = 25'b00011011_11001010_11100101_0;
      patterns[7117] = 25'b00011011_11001011_11100110_0;
      patterns[7118] = 25'b00011011_11001100_11100111_0;
      patterns[7119] = 25'b00011011_11001101_11101000_0;
      patterns[7120] = 25'b00011011_11001110_11101001_0;
      patterns[7121] = 25'b00011011_11001111_11101010_0;
      patterns[7122] = 25'b00011011_11010000_11101011_0;
      patterns[7123] = 25'b00011011_11010001_11101100_0;
      patterns[7124] = 25'b00011011_11010010_11101101_0;
      patterns[7125] = 25'b00011011_11010011_11101110_0;
      patterns[7126] = 25'b00011011_11010100_11101111_0;
      patterns[7127] = 25'b00011011_11010101_11110000_0;
      patterns[7128] = 25'b00011011_11010110_11110001_0;
      patterns[7129] = 25'b00011011_11010111_11110010_0;
      patterns[7130] = 25'b00011011_11011000_11110011_0;
      patterns[7131] = 25'b00011011_11011001_11110100_0;
      patterns[7132] = 25'b00011011_11011010_11110101_0;
      patterns[7133] = 25'b00011011_11011011_11110110_0;
      patterns[7134] = 25'b00011011_11011100_11110111_0;
      patterns[7135] = 25'b00011011_11011101_11111000_0;
      patterns[7136] = 25'b00011011_11011110_11111001_0;
      patterns[7137] = 25'b00011011_11011111_11111010_0;
      patterns[7138] = 25'b00011011_11100000_11111011_0;
      patterns[7139] = 25'b00011011_11100001_11111100_0;
      patterns[7140] = 25'b00011011_11100010_11111101_0;
      patterns[7141] = 25'b00011011_11100011_11111110_0;
      patterns[7142] = 25'b00011011_11100100_11111111_0;
      patterns[7143] = 25'b00011011_11100101_00000000_1;
      patterns[7144] = 25'b00011011_11100110_00000001_1;
      patterns[7145] = 25'b00011011_11100111_00000010_1;
      patterns[7146] = 25'b00011011_11101000_00000011_1;
      patterns[7147] = 25'b00011011_11101001_00000100_1;
      patterns[7148] = 25'b00011011_11101010_00000101_1;
      patterns[7149] = 25'b00011011_11101011_00000110_1;
      patterns[7150] = 25'b00011011_11101100_00000111_1;
      patterns[7151] = 25'b00011011_11101101_00001000_1;
      patterns[7152] = 25'b00011011_11101110_00001001_1;
      patterns[7153] = 25'b00011011_11101111_00001010_1;
      patterns[7154] = 25'b00011011_11110000_00001011_1;
      patterns[7155] = 25'b00011011_11110001_00001100_1;
      patterns[7156] = 25'b00011011_11110010_00001101_1;
      patterns[7157] = 25'b00011011_11110011_00001110_1;
      patterns[7158] = 25'b00011011_11110100_00001111_1;
      patterns[7159] = 25'b00011011_11110101_00010000_1;
      patterns[7160] = 25'b00011011_11110110_00010001_1;
      patterns[7161] = 25'b00011011_11110111_00010010_1;
      patterns[7162] = 25'b00011011_11111000_00010011_1;
      patterns[7163] = 25'b00011011_11111001_00010100_1;
      patterns[7164] = 25'b00011011_11111010_00010101_1;
      patterns[7165] = 25'b00011011_11111011_00010110_1;
      patterns[7166] = 25'b00011011_11111100_00010111_1;
      patterns[7167] = 25'b00011011_11111101_00011000_1;
      patterns[7168] = 25'b00011011_11111110_00011001_1;
      patterns[7169] = 25'b00011011_11111111_00011010_1;
      patterns[7170] = 25'b00011100_00000000_00011100_0;
      patterns[7171] = 25'b00011100_00000001_00011101_0;
      patterns[7172] = 25'b00011100_00000010_00011110_0;
      patterns[7173] = 25'b00011100_00000011_00011111_0;
      patterns[7174] = 25'b00011100_00000100_00100000_0;
      patterns[7175] = 25'b00011100_00000101_00100001_0;
      patterns[7176] = 25'b00011100_00000110_00100010_0;
      patterns[7177] = 25'b00011100_00000111_00100011_0;
      patterns[7178] = 25'b00011100_00001000_00100100_0;
      patterns[7179] = 25'b00011100_00001001_00100101_0;
      patterns[7180] = 25'b00011100_00001010_00100110_0;
      patterns[7181] = 25'b00011100_00001011_00100111_0;
      patterns[7182] = 25'b00011100_00001100_00101000_0;
      patterns[7183] = 25'b00011100_00001101_00101001_0;
      patterns[7184] = 25'b00011100_00001110_00101010_0;
      patterns[7185] = 25'b00011100_00001111_00101011_0;
      patterns[7186] = 25'b00011100_00010000_00101100_0;
      patterns[7187] = 25'b00011100_00010001_00101101_0;
      patterns[7188] = 25'b00011100_00010010_00101110_0;
      patterns[7189] = 25'b00011100_00010011_00101111_0;
      patterns[7190] = 25'b00011100_00010100_00110000_0;
      patterns[7191] = 25'b00011100_00010101_00110001_0;
      patterns[7192] = 25'b00011100_00010110_00110010_0;
      patterns[7193] = 25'b00011100_00010111_00110011_0;
      patterns[7194] = 25'b00011100_00011000_00110100_0;
      patterns[7195] = 25'b00011100_00011001_00110101_0;
      patterns[7196] = 25'b00011100_00011010_00110110_0;
      patterns[7197] = 25'b00011100_00011011_00110111_0;
      patterns[7198] = 25'b00011100_00011100_00111000_0;
      patterns[7199] = 25'b00011100_00011101_00111001_0;
      patterns[7200] = 25'b00011100_00011110_00111010_0;
      patterns[7201] = 25'b00011100_00011111_00111011_0;
      patterns[7202] = 25'b00011100_00100000_00111100_0;
      patterns[7203] = 25'b00011100_00100001_00111101_0;
      patterns[7204] = 25'b00011100_00100010_00111110_0;
      patterns[7205] = 25'b00011100_00100011_00111111_0;
      patterns[7206] = 25'b00011100_00100100_01000000_0;
      patterns[7207] = 25'b00011100_00100101_01000001_0;
      patterns[7208] = 25'b00011100_00100110_01000010_0;
      patterns[7209] = 25'b00011100_00100111_01000011_0;
      patterns[7210] = 25'b00011100_00101000_01000100_0;
      patterns[7211] = 25'b00011100_00101001_01000101_0;
      patterns[7212] = 25'b00011100_00101010_01000110_0;
      patterns[7213] = 25'b00011100_00101011_01000111_0;
      patterns[7214] = 25'b00011100_00101100_01001000_0;
      patterns[7215] = 25'b00011100_00101101_01001001_0;
      patterns[7216] = 25'b00011100_00101110_01001010_0;
      patterns[7217] = 25'b00011100_00101111_01001011_0;
      patterns[7218] = 25'b00011100_00110000_01001100_0;
      patterns[7219] = 25'b00011100_00110001_01001101_0;
      patterns[7220] = 25'b00011100_00110010_01001110_0;
      patterns[7221] = 25'b00011100_00110011_01001111_0;
      patterns[7222] = 25'b00011100_00110100_01010000_0;
      patterns[7223] = 25'b00011100_00110101_01010001_0;
      patterns[7224] = 25'b00011100_00110110_01010010_0;
      patterns[7225] = 25'b00011100_00110111_01010011_0;
      patterns[7226] = 25'b00011100_00111000_01010100_0;
      patterns[7227] = 25'b00011100_00111001_01010101_0;
      patterns[7228] = 25'b00011100_00111010_01010110_0;
      patterns[7229] = 25'b00011100_00111011_01010111_0;
      patterns[7230] = 25'b00011100_00111100_01011000_0;
      patterns[7231] = 25'b00011100_00111101_01011001_0;
      patterns[7232] = 25'b00011100_00111110_01011010_0;
      patterns[7233] = 25'b00011100_00111111_01011011_0;
      patterns[7234] = 25'b00011100_01000000_01011100_0;
      patterns[7235] = 25'b00011100_01000001_01011101_0;
      patterns[7236] = 25'b00011100_01000010_01011110_0;
      patterns[7237] = 25'b00011100_01000011_01011111_0;
      patterns[7238] = 25'b00011100_01000100_01100000_0;
      patterns[7239] = 25'b00011100_01000101_01100001_0;
      patterns[7240] = 25'b00011100_01000110_01100010_0;
      patterns[7241] = 25'b00011100_01000111_01100011_0;
      patterns[7242] = 25'b00011100_01001000_01100100_0;
      patterns[7243] = 25'b00011100_01001001_01100101_0;
      patterns[7244] = 25'b00011100_01001010_01100110_0;
      patterns[7245] = 25'b00011100_01001011_01100111_0;
      patterns[7246] = 25'b00011100_01001100_01101000_0;
      patterns[7247] = 25'b00011100_01001101_01101001_0;
      patterns[7248] = 25'b00011100_01001110_01101010_0;
      patterns[7249] = 25'b00011100_01001111_01101011_0;
      patterns[7250] = 25'b00011100_01010000_01101100_0;
      patterns[7251] = 25'b00011100_01010001_01101101_0;
      patterns[7252] = 25'b00011100_01010010_01101110_0;
      patterns[7253] = 25'b00011100_01010011_01101111_0;
      patterns[7254] = 25'b00011100_01010100_01110000_0;
      patterns[7255] = 25'b00011100_01010101_01110001_0;
      patterns[7256] = 25'b00011100_01010110_01110010_0;
      patterns[7257] = 25'b00011100_01010111_01110011_0;
      patterns[7258] = 25'b00011100_01011000_01110100_0;
      patterns[7259] = 25'b00011100_01011001_01110101_0;
      patterns[7260] = 25'b00011100_01011010_01110110_0;
      patterns[7261] = 25'b00011100_01011011_01110111_0;
      patterns[7262] = 25'b00011100_01011100_01111000_0;
      patterns[7263] = 25'b00011100_01011101_01111001_0;
      patterns[7264] = 25'b00011100_01011110_01111010_0;
      patterns[7265] = 25'b00011100_01011111_01111011_0;
      patterns[7266] = 25'b00011100_01100000_01111100_0;
      patterns[7267] = 25'b00011100_01100001_01111101_0;
      patterns[7268] = 25'b00011100_01100010_01111110_0;
      patterns[7269] = 25'b00011100_01100011_01111111_0;
      patterns[7270] = 25'b00011100_01100100_10000000_0;
      patterns[7271] = 25'b00011100_01100101_10000001_0;
      patterns[7272] = 25'b00011100_01100110_10000010_0;
      patterns[7273] = 25'b00011100_01100111_10000011_0;
      patterns[7274] = 25'b00011100_01101000_10000100_0;
      patterns[7275] = 25'b00011100_01101001_10000101_0;
      patterns[7276] = 25'b00011100_01101010_10000110_0;
      patterns[7277] = 25'b00011100_01101011_10000111_0;
      patterns[7278] = 25'b00011100_01101100_10001000_0;
      patterns[7279] = 25'b00011100_01101101_10001001_0;
      patterns[7280] = 25'b00011100_01101110_10001010_0;
      patterns[7281] = 25'b00011100_01101111_10001011_0;
      patterns[7282] = 25'b00011100_01110000_10001100_0;
      patterns[7283] = 25'b00011100_01110001_10001101_0;
      patterns[7284] = 25'b00011100_01110010_10001110_0;
      patterns[7285] = 25'b00011100_01110011_10001111_0;
      patterns[7286] = 25'b00011100_01110100_10010000_0;
      patterns[7287] = 25'b00011100_01110101_10010001_0;
      patterns[7288] = 25'b00011100_01110110_10010010_0;
      patterns[7289] = 25'b00011100_01110111_10010011_0;
      patterns[7290] = 25'b00011100_01111000_10010100_0;
      patterns[7291] = 25'b00011100_01111001_10010101_0;
      patterns[7292] = 25'b00011100_01111010_10010110_0;
      patterns[7293] = 25'b00011100_01111011_10010111_0;
      patterns[7294] = 25'b00011100_01111100_10011000_0;
      patterns[7295] = 25'b00011100_01111101_10011001_0;
      patterns[7296] = 25'b00011100_01111110_10011010_0;
      patterns[7297] = 25'b00011100_01111111_10011011_0;
      patterns[7298] = 25'b00011100_10000000_10011100_0;
      patterns[7299] = 25'b00011100_10000001_10011101_0;
      patterns[7300] = 25'b00011100_10000010_10011110_0;
      patterns[7301] = 25'b00011100_10000011_10011111_0;
      patterns[7302] = 25'b00011100_10000100_10100000_0;
      patterns[7303] = 25'b00011100_10000101_10100001_0;
      patterns[7304] = 25'b00011100_10000110_10100010_0;
      patterns[7305] = 25'b00011100_10000111_10100011_0;
      patterns[7306] = 25'b00011100_10001000_10100100_0;
      patterns[7307] = 25'b00011100_10001001_10100101_0;
      patterns[7308] = 25'b00011100_10001010_10100110_0;
      patterns[7309] = 25'b00011100_10001011_10100111_0;
      patterns[7310] = 25'b00011100_10001100_10101000_0;
      patterns[7311] = 25'b00011100_10001101_10101001_0;
      patterns[7312] = 25'b00011100_10001110_10101010_0;
      patterns[7313] = 25'b00011100_10001111_10101011_0;
      patterns[7314] = 25'b00011100_10010000_10101100_0;
      patterns[7315] = 25'b00011100_10010001_10101101_0;
      patterns[7316] = 25'b00011100_10010010_10101110_0;
      patterns[7317] = 25'b00011100_10010011_10101111_0;
      patterns[7318] = 25'b00011100_10010100_10110000_0;
      patterns[7319] = 25'b00011100_10010101_10110001_0;
      patterns[7320] = 25'b00011100_10010110_10110010_0;
      patterns[7321] = 25'b00011100_10010111_10110011_0;
      patterns[7322] = 25'b00011100_10011000_10110100_0;
      patterns[7323] = 25'b00011100_10011001_10110101_0;
      patterns[7324] = 25'b00011100_10011010_10110110_0;
      patterns[7325] = 25'b00011100_10011011_10110111_0;
      patterns[7326] = 25'b00011100_10011100_10111000_0;
      patterns[7327] = 25'b00011100_10011101_10111001_0;
      patterns[7328] = 25'b00011100_10011110_10111010_0;
      patterns[7329] = 25'b00011100_10011111_10111011_0;
      patterns[7330] = 25'b00011100_10100000_10111100_0;
      patterns[7331] = 25'b00011100_10100001_10111101_0;
      patterns[7332] = 25'b00011100_10100010_10111110_0;
      patterns[7333] = 25'b00011100_10100011_10111111_0;
      patterns[7334] = 25'b00011100_10100100_11000000_0;
      patterns[7335] = 25'b00011100_10100101_11000001_0;
      patterns[7336] = 25'b00011100_10100110_11000010_0;
      patterns[7337] = 25'b00011100_10100111_11000011_0;
      patterns[7338] = 25'b00011100_10101000_11000100_0;
      patterns[7339] = 25'b00011100_10101001_11000101_0;
      patterns[7340] = 25'b00011100_10101010_11000110_0;
      patterns[7341] = 25'b00011100_10101011_11000111_0;
      patterns[7342] = 25'b00011100_10101100_11001000_0;
      patterns[7343] = 25'b00011100_10101101_11001001_0;
      patterns[7344] = 25'b00011100_10101110_11001010_0;
      patterns[7345] = 25'b00011100_10101111_11001011_0;
      patterns[7346] = 25'b00011100_10110000_11001100_0;
      patterns[7347] = 25'b00011100_10110001_11001101_0;
      patterns[7348] = 25'b00011100_10110010_11001110_0;
      patterns[7349] = 25'b00011100_10110011_11001111_0;
      patterns[7350] = 25'b00011100_10110100_11010000_0;
      patterns[7351] = 25'b00011100_10110101_11010001_0;
      patterns[7352] = 25'b00011100_10110110_11010010_0;
      patterns[7353] = 25'b00011100_10110111_11010011_0;
      patterns[7354] = 25'b00011100_10111000_11010100_0;
      patterns[7355] = 25'b00011100_10111001_11010101_0;
      patterns[7356] = 25'b00011100_10111010_11010110_0;
      patterns[7357] = 25'b00011100_10111011_11010111_0;
      patterns[7358] = 25'b00011100_10111100_11011000_0;
      patterns[7359] = 25'b00011100_10111101_11011001_0;
      patterns[7360] = 25'b00011100_10111110_11011010_0;
      patterns[7361] = 25'b00011100_10111111_11011011_0;
      patterns[7362] = 25'b00011100_11000000_11011100_0;
      patterns[7363] = 25'b00011100_11000001_11011101_0;
      patterns[7364] = 25'b00011100_11000010_11011110_0;
      patterns[7365] = 25'b00011100_11000011_11011111_0;
      patterns[7366] = 25'b00011100_11000100_11100000_0;
      patterns[7367] = 25'b00011100_11000101_11100001_0;
      patterns[7368] = 25'b00011100_11000110_11100010_0;
      patterns[7369] = 25'b00011100_11000111_11100011_0;
      patterns[7370] = 25'b00011100_11001000_11100100_0;
      patterns[7371] = 25'b00011100_11001001_11100101_0;
      patterns[7372] = 25'b00011100_11001010_11100110_0;
      patterns[7373] = 25'b00011100_11001011_11100111_0;
      patterns[7374] = 25'b00011100_11001100_11101000_0;
      patterns[7375] = 25'b00011100_11001101_11101001_0;
      patterns[7376] = 25'b00011100_11001110_11101010_0;
      patterns[7377] = 25'b00011100_11001111_11101011_0;
      patterns[7378] = 25'b00011100_11010000_11101100_0;
      patterns[7379] = 25'b00011100_11010001_11101101_0;
      patterns[7380] = 25'b00011100_11010010_11101110_0;
      patterns[7381] = 25'b00011100_11010011_11101111_0;
      patterns[7382] = 25'b00011100_11010100_11110000_0;
      patterns[7383] = 25'b00011100_11010101_11110001_0;
      patterns[7384] = 25'b00011100_11010110_11110010_0;
      patterns[7385] = 25'b00011100_11010111_11110011_0;
      patterns[7386] = 25'b00011100_11011000_11110100_0;
      patterns[7387] = 25'b00011100_11011001_11110101_0;
      patterns[7388] = 25'b00011100_11011010_11110110_0;
      patterns[7389] = 25'b00011100_11011011_11110111_0;
      patterns[7390] = 25'b00011100_11011100_11111000_0;
      patterns[7391] = 25'b00011100_11011101_11111001_0;
      patterns[7392] = 25'b00011100_11011110_11111010_0;
      patterns[7393] = 25'b00011100_11011111_11111011_0;
      patterns[7394] = 25'b00011100_11100000_11111100_0;
      patterns[7395] = 25'b00011100_11100001_11111101_0;
      patterns[7396] = 25'b00011100_11100010_11111110_0;
      patterns[7397] = 25'b00011100_11100011_11111111_0;
      patterns[7398] = 25'b00011100_11100100_00000000_1;
      patterns[7399] = 25'b00011100_11100101_00000001_1;
      patterns[7400] = 25'b00011100_11100110_00000010_1;
      patterns[7401] = 25'b00011100_11100111_00000011_1;
      patterns[7402] = 25'b00011100_11101000_00000100_1;
      patterns[7403] = 25'b00011100_11101001_00000101_1;
      patterns[7404] = 25'b00011100_11101010_00000110_1;
      patterns[7405] = 25'b00011100_11101011_00000111_1;
      patterns[7406] = 25'b00011100_11101100_00001000_1;
      patterns[7407] = 25'b00011100_11101101_00001001_1;
      patterns[7408] = 25'b00011100_11101110_00001010_1;
      patterns[7409] = 25'b00011100_11101111_00001011_1;
      patterns[7410] = 25'b00011100_11110000_00001100_1;
      patterns[7411] = 25'b00011100_11110001_00001101_1;
      patterns[7412] = 25'b00011100_11110010_00001110_1;
      patterns[7413] = 25'b00011100_11110011_00001111_1;
      patterns[7414] = 25'b00011100_11110100_00010000_1;
      patterns[7415] = 25'b00011100_11110101_00010001_1;
      patterns[7416] = 25'b00011100_11110110_00010010_1;
      patterns[7417] = 25'b00011100_11110111_00010011_1;
      patterns[7418] = 25'b00011100_11111000_00010100_1;
      patterns[7419] = 25'b00011100_11111001_00010101_1;
      patterns[7420] = 25'b00011100_11111010_00010110_1;
      patterns[7421] = 25'b00011100_11111011_00010111_1;
      patterns[7422] = 25'b00011100_11111100_00011000_1;
      patterns[7423] = 25'b00011100_11111101_00011001_1;
      patterns[7424] = 25'b00011100_11111110_00011010_1;
      patterns[7425] = 25'b00011100_11111111_00011011_1;
      patterns[7426] = 25'b00011101_00000000_00011101_0;
      patterns[7427] = 25'b00011101_00000001_00011110_0;
      patterns[7428] = 25'b00011101_00000010_00011111_0;
      patterns[7429] = 25'b00011101_00000011_00100000_0;
      patterns[7430] = 25'b00011101_00000100_00100001_0;
      patterns[7431] = 25'b00011101_00000101_00100010_0;
      patterns[7432] = 25'b00011101_00000110_00100011_0;
      patterns[7433] = 25'b00011101_00000111_00100100_0;
      patterns[7434] = 25'b00011101_00001000_00100101_0;
      patterns[7435] = 25'b00011101_00001001_00100110_0;
      patterns[7436] = 25'b00011101_00001010_00100111_0;
      patterns[7437] = 25'b00011101_00001011_00101000_0;
      patterns[7438] = 25'b00011101_00001100_00101001_0;
      patterns[7439] = 25'b00011101_00001101_00101010_0;
      patterns[7440] = 25'b00011101_00001110_00101011_0;
      patterns[7441] = 25'b00011101_00001111_00101100_0;
      patterns[7442] = 25'b00011101_00010000_00101101_0;
      patterns[7443] = 25'b00011101_00010001_00101110_0;
      patterns[7444] = 25'b00011101_00010010_00101111_0;
      patterns[7445] = 25'b00011101_00010011_00110000_0;
      patterns[7446] = 25'b00011101_00010100_00110001_0;
      patterns[7447] = 25'b00011101_00010101_00110010_0;
      patterns[7448] = 25'b00011101_00010110_00110011_0;
      patterns[7449] = 25'b00011101_00010111_00110100_0;
      patterns[7450] = 25'b00011101_00011000_00110101_0;
      patterns[7451] = 25'b00011101_00011001_00110110_0;
      patterns[7452] = 25'b00011101_00011010_00110111_0;
      patterns[7453] = 25'b00011101_00011011_00111000_0;
      patterns[7454] = 25'b00011101_00011100_00111001_0;
      patterns[7455] = 25'b00011101_00011101_00111010_0;
      patterns[7456] = 25'b00011101_00011110_00111011_0;
      patterns[7457] = 25'b00011101_00011111_00111100_0;
      patterns[7458] = 25'b00011101_00100000_00111101_0;
      patterns[7459] = 25'b00011101_00100001_00111110_0;
      patterns[7460] = 25'b00011101_00100010_00111111_0;
      patterns[7461] = 25'b00011101_00100011_01000000_0;
      patterns[7462] = 25'b00011101_00100100_01000001_0;
      patterns[7463] = 25'b00011101_00100101_01000010_0;
      patterns[7464] = 25'b00011101_00100110_01000011_0;
      patterns[7465] = 25'b00011101_00100111_01000100_0;
      patterns[7466] = 25'b00011101_00101000_01000101_0;
      patterns[7467] = 25'b00011101_00101001_01000110_0;
      patterns[7468] = 25'b00011101_00101010_01000111_0;
      patterns[7469] = 25'b00011101_00101011_01001000_0;
      patterns[7470] = 25'b00011101_00101100_01001001_0;
      patterns[7471] = 25'b00011101_00101101_01001010_0;
      patterns[7472] = 25'b00011101_00101110_01001011_0;
      patterns[7473] = 25'b00011101_00101111_01001100_0;
      patterns[7474] = 25'b00011101_00110000_01001101_0;
      patterns[7475] = 25'b00011101_00110001_01001110_0;
      patterns[7476] = 25'b00011101_00110010_01001111_0;
      patterns[7477] = 25'b00011101_00110011_01010000_0;
      patterns[7478] = 25'b00011101_00110100_01010001_0;
      patterns[7479] = 25'b00011101_00110101_01010010_0;
      patterns[7480] = 25'b00011101_00110110_01010011_0;
      patterns[7481] = 25'b00011101_00110111_01010100_0;
      patterns[7482] = 25'b00011101_00111000_01010101_0;
      patterns[7483] = 25'b00011101_00111001_01010110_0;
      patterns[7484] = 25'b00011101_00111010_01010111_0;
      patterns[7485] = 25'b00011101_00111011_01011000_0;
      patterns[7486] = 25'b00011101_00111100_01011001_0;
      patterns[7487] = 25'b00011101_00111101_01011010_0;
      patterns[7488] = 25'b00011101_00111110_01011011_0;
      patterns[7489] = 25'b00011101_00111111_01011100_0;
      patterns[7490] = 25'b00011101_01000000_01011101_0;
      patterns[7491] = 25'b00011101_01000001_01011110_0;
      patterns[7492] = 25'b00011101_01000010_01011111_0;
      patterns[7493] = 25'b00011101_01000011_01100000_0;
      patterns[7494] = 25'b00011101_01000100_01100001_0;
      patterns[7495] = 25'b00011101_01000101_01100010_0;
      patterns[7496] = 25'b00011101_01000110_01100011_0;
      patterns[7497] = 25'b00011101_01000111_01100100_0;
      patterns[7498] = 25'b00011101_01001000_01100101_0;
      patterns[7499] = 25'b00011101_01001001_01100110_0;
      patterns[7500] = 25'b00011101_01001010_01100111_0;
      patterns[7501] = 25'b00011101_01001011_01101000_0;
      patterns[7502] = 25'b00011101_01001100_01101001_0;
      patterns[7503] = 25'b00011101_01001101_01101010_0;
      patterns[7504] = 25'b00011101_01001110_01101011_0;
      patterns[7505] = 25'b00011101_01001111_01101100_0;
      patterns[7506] = 25'b00011101_01010000_01101101_0;
      patterns[7507] = 25'b00011101_01010001_01101110_0;
      patterns[7508] = 25'b00011101_01010010_01101111_0;
      patterns[7509] = 25'b00011101_01010011_01110000_0;
      patterns[7510] = 25'b00011101_01010100_01110001_0;
      patterns[7511] = 25'b00011101_01010101_01110010_0;
      patterns[7512] = 25'b00011101_01010110_01110011_0;
      patterns[7513] = 25'b00011101_01010111_01110100_0;
      patterns[7514] = 25'b00011101_01011000_01110101_0;
      patterns[7515] = 25'b00011101_01011001_01110110_0;
      patterns[7516] = 25'b00011101_01011010_01110111_0;
      patterns[7517] = 25'b00011101_01011011_01111000_0;
      patterns[7518] = 25'b00011101_01011100_01111001_0;
      patterns[7519] = 25'b00011101_01011101_01111010_0;
      patterns[7520] = 25'b00011101_01011110_01111011_0;
      patterns[7521] = 25'b00011101_01011111_01111100_0;
      patterns[7522] = 25'b00011101_01100000_01111101_0;
      patterns[7523] = 25'b00011101_01100001_01111110_0;
      patterns[7524] = 25'b00011101_01100010_01111111_0;
      patterns[7525] = 25'b00011101_01100011_10000000_0;
      patterns[7526] = 25'b00011101_01100100_10000001_0;
      patterns[7527] = 25'b00011101_01100101_10000010_0;
      patterns[7528] = 25'b00011101_01100110_10000011_0;
      patterns[7529] = 25'b00011101_01100111_10000100_0;
      patterns[7530] = 25'b00011101_01101000_10000101_0;
      patterns[7531] = 25'b00011101_01101001_10000110_0;
      patterns[7532] = 25'b00011101_01101010_10000111_0;
      patterns[7533] = 25'b00011101_01101011_10001000_0;
      patterns[7534] = 25'b00011101_01101100_10001001_0;
      patterns[7535] = 25'b00011101_01101101_10001010_0;
      patterns[7536] = 25'b00011101_01101110_10001011_0;
      patterns[7537] = 25'b00011101_01101111_10001100_0;
      patterns[7538] = 25'b00011101_01110000_10001101_0;
      patterns[7539] = 25'b00011101_01110001_10001110_0;
      patterns[7540] = 25'b00011101_01110010_10001111_0;
      patterns[7541] = 25'b00011101_01110011_10010000_0;
      patterns[7542] = 25'b00011101_01110100_10010001_0;
      patterns[7543] = 25'b00011101_01110101_10010010_0;
      patterns[7544] = 25'b00011101_01110110_10010011_0;
      patterns[7545] = 25'b00011101_01110111_10010100_0;
      patterns[7546] = 25'b00011101_01111000_10010101_0;
      patterns[7547] = 25'b00011101_01111001_10010110_0;
      patterns[7548] = 25'b00011101_01111010_10010111_0;
      patterns[7549] = 25'b00011101_01111011_10011000_0;
      patterns[7550] = 25'b00011101_01111100_10011001_0;
      patterns[7551] = 25'b00011101_01111101_10011010_0;
      patterns[7552] = 25'b00011101_01111110_10011011_0;
      patterns[7553] = 25'b00011101_01111111_10011100_0;
      patterns[7554] = 25'b00011101_10000000_10011101_0;
      patterns[7555] = 25'b00011101_10000001_10011110_0;
      patterns[7556] = 25'b00011101_10000010_10011111_0;
      patterns[7557] = 25'b00011101_10000011_10100000_0;
      patterns[7558] = 25'b00011101_10000100_10100001_0;
      patterns[7559] = 25'b00011101_10000101_10100010_0;
      patterns[7560] = 25'b00011101_10000110_10100011_0;
      patterns[7561] = 25'b00011101_10000111_10100100_0;
      patterns[7562] = 25'b00011101_10001000_10100101_0;
      patterns[7563] = 25'b00011101_10001001_10100110_0;
      patterns[7564] = 25'b00011101_10001010_10100111_0;
      patterns[7565] = 25'b00011101_10001011_10101000_0;
      patterns[7566] = 25'b00011101_10001100_10101001_0;
      patterns[7567] = 25'b00011101_10001101_10101010_0;
      patterns[7568] = 25'b00011101_10001110_10101011_0;
      patterns[7569] = 25'b00011101_10001111_10101100_0;
      patterns[7570] = 25'b00011101_10010000_10101101_0;
      patterns[7571] = 25'b00011101_10010001_10101110_0;
      patterns[7572] = 25'b00011101_10010010_10101111_0;
      patterns[7573] = 25'b00011101_10010011_10110000_0;
      patterns[7574] = 25'b00011101_10010100_10110001_0;
      patterns[7575] = 25'b00011101_10010101_10110010_0;
      patterns[7576] = 25'b00011101_10010110_10110011_0;
      patterns[7577] = 25'b00011101_10010111_10110100_0;
      patterns[7578] = 25'b00011101_10011000_10110101_0;
      patterns[7579] = 25'b00011101_10011001_10110110_0;
      patterns[7580] = 25'b00011101_10011010_10110111_0;
      patterns[7581] = 25'b00011101_10011011_10111000_0;
      patterns[7582] = 25'b00011101_10011100_10111001_0;
      patterns[7583] = 25'b00011101_10011101_10111010_0;
      patterns[7584] = 25'b00011101_10011110_10111011_0;
      patterns[7585] = 25'b00011101_10011111_10111100_0;
      patterns[7586] = 25'b00011101_10100000_10111101_0;
      patterns[7587] = 25'b00011101_10100001_10111110_0;
      patterns[7588] = 25'b00011101_10100010_10111111_0;
      patterns[7589] = 25'b00011101_10100011_11000000_0;
      patterns[7590] = 25'b00011101_10100100_11000001_0;
      patterns[7591] = 25'b00011101_10100101_11000010_0;
      patterns[7592] = 25'b00011101_10100110_11000011_0;
      patterns[7593] = 25'b00011101_10100111_11000100_0;
      patterns[7594] = 25'b00011101_10101000_11000101_0;
      patterns[7595] = 25'b00011101_10101001_11000110_0;
      patterns[7596] = 25'b00011101_10101010_11000111_0;
      patterns[7597] = 25'b00011101_10101011_11001000_0;
      patterns[7598] = 25'b00011101_10101100_11001001_0;
      patterns[7599] = 25'b00011101_10101101_11001010_0;
      patterns[7600] = 25'b00011101_10101110_11001011_0;
      patterns[7601] = 25'b00011101_10101111_11001100_0;
      patterns[7602] = 25'b00011101_10110000_11001101_0;
      patterns[7603] = 25'b00011101_10110001_11001110_0;
      patterns[7604] = 25'b00011101_10110010_11001111_0;
      patterns[7605] = 25'b00011101_10110011_11010000_0;
      patterns[7606] = 25'b00011101_10110100_11010001_0;
      patterns[7607] = 25'b00011101_10110101_11010010_0;
      patterns[7608] = 25'b00011101_10110110_11010011_0;
      patterns[7609] = 25'b00011101_10110111_11010100_0;
      patterns[7610] = 25'b00011101_10111000_11010101_0;
      patterns[7611] = 25'b00011101_10111001_11010110_0;
      patterns[7612] = 25'b00011101_10111010_11010111_0;
      patterns[7613] = 25'b00011101_10111011_11011000_0;
      patterns[7614] = 25'b00011101_10111100_11011001_0;
      patterns[7615] = 25'b00011101_10111101_11011010_0;
      patterns[7616] = 25'b00011101_10111110_11011011_0;
      patterns[7617] = 25'b00011101_10111111_11011100_0;
      patterns[7618] = 25'b00011101_11000000_11011101_0;
      patterns[7619] = 25'b00011101_11000001_11011110_0;
      patterns[7620] = 25'b00011101_11000010_11011111_0;
      patterns[7621] = 25'b00011101_11000011_11100000_0;
      patterns[7622] = 25'b00011101_11000100_11100001_0;
      patterns[7623] = 25'b00011101_11000101_11100010_0;
      patterns[7624] = 25'b00011101_11000110_11100011_0;
      patterns[7625] = 25'b00011101_11000111_11100100_0;
      patterns[7626] = 25'b00011101_11001000_11100101_0;
      patterns[7627] = 25'b00011101_11001001_11100110_0;
      patterns[7628] = 25'b00011101_11001010_11100111_0;
      patterns[7629] = 25'b00011101_11001011_11101000_0;
      patterns[7630] = 25'b00011101_11001100_11101001_0;
      patterns[7631] = 25'b00011101_11001101_11101010_0;
      patterns[7632] = 25'b00011101_11001110_11101011_0;
      patterns[7633] = 25'b00011101_11001111_11101100_0;
      patterns[7634] = 25'b00011101_11010000_11101101_0;
      patterns[7635] = 25'b00011101_11010001_11101110_0;
      patterns[7636] = 25'b00011101_11010010_11101111_0;
      patterns[7637] = 25'b00011101_11010011_11110000_0;
      patterns[7638] = 25'b00011101_11010100_11110001_0;
      patterns[7639] = 25'b00011101_11010101_11110010_0;
      patterns[7640] = 25'b00011101_11010110_11110011_0;
      patterns[7641] = 25'b00011101_11010111_11110100_0;
      patterns[7642] = 25'b00011101_11011000_11110101_0;
      patterns[7643] = 25'b00011101_11011001_11110110_0;
      patterns[7644] = 25'b00011101_11011010_11110111_0;
      patterns[7645] = 25'b00011101_11011011_11111000_0;
      patterns[7646] = 25'b00011101_11011100_11111001_0;
      patterns[7647] = 25'b00011101_11011101_11111010_0;
      patterns[7648] = 25'b00011101_11011110_11111011_0;
      patterns[7649] = 25'b00011101_11011111_11111100_0;
      patterns[7650] = 25'b00011101_11100000_11111101_0;
      patterns[7651] = 25'b00011101_11100001_11111110_0;
      patterns[7652] = 25'b00011101_11100010_11111111_0;
      patterns[7653] = 25'b00011101_11100011_00000000_1;
      patterns[7654] = 25'b00011101_11100100_00000001_1;
      patterns[7655] = 25'b00011101_11100101_00000010_1;
      patterns[7656] = 25'b00011101_11100110_00000011_1;
      patterns[7657] = 25'b00011101_11100111_00000100_1;
      patterns[7658] = 25'b00011101_11101000_00000101_1;
      patterns[7659] = 25'b00011101_11101001_00000110_1;
      patterns[7660] = 25'b00011101_11101010_00000111_1;
      patterns[7661] = 25'b00011101_11101011_00001000_1;
      patterns[7662] = 25'b00011101_11101100_00001001_1;
      patterns[7663] = 25'b00011101_11101101_00001010_1;
      patterns[7664] = 25'b00011101_11101110_00001011_1;
      patterns[7665] = 25'b00011101_11101111_00001100_1;
      patterns[7666] = 25'b00011101_11110000_00001101_1;
      patterns[7667] = 25'b00011101_11110001_00001110_1;
      patterns[7668] = 25'b00011101_11110010_00001111_1;
      patterns[7669] = 25'b00011101_11110011_00010000_1;
      patterns[7670] = 25'b00011101_11110100_00010001_1;
      patterns[7671] = 25'b00011101_11110101_00010010_1;
      patterns[7672] = 25'b00011101_11110110_00010011_1;
      patterns[7673] = 25'b00011101_11110111_00010100_1;
      patterns[7674] = 25'b00011101_11111000_00010101_1;
      patterns[7675] = 25'b00011101_11111001_00010110_1;
      patterns[7676] = 25'b00011101_11111010_00010111_1;
      patterns[7677] = 25'b00011101_11111011_00011000_1;
      patterns[7678] = 25'b00011101_11111100_00011001_1;
      patterns[7679] = 25'b00011101_11111101_00011010_1;
      patterns[7680] = 25'b00011101_11111110_00011011_1;
      patterns[7681] = 25'b00011101_11111111_00011100_1;
      patterns[7682] = 25'b00011110_00000000_00011110_0;
      patterns[7683] = 25'b00011110_00000001_00011111_0;
      patterns[7684] = 25'b00011110_00000010_00100000_0;
      patterns[7685] = 25'b00011110_00000011_00100001_0;
      patterns[7686] = 25'b00011110_00000100_00100010_0;
      patterns[7687] = 25'b00011110_00000101_00100011_0;
      patterns[7688] = 25'b00011110_00000110_00100100_0;
      patterns[7689] = 25'b00011110_00000111_00100101_0;
      patterns[7690] = 25'b00011110_00001000_00100110_0;
      patterns[7691] = 25'b00011110_00001001_00100111_0;
      patterns[7692] = 25'b00011110_00001010_00101000_0;
      patterns[7693] = 25'b00011110_00001011_00101001_0;
      patterns[7694] = 25'b00011110_00001100_00101010_0;
      patterns[7695] = 25'b00011110_00001101_00101011_0;
      patterns[7696] = 25'b00011110_00001110_00101100_0;
      patterns[7697] = 25'b00011110_00001111_00101101_0;
      patterns[7698] = 25'b00011110_00010000_00101110_0;
      patterns[7699] = 25'b00011110_00010001_00101111_0;
      patterns[7700] = 25'b00011110_00010010_00110000_0;
      patterns[7701] = 25'b00011110_00010011_00110001_0;
      patterns[7702] = 25'b00011110_00010100_00110010_0;
      patterns[7703] = 25'b00011110_00010101_00110011_0;
      patterns[7704] = 25'b00011110_00010110_00110100_0;
      patterns[7705] = 25'b00011110_00010111_00110101_0;
      patterns[7706] = 25'b00011110_00011000_00110110_0;
      patterns[7707] = 25'b00011110_00011001_00110111_0;
      patterns[7708] = 25'b00011110_00011010_00111000_0;
      patterns[7709] = 25'b00011110_00011011_00111001_0;
      patterns[7710] = 25'b00011110_00011100_00111010_0;
      patterns[7711] = 25'b00011110_00011101_00111011_0;
      patterns[7712] = 25'b00011110_00011110_00111100_0;
      patterns[7713] = 25'b00011110_00011111_00111101_0;
      patterns[7714] = 25'b00011110_00100000_00111110_0;
      patterns[7715] = 25'b00011110_00100001_00111111_0;
      patterns[7716] = 25'b00011110_00100010_01000000_0;
      patterns[7717] = 25'b00011110_00100011_01000001_0;
      patterns[7718] = 25'b00011110_00100100_01000010_0;
      patterns[7719] = 25'b00011110_00100101_01000011_0;
      patterns[7720] = 25'b00011110_00100110_01000100_0;
      patterns[7721] = 25'b00011110_00100111_01000101_0;
      patterns[7722] = 25'b00011110_00101000_01000110_0;
      patterns[7723] = 25'b00011110_00101001_01000111_0;
      patterns[7724] = 25'b00011110_00101010_01001000_0;
      patterns[7725] = 25'b00011110_00101011_01001001_0;
      patterns[7726] = 25'b00011110_00101100_01001010_0;
      patterns[7727] = 25'b00011110_00101101_01001011_0;
      patterns[7728] = 25'b00011110_00101110_01001100_0;
      patterns[7729] = 25'b00011110_00101111_01001101_0;
      patterns[7730] = 25'b00011110_00110000_01001110_0;
      patterns[7731] = 25'b00011110_00110001_01001111_0;
      patterns[7732] = 25'b00011110_00110010_01010000_0;
      patterns[7733] = 25'b00011110_00110011_01010001_0;
      patterns[7734] = 25'b00011110_00110100_01010010_0;
      patterns[7735] = 25'b00011110_00110101_01010011_0;
      patterns[7736] = 25'b00011110_00110110_01010100_0;
      patterns[7737] = 25'b00011110_00110111_01010101_0;
      patterns[7738] = 25'b00011110_00111000_01010110_0;
      patterns[7739] = 25'b00011110_00111001_01010111_0;
      patterns[7740] = 25'b00011110_00111010_01011000_0;
      patterns[7741] = 25'b00011110_00111011_01011001_0;
      patterns[7742] = 25'b00011110_00111100_01011010_0;
      patterns[7743] = 25'b00011110_00111101_01011011_0;
      patterns[7744] = 25'b00011110_00111110_01011100_0;
      patterns[7745] = 25'b00011110_00111111_01011101_0;
      patterns[7746] = 25'b00011110_01000000_01011110_0;
      patterns[7747] = 25'b00011110_01000001_01011111_0;
      patterns[7748] = 25'b00011110_01000010_01100000_0;
      patterns[7749] = 25'b00011110_01000011_01100001_0;
      patterns[7750] = 25'b00011110_01000100_01100010_0;
      patterns[7751] = 25'b00011110_01000101_01100011_0;
      patterns[7752] = 25'b00011110_01000110_01100100_0;
      patterns[7753] = 25'b00011110_01000111_01100101_0;
      patterns[7754] = 25'b00011110_01001000_01100110_0;
      patterns[7755] = 25'b00011110_01001001_01100111_0;
      patterns[7756] = 25'b00011110_01001010_01101000_0;
      patterns[7757] = 25'b00011110_01001011_01101001_0;
      patterns[7758] = 25'b00011110_01001100_01101010_0;
      patterns[7759] = 25'b00011110_01001101_01101011_0;
      patterns[7760] = 25'b00011110_01001110_01101100_0;
      patterns[7761] = 25'b00011110_01001111_01101101_0;
      patterns[7762] = 25'b00011110_01010000_01101110_0;
      patterns[7763] = 25'b00011110_01010001_01101111_0;
      patterns[7764] = 25'b00011110_01010010_01110000_0;
      patterns[7765] = 25'b00011110_01010011_01110001_0;
      patterns[7766] = 25'b00011110_01010100_01110010_0;
      patterns[7767] = 25'b00011110_01010101_01110011_0;
      patterns[7768] = 25'b00011110_01010110_01110100_0;
      patterns[7769] = 25'b00011110_01010111_01110101_0;
      patterns[7770] = 25'b00011110_01011000_01110110_0;
      patterns[7771] = 25'b00011110_01011001_01110111_0;
      patterns[7772] = 25'b00011110_01011010_01111000_0;
      patterns[7773] = 25'b00011110_01011011_01111001_0;
      patterns[7774] = 25'b00011110_01011100_01111010_0;
      patterns[7775] = 25'b00011110_01011101_01111011_0;
      patterns[7776] = 25'b00011110_01011110_01111100_0;
      patterns[7777] = 25'b00011110_01011111_01111101_0;
      patterns[7778] = 25'b00011110_01100000_01111110_0;
      patterns[7779] = 25'b00011110_01100001_01111111_0;
      patterns[7780] = 25'b00011110_01100010_10000000_0;
      patterns[7781] = 25'b00011110_01100011_10000001_0;
      patterns[7782] = 25'b00011110_01100100_10000010_0;
      patterns[7783] = 25'b00011110_01100101_10000011_0;
      patterns[7784] = 25'b00011110_01100110_10000100_0;
      patterns[7785] = 25'b00011110_01100111_10000101_0;
      patterns[7786] = 25'b00011110_01101000_10000110_0;
      patterns[7787] = 25'b00011110_01101001_10000111_0;
      patterns[7788] = 25'b00011110_01101010_10001000_0;
      patterns[7789] = 25'b00011110_01101011_10001001_0;
      patterns[7790] = 25'b00011110_01101100_10001010_0;
      patterns[7791] = 25'b00011110_01101101_10001011_0;
      patterns[7792] = 25'b00011110_01101110_10001100_0;
      patterns[7793] = 25'b00011110_01101111_10001101_0;
      patterns[7794] = 25'b00011110_01110000_10001110_0;
      patterns[7795] = 25'b00011110_01110001_10001111_0;
      patterns[7796] = 25'b00011110_01110010_10010000_0;
      patterns[7797] = 25'b00011110_01110011_10010001_0;
      patterns[7798] = 25'b00011110_01110100_10010010_0;
      patterns[7799] = 25'b00011110_01110101_10010011_0;
      patterns[7800] = 25'b00011110_01110110_10010100_0;
      patterns[7801] = 25'b00011110_01110111_10010101_0;
      patterns[7802] = 25'b00011110_01111000_10010110_0;
      patterns[7803] = 25'b00011110_01111001_10010111_0;
      patterns[7804] = 25'b00011110_01111010_10011000_0;
      patterns[7805] = 25'b00011110_01111011_10011001_0;
      patterns[7806] = 25'b00011110_01111100_10011010_0;
      patterns[7807] = 25'b00011110_01111101_10011011_0;
      patterns[7808] = 25'b00011110_01111110_10011100_0;
      patterns[7809] = 25'b00011110_01111111_10011101_0;
      patterns[7810] = 25'b00011110_10000000_10011110_0;
      patterns[7811] = 25'b00011110_10000001_10011111_0;
      patterns[7812] = 25'b00011110_10000010_10100000_0;
      patterns[7813] = 25'b00011110_10000011_10100001_0;
      patterns[7814] = 25'b00011110_10000100_10100010_0;
      patterns[7815] = 25'b00011110_10000101_10100011_0;
      patterns[7816] = 25'b00011110_10000110_10100100_0;
      patterns[7817] = 25'b00011110_10000111_10100101_0;
      patterns[7818] = 25'b00011110_10001000_10100110_0;
      patterns[7819] = 25'b00011110_10001001_10100111_0;
      patterns[7820] = 25'b00011110_10001010_10101000_0;
      patterns[7821] = 25'b00011110_10001011_10101001_0;
      patterns[7822] = 25'b00011110_10001100_10101010_0;
      patterns[7823] = 25'b00011110_10001101_10101011_0;
      patterns[7824] = 25'b00011110_10001110_10101100_0;
      patterns[7825] = 25'b00011110_10001111_10101101_0;
      patterns[7826] = 25'b00011110_10010000_10101110_0;
      patterns[7827] = 25'b00011110_10010001_10101111_0;
      patterns[7828] = 25'b00011110_10010010_10110000_0;
      patterns[7829] = 25'b00011110_10010011_10110001_0;
      patterns[7830] = 25'b00011110_10010100_10110010_0;
      patterns[7831] = 25'b00011110_10010101_10110011_0;
      patterns[7832] = 25'b00011110_10010110_10110100_0;
      patterns[7833] = 25'b00011110_10010111_10110101_0;
      patterns[7834] = 25'b00011110_10011000_10110110_0;
      patterns[7835] = 25'b00011110_10011001_10110111_0;
      patterns[7836] = 25'b00011110_10011010_10111000_0;
      patterns[7837] = 25'b00011110_10011011_10111001_0;
      patterns[7838] = 25'b00011110_10011100_10111010_0;
      patterns[7839] = 25'b00011110_10011101_10111011_0;
      patterns[7840] = 25'b00011110_10011110_10111100_0;
      patterns[7841] = 25'b00011110_10011111_10111101_0;
      patterns[7842] = 25'b00011110_10100000_10111110_0;
      patterns[7843] = 25'b00011110_10100001_10111111_0;
      patterns[7844] = 25'b00011110_10100010_11000000_0;
      patterns[7845] = 25'b00011110_10100011_11000001_0;
      patterns[7846] = 25'b00011110_10100100_11000010_0;
      patterns[7847] = 25'b00011110_10100101_11000011_0;
      patterns[7848] = 25'b00011110_10100110_11000100_0;
      patterns[7849] = 25'b00011110_10100111_11000101_0;
      patterns[7850] = 25'b00011110_10101000_11000110_0;
      patterns[7851] = 25'b00011110_10101001_11000111_0;
      patterns[7852] = 25'b00011110_10101010_11001000_0;
      patterns[7853] = 25'b00011110_10101011_11001001_0;
      patterns[7854] = 25'b00011110_10101100_11001010_0;
      patterns[7855] = 25'b00011110_10101101_11001011_0;
      patterns[7856] = 25'b00011110_10101110_11001100_0;
      patterns[7857] = 25'b00011110_10101111_11001101_0;
      patterns[7858] = 25'b00011110_10110000_11001110_0;
      patterns[7859] = 25'b00011110_10110001_11001111_0;
      patterns[7860] = 25'b00011110_10110010_11010000_0;
      patterns[7861] = 25'b00011110_10110011_11010001_0;
      patterns[7862] = 25'b00011110_10110100_11010010_0;
      patterns[7863] = 25'b00011110_10110101_11010011_0;
      patterns[7864] = 25'b00011110_10110110_11010100_0;
      patterns[7865] = 25'b00011110_10110111_11010101_0;
      patterns[7866] = 25'b00011110_10111000_11010110_0;
      patterns[7867] = 25'b00011110_10111001_11010111_0;
      patterns[7868] = 25'b00011110_10111010_11011000_0;
      patterns[7869] = 25'b00011110_10111011_11011001_0;
      patterns[7870] = 25'b00011110_10111100_11011010_0;
      patterns[7871] = 25'b00011110_10111101_11011011_0;
      patterns[7872] = 25'b00011110_10111110_11011100_0;
      patterns[7873] = 25'b00011110_10111111_11011101_0;
      patterns[7874] = 25'b00011110_11000000_11011110_0;
      patterns[7875] = 25'b00011110_11000001_11011111_0;
      patterns[7876] = 25'b00011110_11000010_11100000_0;
      patterns[7877] = 25'b00011110_11000011_11100001_0;
      patterns[7878] = 25'b00011110_11000100_11100010_0;
      patterns[7879] = 25'b00011110_11000101_11100011_0;
      patterns[7880] = 25'b00011110_11000110_11100100_0;
      patterns[7881] = 25'b00011110_11000111_11100101_0;
      patterns[7882] = 25'b00011110_11001000_11100110_0;
      patterns[7883] = 25'b00011110_11001001_11100111_0;
      patterns[7884] = 25'b00011110_11001010_11101000_0;
      patterns[7885] = 25'b00011110_11001011_11101001_0;
      patterns[7886] = 25'b00011110_11001100_11101010_0;
      patterns[7887] = 25'b00011110_11001101_11101011_0;
      patterns[7888] = 25'b00011110_11001110_11101100_0;
      patterns[7889] = 25'b00011110_11001111_11101101_0;
      patterns[7890] = 25'b00011110_11010000_11101110_0;
      patterns[7891] = 25'b00011110_11010001_11101111_0;
      patterns[7892] = 25'b00011110_11010010_11110000_0;
      patterns[7893] = 25'b00011110_11010011_11110001_0;
      patterns[7894] = 25'b00011110_11010100_11110010_0;
      patterns[7895] = 25'b00011110_11010101_11110011_0;
      patterns[7896] = 25'b00011110_11010110_11110100_0;
      patterns[7897] = 25'b00011110_11010111_11110101_0;
      patterns[7898] = 25'b00011110_11011000_11110110_0;
      patterns[7899] = 25'b00011110_11011001_11110111_0;
      patterns[7900] = 25'b00011110_11011010_11111000_0;
      patterns[7901] = 25'b00011110_11011011_11111001_0;
      patterns[7902] = 25'b00011110_11011100_11111010_0;
      patterns[7903] = 25'b00011110_11011101_11111011_0;
      patterns[7904] = 25'b00011110_11011110_11111100_0;
      patterns[7905] = 25'b00011110_11011111_11111101_0;
      patterns[7906] = 25'b00011110_11100000_11111110_0;
      patterns[7907] = 25'b00011110_11100001_11111111_0;
      patterns[7908] = 25'b00011110_11100010_00000000_1;
      patterns[7909] = 25'b00011110_11100011_00000001_1;
      patterns[7910] = 25'b00011110_11100100_00000010_1;
      patterns[7911] = 25'b00011110_11100101_00000011_1;
      patterns[7912] = 25'b00011110_11100110_00000100_1;
      patterns[7913] = 25'b00011110_11100111_00000101_1;
      patterns[7914] = 25'b00011110_11101000_00000110_1;
      patterns[7915] = 25'b00011110_11101001_00000111_1;
      patterns[7916] = 25'b00011110_11101010_00001000_1;
      patterns[7917] = 25'b00011110_11101011_00001001_1;
      patterns[7918] = 25'b00011110_11101100_00001010_1;
      patterns[7919] = 25'b00011110_11101101_00001011_1;
      patterns[7920] = 25'b00011110_11101110_00001100_1;
      patterns[7921] = 25'b00011110_11101111_00001101_1;
      patterns[7922] = 25'b00011110_11110000_00001110_1;
      patterns[7923] = 25'b00011110_11110001_00001111_1;
      patterns[7924] = 25'b00011110_11110010_00010000_1;
      patterns[7925] = 25'b00011110_11110011_00010001_1;
      patterns[7926] = 25'b00011110_11110100_00010010_1;
      patterns[7927] = 25'b00011110_11110101_00010011_1;
      patterns[7928] = 25'b00011110_11110110_00010100_1;
      patterns[7929] = 25'b00011110_11110111_00010101_1;
      patterns[7930] = 25'b00011110_11111000_00010110_1;
      patterns[7931] = 25'b00011110_11111001_00010111_1;
      patterns[7932] = 25'b00011110_11111010_00011000_1;
      patterns[7933] = 25'b00011110_11111011_00011001_1;
      patterns[7934] = 25'b00011110_11111100_00011010_1;
      patterns[7935] = 25'b00011110_11111101_00011011_1;
      patterns[7936] = 25'b00011110_11111110_00011100_1;
      patterns[7937] = 25'b00011110_11111111_00011101_1;
      patterns[7938] = 25'b00011111_00000000_00011111_0;
      patterns[7939] = 25'b00011111_00000001_00100000_0;
      patterns[7940] = 25'b00011111_00000010_00100001_0;
      patterns[7941] = 25'b00011111_00000011_00100010_0;
      patterns[7942] = 25'b00011111_00000100_00100011_0;
      patterns[7943] = 25'b00011111_00000101_00100100_0;
      patterns[7944] = 25'b00011111_00000110_00100101_0;
      patterns[7945] = 25'b00011111_00000111_00100110_0;
      patterns[7946] = 25'b00011111_00001000_00100111_0;
      patterns[7947] = 25'b00011111_00001001_00101000_0;
      patterns[7948] = 25'b00011111_00001010_00101001_0;
      patterns[7949] = 25'b00011111_00001011_00101010_0;
      patterns[7950] = 25'b00011111_00001100_00101011_0;
      patterns[7951] = 25'b00011111_00001101_00101100_0;
      patterns[7952] = 25'b00011111_00001110_00101101_0;
      patterns[7953] = 25'b00011111_00001111_00101110_0;
      patterns[7954] = 25'b00011111_00010000_00101111_0;
      patterns[7955] = 25'b00011111_00010001_00110000_0;
      patterns[7956] = 25'b00011111_00010010_00110001_0;
      patterns[7957] = 25'b00011111_00010011_00110010_0;
      patterns[7958] = 25'b00011111_00010100_00110011_0;
      patterns[7959] = 25'b00011111_00010101_00110100_0;
      patterns[7960] = 25'b00011111_00010110_00110101_0;
      patterns[7961] = 25'b00011111_00010111_00110110_0;
      patterns[7962] = 25'b00011111_00011000_00110111_0;
      patterns[7963] = 25'b00011111_00011001_00111000_0;
      patterns[7964] = 25'b00011111_00011010_00111001_0;
      patterns[7965] = 25'b00011111_00011011_00111010_0;
      patterns[7966] = 25'b00011111_00011100_00111011_0;
      patterns[7967] = 25'b00011111_00011101_00111100_0;
      patterns[7968] = 25'b00011111_00011110_00111101_0;
      patterns[7969] = 25'b00011111_00011111_00111110_0;
      patterns[7970] = 25'b00011111_00100000_00111111_0;
      patterns[7971] = 25'b00011111_00100001_01000000_0;
      patterns[7972] = 25'b00011111_00100010_01000001_0;
      patterns[7973] = 25'b00011111_00100011_01000010_0;
      patterns[7974] = 25'b00011111_00100100_01000011_0;
      patterns[7975] = 25'b00011111_00100101_01000100_0;
      patterns[7976] = 25'b00011111_00100110_01000101_0;
      patterns[7977] = 25'b00011111_00100111_01000110_0;
      patterns[7978] = 25'b00011111_00101000_01000111_0;
      patterns[7979] = 25'b00011111_00101001_01001000_0;
      patterns[7980] = 25'b00011111_00101010_01001001_0;
      patterns[7981] = 25'b00011111_00101011_01001010_0;
      patterns[7982] = 25'b00011111_00101100_01001011_0;
      patterns[7983] = 25'b00011111_00101101_01001100_0;
      patterns[7984] = 25'b00011111_00101110_01001101_0;
      patterns[7985] = 25'b00011111_00101111_01001110_0;
      patterns[7986] = 25'b00011111_00110000_01001111_0;
      patterns[7987] = 25'b00011111_00110001_01010000_0;
      patterns[7988] = 25'b00011111_00110010_01010001_0;
      patterns[7989] = 25'b00011111_00110011_01010010_0;
      patterns[7990] = 25'b00011111_00110100_01010011_0;
      patterns[7991] = 25'b00011111_00110101_01010100_0;
      patterns[7992] = 25'b00011111_00110110_01010101_0;
      patterns[7993] = 25'b00011111_00110111_01010110_0;
      patterns[7994] = 25'b00011111_00111000_01010111_0;
      patterns[7995] = 25'b00011111_00111001_01011000_0;
      patterns[7996] = 25'b00011111_00111010_01011001_0;
      patterns[7997] = 25'b00011111_00111011_01011010_0;
      patterns[7998] = 25'b00011111_00111100_01011011_0;
      patterns[7999] = 25'b00011111_00111101_01011100_0;
      patterns[8000] = 25'b00011111_00111110_01011101_0;
      patterns[8001] = 25'b00011111_00111111_01011110_0;
      patterns[8002] = 25'b00011111_01000000_01011111_0;
      patterns[8003] = 25'b00011111_01000001_01100000_0;
      patterns[8004] = 25'b00011111_01000010_01100001_0;
      patterns[8005] = 25'b00011111_01000011_01100010_0;
      patterns[8006] = 25'b00011111_01000100_01100011_0;
      patterns[8007] = 25'b00011111_01000101_01100100_0;
      patterns[8008] = 25'b00011111_01000110_01100101_0;
      patterns[8009] = 25'b00011111_01000111_01100110_0;
      patterns[8010] = 25'b00011111_01001000_01100111_0;
      patterns[8011] = 25'b00011111_01001001_01101000_0;
      patterns[8012] = 25'b00011111_01001010_01101001_0;
      patterns[8013] = 25'b00011111_01001011_01101010_0;
      patterns[8014] = 25'b00011111_01001100_01101011_0;
      patterns[8015] = 25'b00011111_01001101_01101100_0;
      patterns[8016] = 25'b00011111_01001110_01101101_0;
      patterns[8017] = 25'b00011111_01001111_01101110_0;
      patterns[8018] = 25'b00011111_01010000_01101111_0;
      patterns[8019] = 25'b00011111_01010001_01110000_0;
      patterns[8020] = 25'b00011111_01010010_01110001_0;
      patterns[8021] = 25'b00011111_01010011_01110010_0;
      patterns[8022] = 25'b00011111_01010100_01110011_0;
      patterns[8023] = 25'b00011111_01010101_01110100_0;
      patterns[8024] = 25'b00011111_01010110_01110101_0;
      patterns[8025] = 25'b00011111_01010111_01110110_0;
      patterns[8026] = 25'b00011111_01011000_01110111_0;
      patterns[8027] = 25'b00011111_01011001_01111000_0;
      patterns[8028] = 25'b00011111_01011010_01111001_0;
      patterns[8029] = 25'b00011111_01011011_01111010_0;
      patterns[8030] = 25'b00011111_01011100_01111011_0;
      patterns[8031] = 25'b00011111_01011101_01111100_0;
      patterns[8032] = 25'b00011111_01011110_01111101_0;
      patterns[8033] = 25'b00011111_01011111_01111110_0;
      patterns[8034] = 25'b00011111_01100000_01111111_0;
      patterns[8035] = 25'b00011111_01100001_10000000_0;
      patterns[8036] = 25'b00011111_01100010_10000001_0;
      patterns[8037] = 25'b00011111_01100011_10000010_0;
      patterns[8038] = 25'b00011111_01100100_10000011_0;
      patterns[8039] = 25'b00011111_01100101_10000100_0;
      patterns[8040] = 25'b00011111_01100110_10000101_0;
      patterns[8041] = 25'b00011111_01100111_10000110_0;
      patterns[8042] = 25'b00011111_01101000_10000111_0;
      patterns[8043] = 25'b00011111_01101001_10001000_0;
      patterns[8044] = 25'b00011111_01101010_10001001_0;
      patterns[8045] = 25'b00011111_01101011_10001010_0;
      patterns[8046] = 25'b00011111_01101100_10001011_0;
      patterns[8047] = 25'b00011111_01101101_10001100_0;
      patterns[8048] = 25'b00011111_01101110_10001101_0;
      patterns[8049] = 25'b00011111_01101111_10001110_0;
      patterns[8050] = 25'b00011111_01110000_10001111_0;
      patterns[8051] = 25'b00011111_01110001_10010000_0;
      patterns[8052] = 25'b00011111_01110010_10010001_0;
      patterns[8053] = 25'b00011111_01110011_10010010_0;
      patterns[8054] = 25'b00011111_01110100_10010011_0;
      patterns[8055] = 25'b00011111_01110101_10010100_0;
      patterns[8056] = 25'b00011111_01110110_10010101_0;
      patterns[8057] = 25'b00011111_01110111_10010110_0;
      patterns[8058] = 25'b00011111_01111000_10010111_0;
      patterns[8059] = 25'b00011111_01111001_10011000_0;
      patterns[8060] = 25'b00011111_01111010_10011001_0;
      patterns[8061] = 25'b00011111_01111011_10011010_0;
      patterns[8062] = 25'b00011111_01111100_10011011_0;
      patterns[8063] = 25'b00011111_01111101_10011100_0;
      patterns[8064] = 25'b00011111_01111110_10011101_0;
      patterns[8065] = 25'b00011111_01111111_10011110_0;
      patterns[8066] = 25'b00011111_10000000_10011111_0;
      patterns[8067] = 25'b00011111_10000001_10100000_0;
      patterns[8068] = 25'b00011111_10000010_10100001_0;
      patterns[8069] = 25'b00011111_10000011_10100010_0;
      patterns[8070] = 25'b00011111_10000100_10100011_0;
      patterns[8071] = 25'b00011111_10000101_10100100_0;
      patterns[8072] = 25'b00011111_10000110_10100101_0;
      patterns[8073] = 25'b00011111_10000111_10100110_0;
      patterns[8074] = 25'b00011111_10001000_10100111_0;
      patterns[8075] = 25'b00011111_10001001_10101000_0;
      patterns[8076] = 25'b00011111_10001010_10101001_0;
      patterns[8077] = 25'b00011111_10001011_10101010_0;
      patterns[8078] = 25'b00011111_10001100_10101011_0;
      patterns[8079] = 25'b00011111_10001101_10101100_0;
      patterns[8080] = 25'b00011111_10001110_10101101_0;
      patterns[8081] = 25'b00011111_10001111_10101110_0;
      patterns[8082] = 25'b00011111_10010000_10101111_0;
      patterns[8083] = 25'b00011111_10010001_10110000_0;
      patterns[8084] = 25'b00011111_10010010_10110001_0;
      patterns[8085] = 25'b00011111_10010011_10110010_0;
      patterns[8086] = 25'b00011111_10010100_10110011_0;
      patterns[8087] = 25'b00011111_10010101_10110100_0;
      patterns[8088] = 25'b00011111_10010110_10110101_0;
      patterns[8089] = 25'b00011111_10010111_10110110_0;
      patterns[8090] = 25'b00011111_10011000_10110111_0;
      patterns[8091] = 25'b00011111_10011001_10111000_0;
      patterns[8092] = 25'b00011111_10011010_10111001_0;
      patterns[8093] = 25'b00011111_10011011_10111010_0;
      patterns[8094] = 25'b00011111_10011100_10111011_0;
      patterns[8095] = 25'b00011111_10011101_10111100_0;
      patterns[8096] = 25'b00011111_10011110_10111101_0;
      patterns[8097] = 25'b00011111_10011111_10111110_0;
      patterns[8098] = 25'b00011111_10100000_10111111_0;
      patterns[8099] = 25'b00011111_10100001_11000000_0;
      patterns[8100] = 25'b00011111_10100010_11000001_0;
      patterns[8101] = 25'b00011111_10100011_11000010_0;
      patterns[8102] = 25'b00011111_10100100_11000011_0;
      patterns[8103] = 25'b00011111_10100101_11000100_0;
      patterns[8104] = 25'b00011111_10100110_11000101_0;
      patterns[8105] = 25'b00011111_10100111_11000110_0;
      patterns[8106] = 25'b00011111_10101000_11000111_0;
      patterns[8107] = 25'b00011111_10101001_11001000_0;
      patterns[8108] = 25'b00011111_10101010_11001001_0;
      patterns[8109] = 25'b00011111_10101011_11001010_0;
      patterns[8110] = 25'b00011111_10101100_11001011_0;
      patterns[8111] = 25'b00011111_10101101_11001100_0;
      patterns[8112] = 25'b00011111_10101110_11001101_0;
      patterns[8113] = 25'b00011111_10101111_11001110_0;
      patterns[8114] = 25'b00011111_10110000_11001111_0;
      patterns[8115] = 25'b00011111_10110001_11010000_0;
      patterns[8116] = 25'b00011111_10110010_11010001_0;
      patterns[8117] = 25'b00011111_10110011_11010010_0;
      patterns[8118] = 25'b00011111_10110100_11010011_0;
      patterns[8119] = 25'b00011111_10110101_11010100_0;
      patterns[8120] = 25'b00011111_10110110_11010101_0;
      patterns[8121] = 25'b00011111_10110111_11010110_0;
      patterns[8122] = 25'b00011111_10111000_11010111_0;
      patterns[8123] = 25'b00011111_10111001_11011000_0;
      patterns[8124] = 25'b00011111_10111010_11011001_0;
      patterns[8125] = 25'b00011111_10111011_11011010_0;
      patterns[8126] = 25'b00011111_10111100_11011011_0;
      patterns[8127] = 25'b00011111_10111101_11011100_0;
      patterns[8128] = 25'b00011111_10111110_11011101_0;
      patterns[8129] = 25'b00011111_10111111_11011110_0;
      patterns[8130] = 25'b00011111_11000000_11011111_0;
      patterns[8131] = 25'b00011111_11000001_11100000_0;
      patterns[8132] = 25'b00011111_11000010_11100001_0;
      patterns[8133] = 25'b00011111_11000011_11100010_0;
      patterns[8134] = 25'b00011111_11000100_11100011_0;
      patterns[8135] = 25'b00011111_11000101_11100100_0;
      patterns[8136] = 25'b00011111_11000110_11100101_0;
      patterns[8137] = 25'b00011111_11000111_11100110_0;
      patterns[8138] = 25'b00011111_11001000_11100111_0;
      patterns[8139] = 25'b00011111_11001001_11101000_0;
      patterns[8140] = 25'b00011111_11001010_11101001_0;
      patterns[8141] = 25'b00011111_11001011_11101010_0;
      patterns[8142] = 25'b00011111_11001100_11101011_0;
      patterns[8143] = 25'b00011111_11001101_11101100_0;
      patterns[8144] = 25'b00011111_11001110_11101101_0;
      patterns[8145] = 25'b00011111_11001111_11101110_0;
      patterns[8146] = 25'b00011111_11010000_11101111_0;
      patterns[8147] = 25'b00011111_11010001_11110000_0;
      patterns[8148] = 25'b00011111_11010010_11110001_0;
      patterns[8149] = 25'b00011111_11010011_11110010_0;
      patterns[8150] = 25'b00011111_11010100_11110011_0;
      patterns[8151] = 25'b00011111_11010101_11110100_0;
      patterns[8152] = 25'b00011111_11010110_11110101_0;
      patterns[8153] = 25'b00011111_11010111_11110110_0;
      patterns[8154] = 25'b00011111_11011000_11110111_0;
      patterns[8155] = 25'b00011111_11011001_11111000_0;
      patterns[8156] = 25'b00011111_11011010_11111001_0;
      patterns[8157] = 25'b00011111_11011011_11111010_0;
      patterns[8158] = 25'b00011111_11011100_11111011_0;
      patterns[8159] = 25'b00011111_11011101_11111100_0;
      patterns[8160] = 25'b00011111_11011110_11111101_0;
      patterns[8161] = 25'b00011111_11011111_11111110_0;
      patterns[8162] = 25'b00011111_11100000_11111111_0;
      patterns[8163] = 25'b00011111_11100001_00000000_1;
      patterns[8164] = 25'b00011111_11100010_00000001_1;
      patterns[8165] = 25'b00011111_11100011_00000010_1;
      patterns[8166] = 25'b00011111_11100100_00000011_1;
      patterns[8167] = 25'b00011111_11100101_00000100_1;
      patterns[8168] = 25'b00011111_11100110_00000101_1;
      patterns[8169] = 25'b00011111_11100111_00000110_1;
      patterns[8170] = 25'b00011111_11101000_00000111_1;
      patterns[8171] = 25'b00011111_11101001_00001000_1;
      patterns[8172] = 25'b00011111_11101010_00001001_1;
      patterns[8173] = 25'b00011111_11101011_00001010_1;
      patterns[8174] = 25'b00011111_11101100_00001011_1;
      patterns[8175] = 25'b00011111_11101101_00001100_1;
      patterns[8176] = 25'b00011111_11101110_00001101_1;
      patterns[8177] = 25'b00011111_11101111_00001110_1;
      patterns[8178] = 25'b00011111_11110000_00001111_1;
      patterns[8179] = 25'b00011111_11110001_00010000_1;
      patterns[8180] = 25'b00011111_11110010_00010001_1;
      patterns[8181] = 25'b00011111_11110011_00010010_1;
      patterns[8182] = 25'b00011111_11110100_00010011_1;
      patterns[8183] = 25'b00011111_11110101_00010100_1;
      patterns[8184] = 25'b00011111_11110110_00010101_1;
      patterns[8185] = 25'b00011111_11110111_00010110_1;
      patterns[8186] = 25'b00011111_11111000_00010111_1;
      patterns[8187] = 25'b00011111_11111001_00011000_1;
      patterns[8188] = 25'b00011111_11111010_00011001_1;
      patterns[8189] = 25'b00011111_11111011_00011010_1;
      patterns[8190] = 25'b00011111_11111100_00011011_1;
      patterns[8191] = 25'b00011111_11111101_00011100_1;
      patterns[8192] = 25'b00011111_11111110_00011101_1;
      patterns[8193] = 25'b00011111_11111111_00011110_1;
      patterns[8194] = 25'b00100000_00000000_00100000_0;
      patterns[8195] = 25'b00100000_00000001_00100001_0;
      patterns[8196] = 25'b00100000_00000010_00100010_0;
      patterns[8197] = 25'b00100000_00000011_00100011_0;
      patterns[8198] = 25'b00100000_00000100_00100100_0;
      patterns[8199] = 25'b00100000_00000101_00100101_0;
      patterns[8200] = 25'b00100000_00000110_00100110_0;
      patterns[8201] = 25'b00100000_00000111_00100111_0;
      patterns[8202] = 25'b00100000_00001000_00101000_0;
      patterns[8203] = 25'b00100000_00001001_00101001_0;
      patterns[8204] = 25'b00100000_00001010_00101010_0;
      patterns[8205] = 25'b00100000_00001011_00101011_0;
      patterns[8206] = 25'b00100000_00001100_00101100_0;
      patterns[8207] = 25'b00100000_00001101_00101101_0;
      patterns[8208] = 25'b00100000_00001110_00101110_0;
      patterns[8209] = 25'b00100000_00001111_00101111_0;
      patterns[8210] = 25'b00100000_00010000_00110000_0;
      patterns[8211] = 25'b00100000_00010001_00110001_0;
      patterns[8212] = 25'b00100000_00010010_00110010_0;
      patterns[8213] = 25'b00100000_00010011_00110011_0;
      patterns[8214] = 25'b00100000_00010100_00110100_0;
      patterns[8215] = 25'b00100000_00010101_00110101_0;
      patterns[8216] = 25'b00100000_00010110_00110110_0;
      patterns[8217] = 25'b00100000_00010111_00110111_0;
      patterns[8218] = 25'b00100000_00011000_00111000_0;
      patterns[8219] = 25'b00100000_00011001_00111001_0;
      patterns[8220] = 25'b00100000_00011010_00111010_0;
      patterns[8221] = 25'b00100000_00011011_00111011_0;
      patterns[8222] = 25'b00100000_00011100_00111100_0;
      patterns[8223] = 25'b00100000_00011101_00111101_0;
      patterns[8224] = 25'b00100000_00011110_00111110_0;
      patterns[8225] = 25'b00100000_00011111_00111111_0;
      patterns[8226] = 25'b00100000_00100000_01000000_0;
      patterns[8227] = 25'b00100000_00100001_01000001_0;
      patterns[8228] = 25'b00100000_00100010_01000010_0;
      patterns[8229] = 25'b00100000_00100011_01000011_0;
      patterns[8230] = 25'b00100000_00100100_01000100_0;
      patterns[8231] = 25'b00100000_00100101_01000101_0;
      patterns[8232] = 25'b00100000_00100110_01000110_0;
      patterns[8233] = 25'b00100000_00100111_01000111_0;
      patterns[8234] = 25'b00100000_00101000_01001000_0;
      patterns[8235] = 25'b00100000_00101001_01001001_0;
      patterns[8236] = 25'b00100000_00101010_01001010_0;
      patterns[8237] = 25'b00100000_00101011_01001011_0;
      patterns[8238] = 25'b00100000_00101100_01001100_0;
      patterns[8239] = 25'b00100000_00101101_01001101_0;
      patterns[8240] = 25'b00100000_00101110_01001110_0;
      patterns[8241] = 25'b00100000_00101111_01001111_0;
      patterns[8242] = 25'b00100000_00110000_01010000_0;
      patterns[8243] = 25'b00100000_00110001_01010001_0;
      patterns[8244] = 25'b00100000_00110010_01010010_0;
      patterns[8245] = 25'b00100000_00110011_01010011_0;
      patterns[8246] = 25'b00100000_00110100_01010100_0;
      patterns[8247] = 25'b00100000_00110101_01010101_0;
      patterns[8248] = 25'b00100000_00110110_01010110_0;
      patterns[8249] = 25'b00100000_00110111_01010111_0;
      patterns[8250] = 25'b00100000_00111000_01011000_0;
      patterns[8251] = 25'b00100000_00111001_01011001_0;
      patterns[8252] = 25'b00100000_00111010_01011010_0;
      patterns[8253] = 25'b00100000_00111011_01011011_0;
      patterns[8254] = 25'b00100000_00111100_01011100_0;
      patterns[8255] = 25'b00100000_00111101_01011101_0;
      patterns[8256] = 25'b00100000_00111110_01011110_0;
      patterns[8257] = 25'b00100000_00111111_01011111_0;
      patterns[8258] = 25'b00100000_01000000_01100000_0;
      patterns[8259] = 25'b00100000_01000001_01100001_0;
      patterns[8260] = 25'b00100000_01000010_01100010_0;
      patterns[8261] = 25'b00100000_01000011_01100011_0;
      patterns[8262] = 25'b00100000_01000100_01100100_0;
      patterns[8263] = 25'b00100000_01000101_01100101_0;
      patterns[8264] = 25'b00100000_01000110_01100110_0;
      patterns[8265] = 25'b00100000_01000111_01100111_0;
      patterns[8266] = 25'b00100000_01001000_01101000_0;
      patterns[8267] = 25'b00100000_01001001_01101001_0;
      patterns[8268] = 25'b00100000_01001010_01101010_0;
      patterns[8269] = 25'b00100000_01001011_01101011_0;
      patterns[8270] = 25'b00100000_01001100_01101100_0;
      patterns[8271] = 25'b00100000_01001101_01101101_0;
      patterns[8272] = 25'b00100000_01001110_01101110_0;
      patterns[8273] = 25'b00100000_01001111_01101111_0;
      patterns[8274] = 25'b00100000_01010000_01110000_0;
      patterns[8275] = 25'b00100000_01010001_01110001_0;
      patterns[8276] = 25'b00100000_01010010_01110010_0;
      patterns[8277] = 25'b00100000_01010011_01110011_0;
      patterns[8278] = 25'b00100000_01010100_01110100_0;
      patterns[8279] = 25'b00100000_01010101_01110101_0;
      patterns[8280] = 25'b00100000_01010110_01110110_0;
      patterns[8281] = 25'b00100000_01010111_01110111_0;
      patterns[8282] = 25'b00100000_01011000_01111000_0;
      patterns[8283] = 25'b00100000_01011001_01111001_0;
      patterns[8284] = 25'b00100000_01011010_01111010_0;
      patterns[8285] = 25'b00100000_01011011_01111011_0;
      patterns[8286] = 25'b00100000_01011100_01111100_0;
      patterns[8287] = 25'b00100000_01011101_01111101_0;
      patterns[8288] = 25'b00100000_01011110_01111110_0;
      patterns[8289] = 25'b00100000_01011111_01111111_0;
      patterns[8290] = 25'b00100000_01100000_10000000_0;
      patterns[8291] = 25'b00100000_01100001_10000001_0;
      patterns[8292] = 25'b00100000_01100010_10000010_0;
      patterns[8293] = 25'b00100000_01100011_10000011_0;
      patterns[8294] = 25'b00100000_01100100_10000100_0;
      patterns[8295] = 25'b00100000_01100101_10000101_0;
      patterns[8296] = 25'b00100000_01100110_10000110_0;
      patterns[8297] = 25'b00100000_01100111_10000111_0;
      patterns[8298] = 25'b00100000_01101000_10001000_0;
      patterns[8299] = 25'b00100000_01101001_10001001_0;
      patterns[8300] = 25'b00100000_01101010_10001010_0;
      patterns[8301] = 25'b00100000_01101011_10001011_0;
      patterns[8302] = 25'b00100000_01101100_10001100_0;
      patterns[8303] = 25'b00100000_01101101_10001101_0;
      patterns[8304] = 25'b00100000_01101110_10001110_0;
      patterns[8305] = 25'b00100000_01101111_10001111_0;
      patterns[8306] = 25'b00100000_01110000_10010000_0;
      patterns[8307] = 25'b00100000_01110001_10010001_0;
      patterns[8308] = 25'b00100000_01110010_10010010_0;
      patterns[8309] = 25'b00100000_01110011_10010011_0;
      patterns[8310] = 25'b00100000_01110100_10010100_0;
      patterns[8311] = 25'b00100000_01110101_10010101_0;
      patterns[8312] = 25'b00100000_01110110_10010110_0;
      patterns[8313] = 25'b00100000_01110111_10010111_0;
      patterns[8314] = 25'b00100000_01111000_10011000_0;
      patterns[8315] = 25'b00100000_01111001_10011001_0;
      patterns[8316] = 25'b00100000_01111010_10011010_0;
      patterns[8317] = 25'b00100000_01111011_10011011_0;
      patterns[8318] = 25'b00100000_01111100_10011100_0;
      patterns[8319] = 25'b00100000_01111101_10011101_0;
      patterns[8320] = 25'b00100000_01111110_10011110_0;
      patterns[8321] = 25'b00100000_01111111_10011111_0;
      patterns[8322] = 25'b00100000_10000000_10100000_0;
      patterns[8323] = 25'b00100000_10000001_10100001_0;
      patterns[8324] = 25'b00100000_10000010_10100010_0;
      patterns[8325] = 25'b00100000_10000011_10100011_0;
      patterns[8326] = 25'b00100000_10000100_10100100_0;
      patterns[8327] = 25'b00100000_10000101_10100101_0;
      patterns[8328] = 25'b00100000_10000110_10100110_0;
      patterns[8329] = 25'b00100000_10000111_10100111_0;
      patterns[8330] = 25'b00100000_10001000_10101000_0;
      patterns[8331] = 25'b00100000_10001001_10101001_0;
      patterns[8332] = 25'b00100000_10001010_10101010_0;
      patterns[8333] = 25'b00100000_10001011_10101011_0;
      patterns[8334] = 25'b00100000_10001100_10101100_0;
      patterns[8335] = 25'b00100000_10001101_10101101_0;
      patterns[8336] = 25'b00100000_10001110_10101110_0;
      patterns[8337] = 25'b00100000_10001111_10101111_0;
      patterns[8338] = 25'b00100000_10010000_10110000_0;
      patterns[8339] = 25'b00100000_10010001_10110001_0;
      patterns[8340] = 25'b00100000_10010010_10110010_0;
      patterns[8341] = 25'b00100000_10010011_10110011_0;
      patterns[8342] = 25'b00100000_10010100_10110100_0;
      patterns[8343] = 25'b00100000_10010101_10110101_0;
      patterns[8344] = 25'b00100000_10010110_10110110_0;
      patterns[8345] = 25'b00100000_10010111_10110111_0;
      patterns[8346] = 25'b00100000_10011000_10111000_0;
      patterns[8347] = 25'b00100000_10011001_10111001_0;
      patterns[8348] = 25'b00100000_10011010_10111010_0;
      patterns[8349] = 25'b00100000_10011011_10111011_0;
      patterns[8350] = 25'b00100000_10011100_10111100_0;
      patterns[8351] = 25'b00100000_10011101_10111101_0;
      patterns[8352] = 25'b00100000_10011110_10111110_0;
      patterns[8353] = 25'b00100000_10011111_10111111_0;
      patterns[8354] = 25'b00100000_10100000_11000000_0;
      patterns[8355] = 25'b00100000_10100001_11000001_0;
      patterns[8356] = 25'b00100000_10100010_11000010_0;
      patterns[8357] = 25'b00100000_10100011_11000011_0;
      patterns[8358] = 25'b00100000_10100100_11000100_0;
      patterns[8359] = 25'b00100000_10100101_11000101_0;
      patterns[8360] = 25'b00100000_10100110_11000110_0;
      patterns[8361] = 25'b00100000_10100111_11000111_0;
      patterns[8362] = 25'b00100000_10101000_11001000_0;
      patterns[8363] = 25'b00100000_10101001_11001001_0;
      patterns[8364] = 25'b00100000_10101010_11001010_0;
      patterns[8365] = 25'b00100000_10101011_11001011_0;
      patterns[8366] = 25'b00100000_10101100_11001100_0;
      patterns[8367] = 25'b00100000_10101101_11001101_0;
      patterns[8368] = 25'b00100000_10101110_11001110_0;
      patterns[8369] = 25'b00100000_10101111_11001111_0;
      patterns[8370] = 25'b00100000_10110000_11010000_0;
      patterns[8371] = 25'b00100000_10110001_11010001_0;
      patterns[8372] = 25'b00100000_10110010_11010010_0;
      patterns[8373] = 25'b00100000_10110011_11010011_0;
      patterns[8374] = 25'b00100000_10110100_11010100_0;
      patterns[8375] = 25'b00100000_10110101_11010101_0;
      patterns[8376] = 25'b00100000_10110110_11010110_0;
      patterns[8377] = 25'b00100000_10110111_11010111_0;
      patterns[8378] = 25'b00100000_10111000_11011000_0;
      patterns[8379] = 25'b00100000_10111001_11011001_0;
      patterns[8380] = 25'b00100000_10111010_11011010_0;
      patterns[8381] = 25'b00100000_10111011_11011011_0;
      patterns[8382] = 25'b00100000_10111100_11011100_0;
      patterns[8383] = 25'b00100000_10111101_11011101_0;
      patterns[8384] = 25'b00100000_10111110_11011110_0;
      patterns[8385] = 25'b00100000_10111111_11011111_0;
      patterns[8386] = 25'b00100000_11000000_11100000_0;
      patterns[8387] = 25'b00100000_11000001_11100001_0;
      patterns[8388] = 25'b00100000_11000010_11100010_0;
      patterns[8389] = 25'b00100000_11000011_11100011_0;
      patterns[8390] = 25'b00100000_11000100_11100100_0;
      patterns[8391] = 25'b00100000_11000101_11100101_0;
      patterns[8392] = 25'b00100000_11000110_11100110_0;
      patterns[8393] = 25'b00100000_11000111_11100111_0;
      patterns[8394] = 25'b00100000_11001000_11101000_0;
      patterns[8395] = 25'b00100000_11001001_11101001_0;
      patterns[8396] = 25'b00100000_11001010_11101010_0;
      patterns[8397] = 25'b00100000_11001011_11101011_0;
      patterns[8398] = 25'b00100000_11001100_11101100_0;
      patterns[8399] = 25'b00100000_11001101_11101101_0;
      patterns[8400] = 25'b00100000_11001110_11101110_0;
      patterns[8401] = 25'b00100000_11001111_11101111_0;
      patterns[8402] = 25'b00100000_11010000_11110000_0;
      patterns[8403] = 25'b00100000_11010001_11110001_0;
      patterns[8404] = 25'b00100000_11010010_11110010_0;
      patterns[8405] = 25'b00100000_11010011_11110011_0;
      patterns[8406] = 25'b00100000_11010100_11110100_0;
      patterns[8407] = 25'b00100000_11010101_11110101_0;
      patterns[8408] = 25'b00100000_11010110_11110110_0;
      patterns[8409] = 25'b00100000_11010111_11110111_0;
      patterns[8410] = 25'b00100000_11011000_11111000_0;
      patterns[8411] = 25'b00100000_11011001_11111001_0;
      patterns[8412] = 25'b00100000_11011010_11111010_0;
      patterns[8413] = 25'b00100000_11011011_11111011_0;
      patterns[8414] = 25'b00100000_11011100_11111100_0;
      patterns[8415] = 25'b00100000_11011101_11111101_0;
      patterns[8416] = 25'b00100000_11011110_11111110_0;
      patterns[8417] = 25'b00100000_11011111_11111111_0;
      patterns[8418] = 25'b00100000_11100000_00000000_1;
      patterns[8419] = 25'b00100000_11100001_00000001_1;
      patterns[8420] = 25'b00100000_11100010_00000010_1;
      patterns[8421] = 25'b00100000_11100011_00000011_1;
      patterns[8422] = 25'b00100000_11100100_00000100_1;
      patterns[8423] = 25'b00100000_11100101_00000101_1;
      patterns[8424] = 25'b00100000_11100110_00000110_1;
      patterns[8425] = 25'b00100000_11100111_00000111_1;
      patterns[8426] = 25'b00100000_11101000_00001000_1;
      patterns[8427] = 25'b00100000_11101001_00001001_1;
      patterns[8428] = 25'b00100000_11101010_00001010_1;
      patterns[8429] = 25'b00100000_11101011_00001011_1;
      patterns[8430] = 25'b00100000_11101100_00001100_1;
      patterns[8431] = 25'b00100000_11101101_00001101_1;
      patterns[8432] = 25'b00100000_11101110_00001110_1;
      patterns[8433] = 25'b00100000_11101111_00001111_1;
      patterns[8434] = 25'b00100000_11110000_00010000_1;
      patterns[8435] = 25'b00100000_11110001_00010001_1;
      patterns[8436] = 25'b00100000_11110010_00010010_1;
      patterns[8437] = 25'b00100000_11110011_00010011_1;
      patterns[8438] = 25'b00100000_11110100_00010100_1;
      patterns[8439] = 25'b00100000_11110101_00010101_1;
      patterns[8440] = 25'b00100000_11110110_00010110_1;
      patterns[8441] = 25'b00100000_11110111_00010111_1;
      patterns[8442] = 25'b00100000_11111000_00011000_1;
      patterns[8443] = 25'b00100000_11111001_00011001_1;
      patterns[8444] = 25'b00100000_11111010_00011010_1;
      patterns[8445] = 25'b00100000_11111011_00011011_1;
      patterns[8446] = 25'b00100000_11111100_00011100_1;
      patterns[8447] = 25'b00100000_11111101_00011101_1;
      patterns[8448] = 25'b00100000_11111110_00011110_1;
      patterns[8449] = 25'b00100000_11111111_00011111_1;
      patterns[8450] = 25'b00100001_00000000_00100001_0;
      patterns[8451] = 25'b00100001_00000001_00100010_0;
      patterns[8452] = 25'b00100001_00000010_00100011_0;
      patterns[8453] = 25'b00100001_00000011_00100100_0;
      patterns[8454] = 25'b00100001_00000100_00100101_0;
      patterns[8455] = 25'b00100001_00000101_00100110_0;
      patterns[8456] = 25'b00100001_00000110_00100111_0;
      patterns[8457] = 25'b00100001_00000111_00101000_0;
      patterns[8458] = 25'b00100001_00001000_00101001_0;
      patterns[8459] = 25'b00100001_00001001_00101010_0;
      patterns[8460] = 25'b00100001_00001010_00101011_0;
      patterns[8461] = 25'b00100001_00001011_00101100_0;
      patterns[8462] = 25'b00100001_00001100_00101101_0;
      patterns[8463] = 25'b00100001_00001101_00101110_0;
      patterns[8464] = 25'b00100001_00001110_00101111_0;
      patterns[8465] = 25'b00100001_00001111_00110000_0;
      patterns[8466] = 25'b00100001_00010000_00110001_0;
      patterns[8467] = 25'b00100001_00010001_00110010_0;
      patterns[8468] = 25'b00100001_00010010_00110011_0;
      patterns[8469] = 25'b00100001_00010011_00110100_0;
      patterns[8470] = 25'b00100001_00010100_00110101_0;
      patterns[8471] = 25'b00100001_00010101_00110110_0;
      patterns[8472] = 25'b00100001_00010110_00110111_0;
      patterns[8473] = 25'b00100001_00010111_00111000_0;
      patterns[8474] = 25'b00100001_00011000_00111001_0;
      patterns[8475] = 25'b00100001_00011001_00111010_0;
      patterns[8476] = 25'b00100001_00011010_00111011_0;
      patterns[8477] = 25'b00100001_00011011_00111100_0;
      patterns[8478] = 25'b00100001_00011100_00111101_0;
      patterns[8479] = 25'b00100001_00011101_00111110_0;
      patterns[8480] = 25'b00100001_00011110_00111111_0;
      patterns[8481] = 25'b00100001_00011111_01000000_0;
      patterns[8482] = 25'b00100001_00100000_01000001_0;
      patterns[8483] = 25'b00100001_00100001_01000010_0;
      patterns[8484] = 25'b00100001_00100010_01000011_0;
      patterns[8485] = 25'b00100001_00100011_01000100_0;
      patterns[8486] = 25'b00100001_00100100_01000101_0;
      patterns[8487] = 25'b00100001_00100101_01000110_0;
      patterns[8488] = 25'b00100001_00100110_01000111_0;
      patterns[8489] = 25'b00100001_00100111_01001000_0;
      patterns[8490] = 25'b00100001_00101000_01001001_0;
      patterns[8491] = 25'b00100001_00101001_01001010_0;
      patterns[8492] = 25'b00100001_00101010_01001011_0;
      patterns[8493] = 25'b00100001_00101011_01001100_0;
      patterns[8494] = 25'b00100001_00101100_01001101_0;
      patterns[8495] = 25'b00100001_00101101_01001110_0;
      patterns[8496] = 25'b00100001_00101110_01001111_0;
      patterns[8497] = 25'b00100001_00101111_01010000_0;
      patterns[8498] = 25'b00100001_00110000_01010001_0;
      patterns[8499] = 25'b00100001_00110001_01010010_0;
      patterns[8500] = 25'b00100001_00110010_01010011_0;
      patterns[8501] = 25'b00100001_00110011_01010100_0;
      patterns[8502] = 25'b00100001_00110100_01010101_0;
      patterns[8503] = 25'b00100001_00110101_01010110_0;
      patterns[8504] = 25'b00100001_00110110_01010111_0;
      patterns[8505] = 25'b00100001_00110111_01011000_0;
      patterns[8506] = 25'b00100001_00111000_01011001_0;
      patterns[8507] = 25'b00100001_00111001_01011010_0;
      patterns[8508] = 25'b00100001_00111010_01011011_0;
      patterns[8509] = 25'b00100001_00111011_01011100_0;
      patterns[8510] = 25'b00100001_00111100_01011101_0;
      patterns[8511] = 25'b00100001_00111101_01011110_0;
      patterns[8512] = 25'b00100001_00111110_01011111_0;
      patterns[8513] = 25'b00100001_00111111_01100000_0;
      patterns[8514] = 25'b00100001_01000000_01100001_0;
      patterns[8515] = 25'b00100001_01000001_01100010_0;
      patterns[8516] = 25'b00100001_01000010_01100011_0;
      patterns[8517] = 25'b00100001_01000011_01100100_0;
      patterns[8518] = 25'b00100001_01000100_01100101_0;
      patterns[8519] = 25'b00100001_01000101_01100110_0;
      patterns[8520] = 25'b00100001_01000110_01100111_0;
      patterns[8521] = 25'b00100001_01000111_01101000_0;
      patterns[8522] = 25'b00100001_01001000_01101001_0;
      patterns[8523] = 25'b00100001_01001001_01101010_0;
      patterns[8524] = 25'b00100001_01001010_01101011_0;
      patterns[8525] = 25'b00100001_01001011_01101100_0;
      patterns[8526] = 25'b00100001_01001100_01101101_0;
      patterns[8527] = 25'b00100001_01001101_01101110_0;
      patterns[8528] = 25'b00100001_01001110_01101111_0;
      patterns[8529] = 25'b00100001_01001111_01110000_0;
      patterns[8530] = 25'b00100001_01010000_01110001_0;
      patterns[8531] = 25'b00100001_01010001_01110010_0;
      patterns[8532] = 25'b00100001_01010010_01110011_0;
      patterns[8533] = 25'b00100001_01010011_01110100_0;
      patterns[8534] = 25'b00100001_01010100_01110101_0;
      patterns[8535] = 25'b00100001_01010101_01110110_0;
      patterns[8536] = 25'b00100001_01010110_01110111_0;
      patterns[8537] = 25'b00100001_01010111_01111000_0;
      patterns[8538] = 25'b00100001_01011000_01111001_0;
      patterns[8539] = 25'b00100001_01011001_01111010_0;
      patterns[8540] = 25'b00100001_01011010_01111011_0;
      patterns[8541] = 25'b00100001_01011011_01111100_0;
      patterns[8542] = 25'b00100001_01011100_01111101_0;
      patterns[8543] = 25'b00100001_01011101_01111110_0;
      patterns[8544] = 25'b00100001_01011110_01111111_0;
      patterns[8545] = 25'b00100001_01011111_10000000_0;
      patterns[8546] = 25'b00100001_01100000_10000001_0;
      patterns[8547] = 25'b00100001_01100001_10000010_0;
      patterns[8548] = 25'b00100001_01100010_10000011_0;
      patterns[8549] = 25'b00100001_01100011_10000100_0;
      patterns[8550] = 25'b00100001_01100100_10000101_0;
      patterns[8551] = 25'b00100001_01100101_10000110_0;
      patterns[8552] = 25'b00100001_01100110_10000111_0;
      patterns[8553] = 25'b00100001_01100111_10001000_0;
      patterns[8554] = 25'b00100001_01101000_10001001_0;
      patterns[8555] = 25'b00100001_01101001_10001010_0;
      patterns[8556] = 25'b00100001_01101010_10001011_0;
      patterns[8557] = 25'b00100001_01101011_10001100_0;
      patterns[8558] = 25'b00100001_01101100_10001101_0;
      patterns[8559] = 25'b00100001_01101101_10001110_0;
      patterns[8560] = 25'b00100001_01101110_10001111_0;
      patterns[8561] = 25'b00100001_01101111_10010000_0;
      patterns[8562] = 25'b00100001_01110000_10010001_0;
      patterns[8563] = 25'b00100001_01110001_10010010_0;
      patterns[8564] = 25'b00100001_01110010_10010011_0;
      patterns[8565] = 25'b00100001_01110011_10010100_0;
      patterns[8566] = 25'b00100001_01110100_10010101_0;
      patterns[8567] = 25'b00100001_01110101_10010110_0;
      patterns[8568] = 25'b00100001_01110110_10010111_0;
      patterns[8569] = 25'b00100001_01110111_10011000_0;
      patterns[8570] = 25'b00100001_01111000_10011001_0;
      patterns[8571] = 25'b00100001_01111001_10011010_0;
      patterns[8572] = 25'b00100001_01111010_10011011_0;
      patterns[8573] = 25'b00100001_01111011_10011100_0;
      patterns[8574] = 25'b00100001_01111100_10011101_0;
      patterns[8575] = 25'b00100001_01111101_10011110_0;
      patterns[8576] = 25'b00100001_01111110_10011111_0;
      patterns[8577] = 25'b00100001_01111111_10100000_0;
      patterns[8578] = 25'b00100001_10000000_10100001_0;
      patterns[8579] = 25'b00100001_10000001_10100010_0;
      patterns[8580] = 25'b00100001_10000010_10100011_0;
      patterns[8581] = 25'b00100001_10000011_10100100_0;
      patterns[8582] = 25'b00100001_10000100_10100101_0;
      patterns[8583] = 25'b00100001_10000101_10100110_0;
      patterns[8584] = 25'b00100001_10000110_10100111_0;
      patterns[8585] = 25'b00100001_10000111_10101000_0;
      patterns[8586] = 25'b00100001_10001000_10101001_0;
      patterns[8587] = 25'b00100001_10001001_10101010_0;
      patterns[8588] = 25'b00100001_10001010_10101011_0;
      patterns[8589] = 25'b00100001_10001011_10101100_0;
      patterns[8590] = 25'b00100001_10001100_10101101_0;
      patterns[8591] = 25'b00100001_10001101_10101110_0;
      patterns[8592] = 25'b00100001_10001110_10101111_0;
      patterns[8593] = 25'b00100001_10001111_10110000_0;
      patterns[8594] = 25'b00100001_10010000_10110001_0;
      patterns[8595] = 25'b00100001_10010001_10110010_0;
      patterns[8596] = 25'b00100001_10010010_10110011_0;
      patterns[8597] = 25'b00100001_10010011_10110100_0;
      patterns[8598] = 25'b00100001_10010100_10110101_0;
      patterns[8599] = 25'b00100001_10010101_10110110_0;
      patterns[8600] = 25'b00100001_10010110_10110111_0;
      patterns[8601] = 25'b00100001_10010111_10111000_0;
      patterns[8602] = 25'b00100001_10011000_10111001_0;
      patterns[8603] = 25'b00100001_10011001_10111010_0;
      patterns[8604] = 25'b00100001_10011010_10111011_0;
      patterns[8605] = 25'b00100001_10011011_10111100_0;
      patterns[8606] = 25'b00100001_10011100_10111101_0;
      patterns[8607] = 25'b00100001_10011101_10111110_0;
      patterns[8608] = 25'b00100001_10011110_10111111_0;
      patterns[8609] = 25'b00100001_10011111_11000000_0;
      patterns[8610] = 25'b00100001_10100000_11000001_0;
      patterns[8611] = 25'b00100001_10100001_11000010_0;
      patterns[8612] = 25'b00100001_10100010_11000011_0;
      patterns[8613] = 25'b00100001_10100011_11000100_0;
      patterns[8614] = 25'b00100001_10100100_11000101_0;
      patterns[8615] = 25'b00100001_10100101_11000110_0;
      patterns[8616] = 25'b00100001_10100110_11000111_0;
      patterns[8617] = 25'b00100001_10100111_11001000_0;
      patterns[8618] = 25'b00100001_10101000_11001001_0;
      patterns[8619] = 25'b00100001_10101001_11001010_0;
      patterns[8620] = 25'b00100001_10101010_11001011_0;
      patterns[8621] = 25'b00100001_10101011_11001100_0;
      patterns[8622] = 25'b00100001_10101100_11001101_0;
      patterns[8623] = 25'b00100001_10101101_11001110_0;
      patterns[8624] = 25'b00100001_10101110_11001111_0;
      patterns[8625] = 25'b00100001_10101111_11010000_0;
      patterns[8626] = 25'b00100001_10110000_11010001_0;
      patterns[8627] = 25'b00100001_10110001_11010010_0;
      patterns[8628] = 25'b00100001_10110010_11010011_0;
      patterns[8629] = 25'b00100001_10110011_11010100_0;
      patterns[8630] = 25'b00100001_10110100_11010101_0;
      patterns[8631] = 25'b00100001_10110101_11010110_0;
      patterns[8632] = 25'b00100001_10110110_11010111_0;
      patterns[8633] = 25'b00100001_10110111_11011000_0;
      patterns[8634] = 25'b00100001_10111000_11011001_0;
      patterns[8635] = 25'b00100001_10111001_11011010_0;
      patterns[8636] = 25'b00100001_10111010_11011011_0;
      patterns[8637] = 25'b00100001_10111011_11011100_0;
      patterns[8638] = 25'b00100001_10111100_11011101_0;
      patterns[8639] = 25'b00100001_10111101_11011110_0;
      patterns[8640] = 25'b00100001_10111110_11011111_0;
      patterns[8641] = 25'b00100001_10111111_11100000_0;
      patterns[8642] = 25'b00100001_11000000_11100001_0;
      patterns[8643] = 25'b00100001_11000001_11100010_0;
      patterns[8644] = 25'b00100001_11000010_11100011_0;
      patterns[8645] = 25'b00100001_11000011_11100100_0;
      patterns[8646] = 25'b00100001_11000100_11100101_0;
      patterns[8647] = 25'b00100001_11000101_11100110_0;
      patterns[8648] = 25'b00100001_11000110_11100111_0;
      patterns[8649] = 25'b00100001_11000111_11101000_0;
      patterns[8650] = 25'b00100001_11001000_11101001_0;
      patterns[8651] = 25'b00100001_11001001_11101010_0;
      patterns[8652] = 25'b00100001_11001010_11101011_0;
      patterns[8653] = 25'b00100001_11001011_11101100_0;
      patterns[8654] = 25'b00100001_11001100_11101101_0;
      patterns[8655] = 25'b00100001_11001101_11101110_0;
      patterns[8656] = 25'b00100001_11001110_11101111_0;
      patterns[8657] = 25'b00100001_11001111_11110000_0;
      patterns[8658] = 25'b00100001_11010000_11110001_0;
      patterns[8659] = 25'b00100001_11010001_11110010_0;
      patterns[8660] = 25'b00100001_11010010_11110011_0;
      patterns[8661] = 25'b00100001_11010011_11110100_0;
      patterns[8662] = 25'b00100001_11010100_11110101_0;
      patterns[8663] = 25'b00100001_11010101_11110110_0;
      patterns[8664] = 25'b00100001_11010110_11110111_0;
      patterns[8665] = 25'b00100001_11010111_11111000_0;
      patterns[8666] = 25'b00100001_11011000_11111001_0;
      patterns[8667] = 25'b00100001_11011001_11111010_0;
      patterns[8668] = 25'b00100001_11011010_11111011_0;
      patterns[8669] = 25'b00100001_11011011_11111100_0;
      patterns[8670] = 25'b00100001_11011100_11111101_0;
      patterns[8671] = 25'b00100001_11011101_11111110_0;
      patterns[8672] = 25'b00100001_11011110_11111111_0;
      patterns[8673] = 25'b00100001_11011111_00000000_1;
      patterns[8674] = 25'b00100001_11100000_00000001_1;
      patterns[8675] = 25'b00100001_11100001_00000010_1;
      patterns[8676] = 25'b00100001_11100010_00000011_1;
      patterns[8677] = 25'b00100001_11100011_00000100_1;
      patterns[8678] = 25'b00100001_11100100_00000101_1;
      patterns[8679] = 25'b00100001_11100101_00000110_1;
      patterns[8680] = 25'b00100001_11100110_00000111_1;
      patterns[8681] = 25'b00100001_11100111_00001000_1;
      patterns[8682] = 25'b00100001_11101000_00001001_1;
      patterns[8683] = 25'b00100001_11101001_00001010_1;
      patterns[8684] = 25'b00100001_11101010_00001011_1;
      patterns[8685] = 25'b00100001_11101011_00001100_1;
      patterns[8686] = 25'b00100001_11101100_00001101_1;
      patterns[8687] = 25'b00100001_11101101_00001110_1;
      patterns[8688] = 25'b00100001_11101110_00001111_1;
      patterns[8689] = 25'b00100001_11101111_00010000_1;
      patterns[8690] = 25'b00100001_11110000_00010001_1;
      patterns[8691] = 25'b00100001_11110001_00010010_1;
      patterns[8692] = 25'b00100001_11110010_00010011_1;
      patterns[8693] = 25'b00100001_11110011_00010100_1;
      patterns[8694] = 25'b00100001_11110100_00010101_1;
      patterns[8695] = 25'b00100001_11110101_00010110_1;
      patterns[8696] = 25'b00100001_11110110_00010111_1;
      patterns[8697] = 25'b00100001_11110111_00011000_1;
      patterns[8698] = 25'b00100001_11111000_00011001_1;
      patterns[8699] = 25'b00100001_11111001_00011010_1;
      patterns[8700] = 25'b00100001_11111010_00011011_1;
      patterns[8701] = 25'b00100001_11111011_00011100_1;
      patterns[8702] = 25'b00100001_11111100_00011101_1;
      patterns[8703] = 25'b00100001_11111101_00011110_1;
      patterns[8704] = 25'b00100001_11111110_00011111_1;
      patterns[8705] = 25'b00100001_11111111_00100000_1;
      patterns[8706] = 25'b00100010_00000000_00100010_0;
      patterns[8707] = 25'b00100010_00000001_00100011_0;
      patterns[8708] = 25'b00100010_00000010_00100100_0;
      patterns[8709] = 25'b00100010_00000011_00100101_0;
      patterns[8710] = 25'b00100010_00000100_00100110_0;
      patterns[8711] = 25'b00100010_00000101_00100111_0;
      patterns[8712] = 25'b00100010_00000110_00101000_0;
      patterns[8713] = 25'b00100010_00000111_00101001_0;
      patterns[8714] = 25'b00100010_00001000_00101010_0;
      patterns[8715] = 25'b00100010_00001001_00101011_0;
      patterns[8716] = 25'b00100010_00001010_00101100_0;
      patterns[8717] = 25'b00100010_00001011_00101101_0;
      patterns[8718] = 25'b00100010_00001100_00101110_0;
      patterns[8719] = 25'b00100010_00001101_00101111_0;
      patterns[8720] = 25'b00100010_00001110_00110000_0;
      patterns[8721] = 25'b00100010_00001111_00110001_0;
      patterns[8722] = 25'b00100010_00010000_00110010_0;
      patterns[8723] = 25'b00100010_00010001_00110011_0;
      patterns[8724] = 25'b00100010_00010010_00110100_0;
      patterns[8725] = 25'b00100010_00010011_00110101_0;
      patterns[8726] = 25'b00100010_00010100_00110110_0;
      patterns[8727] = 25'b00100010_00010101_00110111_0;
      patterns[8728] = 25'b00100010_00010110_00111000_0;
      patterns[8729] = 25'b00100010_00010111_00111001_0;
      patterns[8730] = 25'b00100010_00011000_00111010_0;
      patterns[8731] = 25'b00100010_00011001_00111011_0;
      patterns[8732] = 25'b00100010_00011010_00111100_0;
      patterns[8733] = 25'b00100010_00011011_00111101_0;
      patterns[8734] = 25'b00100010_00011100_00111110_0;
      patterns[8735] = 25'b00100010_00011101_00111111_0;
      patterns[8736] = 25'b00100010_00011110_01000000_0;
      patterns[8737] = 25'b00100010_00011111_01000001_0;
      patterns[8738] = 25'b00100010_00100000_01000010_0;
      patterns[8739] = 25'b00100010_00100001_01000011_0;
      patterns[8740] = 25'b00100010_00100010_01000100_0;
      patterns[8741] = 25'b00100010_00100011_01000101_0;
      patterns[8742] = 25'b00100010_00100100_01000110_0;
      patterns[8743] = 25'b00100010_00100101_01000111_0;
      patterns[8744] = 25'b00100010_00100110_01001000_0;
      patterns[8745] = 25'b00100010_00100111_01001001_0;
      patterns[8746] = 25'b00100010_00101000_01001010_0;
      patterns[8747] = 25'b00100010_00101001_01001011_0;
      patterns[8748] = 25'b00100010_00101010_01001100_0;
      patterns[8749] = 25'b00100010_00101011_01001101_0;
      patterns[8750] = 25'b00100010_00101100_01001110_0;
      patterns[8751] = 25'b00100010_00101101_01001111_0;
      patterns[8752] = 25'b00100010_00101110_01010000_0;
      patterns[8753] = 25'b00100010_00101111_01010001_0;
      patterns[8754] = 25'b00100010_00110000_01010010_0;
      patterns[8755] = 25'b00100010_00110001_01010011_0;
      patterns[8756] = 25'b00100010_00110010_01010100_0;
      patterns[8757] = 25'b00100010_00110011_01010101_0;
      patterns[8758] = 25'b00100010_00110100_01010110_0;
      patterns[8759] = 25'b00100010_00110101_01010111_0;
      patterns[8760] = 25'b00100010_00110110_01011000_0;
      patterns[8761] = 25'b00100010_00110111_01011001_0;
      patterns[8762] = 25'b00100010_00111000_01011010_0;
      patterns[8763] = 25'b00100010_00111001_01011011_0;
      patterns[8764] = 25'b00100010_00111010_01011100_0;
      patterns[8765] = 25'b00100010_00111011_01011101_0;
      patterns[8766] = 25'b00100010_00111100_01011110_0;
      patterns[8767] = 25'b00100010_00111101_01011111_0;
      patterns[8768] = 25'b00100010_00111110_01100000_0;
      patterns[8769] = 25'b00100010_00111111_01100001_0;
      patterns[8770] = 25'b00100010_01000000_01100010_0;
      patterns[8771] = 25'b00100010_01000001_01100011_0;
      patterns[8772] = 25'b00100010_01000010_01100100_0;
      patterns[8773] = 25'b00100010_01000011_01100101_0;
      patterns[8774] = 25'b00100010_01000100_01100110_0;
      patterns[8775] = 25'b00100010_01000101_01100111_0;
      patterns[8776] = 25'b00100010_01000110_01101000_0;
      patterns[8777] = 25'b00100010_01000111_01101001_0;
      patterns[8778] = 25'b00100010_01001000_01101010_0;
      patterns[8779] = 25'b00100010_01001001_01101011_0;
      patterns[8780] = 25'b00100010_01001010_01101100_0;
      patterns[8781] = 25'b00100010_01001011_01101101_0;
      patterns[8782] = 25'b00100010_01001100_01101110_0;
      patterns[8783] = 25'b00100010_01001101_01101111_0;
      patterns[8784] = 25'b00100010_01001110_01110000_0;
      patterns[8785] = 25'b00100010_01001111_01110001_0;
      patterns[8786] = 25'b00100010_01010000_01110010_0;
      patterns[8787] = 25'b00100010_01010001_01110011_0;
      patterns[8788] = 25'b00100010_01010010_01110100_0;
      patterns[8789] = 25'b00100010_01010011_01110101_0;
      patterns[8790] = 25'b00100010_01010100_01110110_0;
      patterns[8791] = 25'b00100010_01010101_01110111_0;
      patterns[8792] = 25'b00100010_01010110_01111000_0;
      patterns[8793] = 25'b00100010_01010111_01111001_0;
      patterns[8794] = 25'b00100010_01011000_01111010_0;
      patterns[8795] = 25'b00100010_01011001_01111011_0;
      patterns[8796] = 25'b00100010_01011010_01111100_0;
      patterns[8797] = 25'b00100010_01011011_01111101_0;
      patterns[8798] = 25'b00100010_01011100_01111110_0;
      patterns[8799] = 25'b00100010_01011101_01111111_0;
      patterns[8800] = 25'b00100010_01011110_10000000_0;
      patterns[8801] = 25'b00100010_01011111_10000001_0;
      patterns[8802] = 25'b00100010_01100000_10000010_0;
      patterns[8803] = 25'b00100010_01100001_10000011_0;
      patterns[8804] = 25'b00100010_01100010_10000100_0;
      patterns[8805] = 25'b00100010_01100011_10000101_0;
      patterns[8806] = 25'b00100010_01100100_10000110_0;
      patterns[8807] = 25'b00100010_01100101_10000111_0;
      patterns[8808] = 25'b00100010_01100110_10001000_0;
      patterns[8809] = 25'b00100010_01100111_10001001_0;
      patterns[8810] = 25'b00100010_01101000_10001010_0;
      patterns[8811] = 25'b00100010_01101001_10001011_0;
      patterns[8812] = 25'b00100010_01101010_10001100_0;
      patterns[8813] = 25'b00100010_01101011_10001101_0;
      patterns[8814] = 25'b00100010_01101100_10001110_0;
      patterns[8815] = 25'b00100010_01101101_10001111_0;
      patterns[8816] = 25'b00100010_01101110_10010000_0;
      patterns[8817] = 25'b00100010_01101111_10010001_0;
      patterns[8818] = 25'b00100010_01110000_10010010_0;
      patterns[8819] = 25'b00100010_01110001_10010011_0;
      patterns[8820] = 25'b00100010_01110010_10010100_0;
      patterns[8821] = 25'b00100010_01110011_10010101_0;
      patterns[8822] = 25'b00100010_01110100_10010110_0;
      patterns[8823] = 25'b00100010_01110101_10010111_0;
      patterns[8824] = 25'b00100010_01110110_10011000_0;
      patterns[8825] = 25'b00100010_01110111_10011001_0;
      patterns[8826] = 25'b00100010_01111000_10011010_0;
      patterns[8827] = 25'b00100010_01111001_10011011_0;
      patterns[8828] = 25'b00100010_01111010_10011100_0;
      patterns[8829] = 25'b00100010_01111011_10011101_0;
      patterns[8830] = 25'b00100010_01111100_10011110_0;
      patterns[8831] = 25'b00100010_01111101_10011111_0;
      patterns[8832] = 25'b00100010_01111110_10100000_0;
      patterns[8833] = 25'b00100010_01111111_10100001_0;
      patterns[8834] = 25'b00100010_10000000_10100010_0;
      patterns[8835] = 25'b00100010_10000001_10100011_0;
      patterns[8836] = 25'b00100010_10000010_10100100_0;
      patterns[8837] = 25'b00100010_10000011_10100101_0;
      patterns[8838] = 25'b00100010_10000100_10100110_0;
      patterns[8839] = 25'b00100010_10000101_10100111_0;
      patterns[8840] = 25'b00100010_10000110_10101000_0;
      patterns[8841] = 25'b00100010_10000111_10101001_0;
      patterns[8842] = 25'b00100010_10001000_10101010_0;
      patterns[8843] = 25'b00100010_10001001_10101011_0;
      patterns[8844] = 25'b00100010_10001010_10101100_0;
      patterns[8845] = 25'b00100010_10001011_10101101_0;
      patterns[8846] = 25'b00100010_10001100_10101110_0;
      patterns[8847] = 25'b00100010_10001101_10101111_0;
      patterns[8848] = 25'b00100010_10001110_10110000_0;
      patterns[8849] = 25'b00100010_10001111_10110001_0;
      patterns[8850] = 25'b00100010_10010000_10110010_0;
      patterns[8851] = 25'b00100010_10010001_10110011_0;
      patterns[8852] = 25'b00100010_10010010_10110100_0;
      patterns[8853] = 25'b00100010_10010011_10110101_0;
      patterns[8854] = 25'b00100010_10010100_10110110_0;
      patterns[8855] = 25'b00100010_10010101_10110111_0;
      patterns[8856] = 25'b00100010_10010110_10111000_0;
      patterns[8857] = 25'b00100010_10010111_10111001_0;
      patterns[8858] = 25'b00100010_10011000_10111010_0;
      patterns[8859] = 25'b00100010_10011001_10111011_0;
      patterns[8860] = 25'b00100010_10011010_10111100_0;
      patterns[8861] = 25'b00100010_10011011_10111101_0;
      patterns[8862] = 25'b00100010_10011100_10111110_0;
      patterns[8863] = 25'b00100010_10011101_10111111_0;
      patterns[8864] = 25'b00100010_10011110_11000000_0;
      patterns[8865] = 25'b00100010_10011111_11000001_0;
      patterns[8866] = 25'b00100010_10100000_11000010_0;
      patterns[8867] = 25'b00100010_10100001_11000011_0;
      patterns[8868] = 25'b00100010_10100010_11000100_0;
      patterns[8869] = 25'b00100010_10100011_11000101_0;
      patterns[8870] = 25'b00100010_10100100_11000110_0;
      patterns[8871] = 25'b00100010_10100101_11000111_0;
      patterns[8872] = 25'b00100010_10100110_11001000_0;
      patterns[8873] = 25'b00100010_10100111_11001001_0;
      patterns[8874] = 25'b00100010_10101000_11001010_0;
      patterns[8875] = 25'b00100010_10101001_11001011_0;
      patterns[8876] = 25'b00100010_10101010_11001100_0;
      patterns[8877] = 25'b00100010_10101011_11001101_0;
      patterns[8878] = 25'b00100010_10101100_11001110_0;
      patterns[8879] = 25'b00100010_10101101_11001111_0;
      patterns[8880] = 25'b00100010_10101110_11010000_0;
      patterns[8881] = 25'b00100010_10101111_11010001_0;
      patterns[8882] = 25'b00100010_10110000_11010010_0;
      patterns[8883] = 25'b00100010_10110001_11010011_0;
      patterns[8884] = 25'b00100010_10110010_11010100_0;
      patterns[8885] = 25'b00100010_10110011_11010101_0;
      patterns[8886] = 25'b00100010_10110100_11010110_0;
      patterns[8887] = 25'b00100010_10110101_11010111_0;
      patterns[8888] = 25'b00100010_10110110_11011000_0;
      patterns[8889] = 25'b00100010_10110111_11011001_0;
      patterns[8890] = 25'b00100010_10111000_11011010_0;
      patterns[8891] = 25'b00100010_10111001_11011011_0;
      patterns[8892] = 25'b00100010_10111010_11011100_0;
      patterns[8893] = 25'b00100010_10111011_11011101_0;
      patterns[8894] = 25'b00100010_10111100_11011110_0;
      patterns[8895] = 25'b00100010_10111101_11011111_0;
      patterns[8896] = 25'b00100010_10111110_11100000_0;
      patterns[8897] = 25'b00100010_10111111_11100001_0;
      patterns[8898] = 25'b00100010_11000000_11100010_0;
      patterns[8899] = 25'b00100010_11000001_11100011_0;
      patterns[8900] = 25'b00100010_11000010_11100100_0;
      patterns[8901] = 25'b00100010_11000011_11100101_0;
      patterns[8902] = 25'b00100010_11000100_11100110_0;
      patterns[8903] = 25'b00100010_11000101_11100111_0;
      patterns[8904] = 25'b00100010_11000110_11101000_0;
      patterns[8905] = 25'b00100010_11000111_11101001_0;
      patterns[8906] = 25'b00100010_11001000_11101010_0;
      patterns[8907] = 25'b00100010_11001001_11101011_0;
      patterns[8908] = 25'b00100010_11001010_11101100_0;
      patterns[8909] = 25'b00100010_11001011_11101101_0;
      patterns[8910] = 25'b00100010_11001100_11101110_0;
      patterns[8911] = 25'b00100010_11001101_11101111_0;
      patterns[8912] = 25'b00100010_11001110_11110000_0;
      patterns[8913] = 25'b00100010_11001111_11110001_0;
      patterns[8914] = 25'b00100010_11010000_11110010_0;
      patterns[8915] = 25'b00100010_11010001_11110011_0;
      patterns[8916] = 25'b00100010_11010010_11110100_0;
      patterns[8917] = 25'b00100010_11010011_11110101_0;
      patterns[8918] = 25'b00100010_11010100_11110110_0;
      patterns[8919] = 25'b00100010_11010101_11110111_0;
      patterns[8920] = 25'b00100010_11010110_11111000_0;
      patterns[8921] = 25'b00100010_11010111_11111001_0;
      patterns[8922] = 25'b00100010_11011000_11111010_0;
      patterns[8923] = 25'b00100010_11011001_11111011_0;
      patterns[8924] = 25'b00100010_11011010_11111100_0;
      patterns[8925] = 25'b00100010_11011011_11111101_0;
      patterns[8926] = 25'b00100010_11011100_11111110_0;
      patterns[8927] = 25'b00100010_11011101_11111111_0;
      patterns[8928] = 25'b00100010_11011110_00000000_1;
      patterns[8929] = 25'b00100010_11011111_00000001_1;
      patterns[8930] = 25'b00100010_11100000_00000010_1;
      patterns[8931] = 25'b00100010_11100001_00000011_1;
      patterns[8932] = 25'b00100010_11100010_00000100_1;
      patterns[8933] = 25'b00100010_11100011_00000101_1;
      patterns[8934] = 25'b00100010_11100100_00000110_1;
      patterns[8935] = 25'b00100010_11100101_00000111_1;
      patterns[8936] = 25'b00100010_11100110_00001000_1;
      patterns[8937] = 25'b00100010_11100111_00001001_1;
      patterns[8938] = 25'b00100010_11101000_00001010_1;
      patterns[8939] = 25'b00100010_11101001_00001011_1;
      patterns[8940] = 25'b00100010_11101010_00001100_1;
      patterns[8941] = 25'b00100010_11101011_00001101_1;
      patterns[8942] = 25'b00100010_11101100_00001110_1;
      patterns[8943] = 25'b00100010_11101101_00001111_1;
      patterns[8944] = 25'b00100010_11101110_00010000_1;
      patterns[8945] = 25'b00100010_11101111_00010001_1;
      patterns[8946] = 25'b00100010_11110000_00010010_1;
      patterns[8947] = 25'b00100010_11110001_00010011_1;
      patterns[8948] = 25'b00100010_11110010_00010100_1;
      patterns[8949] = 25'b00100010_11110011_00010101_1;
      patterns[8950] = 25'b00100010_11110100_00010110_1;
      patterns[8951] = 25'b00100010_11110101_00010111_1;
      patterns[8952] = 25'b00100010_11110110_00011000_1;
      patterns[8953] = 25'b00100010_11110111_00011001_1;
      patterns[8954] = 25'b00100010_11111000_00011010_1;
      patterns[8955] = 25'b00100010_11111001_00011011_1;
      patterns[8956] = 25'b00100010_11111010_00011100_1;
      patterns[8957] = 25'b00100010_11111011_00011101_1;
      patterns[8958] = 25'b00100010_11111100_00011110_1;
      patterns[8959] = 25'b00100010_11111101_00011111_1;
      patterns[8960] = 25'b00100010_11111110_00100000_1;
      patterns[8961] = 25'b00100010_11111111_00100001_1;
      patterns[8962] = 25'b00100011_00000000_00100011_0;
      patterns[8963] = 25'b00100011_00000001_00100100_0;
      patterns[8964] = 25'b00100011_00000010_00100101_0;
      patterns[8965] = 25'b00100011_00000011_00100110_0;
      patterns[8966] = 25'b00100011_00000100_00100111_0;
      patterns[8967] = 25'b00100011_00000101_00101000_0;
      patterns[8968] = 25'b00100011_00000110_00101001_0;
      patterns[8969] = 25'b00100011_00000111_00101010_0;
      patterns[8970] = 25'b00100011_00001000_00101011_0;
      patterns[8971] = 25'b00100011_00001001_00101100_0;
      patterns[8972] = 25'b00100011_00001010_00101101_0;
      patterns[8973] = 25'b00100011_00001011_00101110_0;
      patterns[8974] = 25'b00100011_00001100_00101111_0;
      patterns[8975] = 25'b00100011_00001101_00110000_0;
      patterns[8976] = 25'b00100011_00001110_00110001_0;
      patterns[8977] = 25'b00100011_00001111_00110010_0;
      patterns[8978] = 25'b00100011_00010000_00110011_0;
      patterns[8979] = 25'b00100011_00010001_00110100_0;
      patterns[8980] = 25'b00100011_00010010_00110101_0;
      patterns[8981] = 25'b00100011_00010011_00110110_0;
      patterns[8982] = 25'b00100011_00010100_00110111_0;
      patterns[8983] = 25'b00100011_00010101_00111000_0;
      patterns[8984] = 25'b00100011_00010110_00111001_0;
      patterns[8985] = 25'b00100011_00010111_00111010_0;
      patterns[8986] = 25'b00100011_00011000_00111011_0;
      patterns[8987] = 25'b00100011_00011001_00111100_0;
      patterns[8988] = 25'b00100011_00011010_00111101_0;
      patterns[8989] = 25'b00100011_00011011_00111110_0;
      patterns[8990] = 25'b00100011_00011100_00111111_0;
      patterns[8991] = 25'b00100011_00011101_01000000_0;
      patterns[8992] = 25'b00100011_00011110_01000001_0;
      patterns[8993] = 25'b00100011_00011111_01000010_0;
      patterns[8994] = 25'b00100011_00100000_01000011_0;
      patterns[8995] = 25'b00100011_00100001_01000100_0;
      patterns[8996] = 25'b00100011_00100010_01000101_0;
      patterns[8997] = 25'b00100011_00100011_01000110_0;
      patterns[8998] = 25'b00100011_00100100_01000111_0;
      patterns[8999] = 25'b00100011_00100101_01001000_0;
      patterns[9000] = 25'b00100011_00100110_01001001_0;
      patterns[9001] = 25'b00100011_00100111_01001010_0;
      patterns[9002] = 25'b00100011_00101000_01001011_0;
      patterns[9003] = 25'b00100011_00101001_01001100_0;
      patterns[9004] = 25'b00100011_00101010_01001101_0;
      patterns[9005] = 25'b00100011_00101011_01001110_0;
      patterns[9006] = 25'b00100011_00101100_01001111_0;
      patterns[9007] = 25'b00100011_00101101_01010000_0;
      patterns[9008] = 25'b00100011_00101110_01010001_0;
      patterns[9009] = 25'b00100011_00101111_01010010_0;
      patterns[9010] = 25'b00100011_00110000_01010011_0;
      patterns[9011] = 25'b00100011_00110001_01010100_0;
      patterns[9012] = 25'b00100011_00110010_01010101_0;
      patterns[9013] = 25'b00100011_00110011_01010110_0;
      patterns[9014] = 25'b00100011_00110100_01010111_0;
      patterns[9015] = 25'b00100011_00110101_01011000_0;
      patterns[9016] = 25'b00100011_00110110_01011001_0;
      patterns[9017] = 25'b00100011_00110111_01011010_0;
      patterns[9018] = 25'b00100011_00111000_01011011_0;
      patterns[9019] = 25'b00100011_00111001_01011100_0;
      patterns[9020] = 25'b00100011_00111010_01011101_0;
      patterns[9021] = 25'b00100011_00111011_01011110_0;
      patterns[9022] = 25'b00100011_00111100_01011111_0;
      patterns[9023] = 25'b00100011_00111101_01100000_0;
      patterns[9024] = 25'b00100011_00111110_01100001_0;
      patterns[9025] = 25'b00100011_00111111_01100010_0;
      patterns[9026] = 25'b00100011_01000000_01100011_0;
      patterns[9027] = 25'b00100011_01000001_01100100_0;
      patterns[9028] = 25'b00100011_01000010_01100101_0;
      patterns[9029] = 25'b00100011_01000011_01100110_0;
      patterns[9030] = 25'b00100011_01000100_01100111_0;
      patterns[9031] = 25'b00100011_01000101_01101000_0;
      patterns[9032] = 25'b00100011_01000110_01101001_0;
      patterns[9033] = 25'b00100011_01000111_01101010_0;
      patterns[9034] = 25'b00100011_01001000_01101011_0;
      patterns[9035] = 25'b00100011_01001001_01101100_0;
      patterns[9036] = 25'b00100011_01001010_01101101_0;
      patterns[9037] = 25'b00100011_01001011_01101110_0;
      patterns[9038] = 25'b00100011_01001100_01101111_0;
      patterns[9039] = 25'b00100011_01001101_01110000_0;
      patterns[9040] = 25'b00100011_01001110_01110001_0;
      patterns[9041] = 25'b00100011_01001111_01110010_0;
      patterns[9042] = 25'b00100011_01010000_01110011_0;
      patterns[9043] = 25'b00100011_01010001_01110100_0;
      patterns[9044] = 25'b00100011_01010010_01110101_0;
      patterns[9045] = 25'b00100011_01010011_01110110_0;
      patterns[9046] = 25'b00100011_01010100_01110111_0;
      patterns[9047] = 25'b00100011_01010101_01111000_0;
      patterns[9048] = 25'b00100011_01010110_01111001_0;
      patterns[9049] = 25'b00100011_01010111_01111010_0;
      patterns[9050] = 25'b00100011_01011000_01111011_0;
      patterns[9051] = 25'b00100011_01011001_01111100_0;
      patterns[9052] = 25'b00100011_01011010_01111101_0;
      patterns[9053] = 25'b00100011_01011011_01111110_0;
      patterns[9054] = 25'b00100011_01011100_01111111_0;
      patterns[9055] = 25'b00100011_01011101_10000000_0;
      patterns[9056] = 25'b00100011_01011110_10000001_0;
      patterns[9057] = 25'b00100011_01011111_10000010_0;
      patterns[9058] = 25'b00100011_01100000_10000011_0;
      patterns[9059] = 25'b00100011_01100001_10000100_0;
      patterns[9060] = 25'b00100011_01100010_10000101_0;
      patterns[9061] = 25'b00100011_01100011_10000110_0;
      patterns[9062] = 25'b00100011_01100100_10000111_0;
      patterns[9063] = 25'b00100011_01100101_10001000_0;
      patterns[9064] = 25'b00100011_01100110_10001001_0;
      patterns[9065] = 25'b00100011_01100111_10001010_0;
      patterns[9066] = 25'b00100011_01101000_10001011_0;
      patterns[9067] = 25'b00100011_01101001_10001100_0;
      patterns[9068] = 25'b00100011_01101010_10001101_0;
      patterns[9069] = 25'b00100011_01101011_10001110_0;
      patterns[9070] = 25'b00100011_01101100_10001111_0;
      patterns[9071] = 25'b00100011_01101101_10010000_0;
      patterns[9072] = 25'b00100011_01101110_10010001_0;
      patterns[9073] = 25'b00100011_01101111_10010010_0;
      patterns[9074] = 25'b00100011_01110000_10010011_0;
      patterns[9075] = 25'b00100011_01110001_10010100_0;
      patterns[9076] = 25'b00100011_01110010_10010101_0;
      patterns[9077] = 25'b00100011_01110011_10010110_0;
      patterns[9078] = 25'b00100011_01110100_10010111_0;
      patterns[9079] = 25'b00100011_01110101_10011000_0;
      patterns[9080] = 25'b00100011_01110110_10011001_0;
      patterns[9081] = 25'b00100011_01110111_10011010_0;
      patterns[9082] = 25'b00100011_01111000_10011011_0;
      patterns[9083] = 25'b00100011_01111001_10011100_0;
      patterns[9084] = 25'b00100011_01111010_10011101_0;
      patterns[9085] = 25'b00100011_01111011_10011110_0;
      patterns[9086] = 25'b00100011_01111100_10011111_0;
      patterns[9087] = 25'b00100011_01111101_10100000_0;
      patterns[9088] = 25'b00100011_01111110_10100001_0;
      patterns[9089] = 25'b00100011_01111111_10100010_0;
      patterns[9090] = 25'b00100011_10000000_10100011_0;
      patterns[9091] = 25'b00100011_10000001_10100100_0;
      patterns[9092] = 25'b00100011_10000010_10100101_0;
      patterns[9093] = 25'b00100011_10000011_10100110_0;
      patterns[9094] = 25'b00100011_10000100_10100111_0;
      patterns[9095] = 25'b00100011_10000101_10101000_0;
      patterns[9096] = 25'b00100011_10000110_10101001_0;
      patterns[9097] = 25'b00100011_10000111_10101010_0;
      patterns[9098] = 25'b00100011_10001000_10101011_0;
      patterns[9099] = 25'b00100011_10001001_10101100_0;
      patterns[9100] = 25'b00100011_10001010_10101101_0;
      patterns[9101] = 25'b00100011_10001011_10101110_0;
      patterns[9102] = 25'b00100011_10001100_10101111_0;
      patterns[9103] = 25'b00100011_10001101_10110000_0;
      patterns[9104] = 25'b00100011_10001110_10110001_0;
      patterns[9105] = 25'b00100011_10001111_10110010_0;
      patterns[9106] = 25'b00100011_10010000_10110011_0;
      patterns[9107] = 25'b00100011_10010001_10110100_0;
      patterns[9108] = 25'b00100011_10010010_10110101_0;
      patterns[9109] = 25'b00100011_10010011_10110110_0;
      patterns[9110] = 25'b00100011_10010100_10110111_0;
      patterns[9111] = 25'b00100011_10010101_10111000_0;
      patterns[9112] = 25'b00100011_10010110_10111001_0;
      patterns[9113] = 25'b00100011_10010111_10111010_0;
      patterns[9114] = 25'b00100011_10011000_10111011_0;
      patterns[9115] = 25'b00100011_10011001_10111100_0;
      patterns[9116] = 25'b00100011_10011010_10111101_0;
      patterns[9117] = 25'b00100011_10011011_10111110_0;
      patterns[9118] = 25'b00100011_10011100_10111111_0;
      patterns[9119] = 25'b00100011_10011101_11000000_0;
      patterns[9120] = 25'b00100011_10011110_11000001_0;
      patterns[9121] = 25'b00100011_10011111_11000010_0;
      patterns[9122] = 25'b00100011_10100000_11000011_0;
      patterns[9123] = 25'b00100011_10100001_11000100_0;
      patterns[9124] = 25'b00100011_10100010_11000101_0;
      patterns[9125] = 25'b00100011_10100011_11000110_0;
      patterns[9126] = 25'b00100011_10100100_11000111_0;
      patterns[9127] = 25'b00100011_10100101_11001000_0;
      patterns[9128] = 25'b00100011_10100110_11001001_0;
      patterns[9129] = 25'b00100011_10100111_11001010_0;
      patterns[9130] = 25'b00100011_10101000_11001011_0;
      patterns[9131] = 25'b00100011_10101001_11001100_0;
      patterns[9132] = 25'b00100011_10101010_11001101_0;
      patterns[9133] = 25'b00100011_10101011_11001110_0;
      patterns[9134] = 25'b00100011_10101100_11001111_0;
      patterns[9135] = 25'b00100011_10101101_11010000_0;
      patterns[9136] = 25'b00100011_10101110_11010001_0;
      patterns[9137] = 25'b00100011_10101111_11010010_0;
      patterns[9138] = 25'b00100011_10110000_11010011_0;
      patterns[9139] = 25'b00100011_10110001_11010100_0;
      patterns[9140] = 25'b00100011_10110010_11010101_0;
      patterns[9141] = 25'b00100011_10110011_11010110_0;
      patterns[9142] = 25'b00100011_10110100_11010111_0;
      patterns[9143] = 25'b00100011_10110101_11011000_0;
      patterns[9144] = 25'b00100011_10110110_11011001_0;
      patterns[9145] = 25'b00100011_10110111_11011010_0;
      patterns[9146] = 25'b00100011_10111000_11011011_0;
      patterns[9147] = 25'b00100011_10111001_11011100_0;
      patterns[9148] = 25'b00100011_10111010_11011101_0;
      patterns[9149] = 25'b00100011_10111011_11011110_0;
      patterns[9150] = 25'b00100011_10111100_11011111_0;
      patterns[9151] = 25'b00100011_10111101_11100000_0;
      patterns[9152] = 25'b00100011_10111110_11100001_0;
      patterns[9153] = 25'b00100011_10111111_11100010_0;
      patterns[9154] = 25'b00100011_11000000_11100011_0;
      patterns[9155] = 25'b00100011_11000001_11100100_0;
      patterns[9156] = 25'b00100011_11000010_11100101_0;
      patterns[9157] = 25'b00100011_11000011_11100110_0;
      patterns[9158] = 25'b00100011_11000100_11100111_0;
      patterns[9159] = 25'b00100011_11000101_11101000_0;
      patterns[9160] = 25'b00100011_11000110_11101001_0;
      patterns[9161] = 25'b00100011_11000111_11101010_0;
      patterns[9162] = 25'b00100011_11001000_11101011_0;
      patterns[9163] = 25'b00100011_11001001_11101100_0;
      patterns[9164] = 25'b00100011_11001010_11101101_0;
      patterns[9165] = 25'b00100011_11001011_11101110_0;
      patterns[9166] = 25'b00100011_11001100_11101111_0;
      patterns[9167] = 25'b00100011_11001101_11110000_0;
      patterns[9168] = 25'b00100011_11001110_11110001_0;
      patterns[9169] = 25'b00100011_11001111_11110010_0;
      patterns[9170] = 25'b00100011_11010000_11110011_0;
      patterns[9171] = 25'b00100011_11010001_11110100_0;
      patterns[9172] = 25'b00100011_11010010_11110101_0;
      patterns[9173] = 25'b00100011_11010011_11110110_0;
      patterns[9174] = 25'b00100011_11010100_11110111_0;
      patterns[9175] = 25'b00100011_11010101_11111000_0;
      patterns[9176] = 25'b00100011_11010110_11111001_0;
      patterns[9177] = 25'b00100011_11010111_11111010_0;
      patterns[9178] = 25'b00100011_11011000_11111011_0;
      patterns[9179] = 25'b00100011_11011001_11111100_0;
      patterns[9180] = 25'b00100011_11011010_11111101_0;
      patterns[9181] = 25'b00100011_11011011_11111110_0;
      patterns[9182] = 25'b00100011_11011100_11111111_0;
      patterns[9183] = 25'b00100011_11011101_00000000_1;
      patterns[9184] = 25'b00100011_11011110_00000001_1;
      patterns[9185] = 25'b00100011_11011111_00000010_1;
      patterns[9186] = 25'b00100011_11100000_00000011_1;
      patterns[9187] = 25'b00100011_11100001_00000100_1;
      patterns[9188] = 25'b00100011_11100010_00000101_1;
      patterns[9189] = 25'b00100011_11100011_00000110_1;
      patterns[9190] = 25'b00100011_11100100_00000111_1;
      patterns[9191] = 25'b00100011_11100101_00001000_1;
      patterns[9192] = 25'b00100011_11100110_00001001_1;
      patterns[9193] = 25'b00100011_11100111_00001010_1;
      patterns[9194] = 25'b00100011_11101000_00001011_1;
      patterns[9195] = 25'b00100011_11101001_00001100_1;
      patterns[9196] = 25'b00100011_11101010_00001101_1;
      patterns[9197] = 25'b00100011_11101011_00001110_1;
      patterns[9198] = 25'b00100011_11101100_00001111_1;
      patterns[9199] = 25'b00100011_11101101_00010000_1;
      patterns[9200] = 25'b00100011_11101110_00010001_1;
      patterns[9201] = 25'b00100011_11101111_00010010_1;
      patterns[9202] = 25'b00100011_11110000_00010011_1;
      patterns[9203] = 25'b00100011_11110001_00010100_1;
      patterns[9204] = 25'b00100011_11110010_00010101_1;
      patterns[9205] = 25'b00100011_11110011_00010110_1;
      patterns[9206] = 25'b00100011_11110100_00010111_1;
      patterns[9207] = 25'b00100011_11110101_00011000_1;
      patterns[9208] = 25'b00100011_11110110_00011001_1;
      patterns[9209] = 25'b00100011_11110111_00011010_1;
      patterns[9210] = 25'b00100011_11111000_00011011_1;
      patterns[9211] = 25'b00100011_11111001_00011100_1;
      patterns[9212] = 25'b00100011_11111010_00011101_1;
      patterns[9213] = 25'b00100011_11111011_00011110_1;
      patterns[9214] = 25'b00100011_11111100_00011111_1;
      patterns[9215] = 25'b00100011_11111101_00100000_1;
      patterns[9216] = 25'b00100011_11111110_00100001_1;
      patterns[9217] = 25'b00100011_11111111_00100010_1;
      patterns[9218] = 25'b00100100_00000000_00100100_0;
      patterns[9219] = 25'b00100100_00000001_00100101_0;
      patterns[9220] = 25'b00100100_00000010_00100110_0;
      patterns[9221] = 25'b00100100_00000011_00100111_0;
      patterns[9222] = 25'b00100100_00000100_00101000_0;
      patterns[9223] = 25'b00100100_00000101_00101001_0;
      patterns[9224] = 25'b00100100_00000110_00101010_0;
      patterns[9225] = 25'b00100100_00000111_00101011_0;
      patterns[9226] = 25'b00100100_00001000_00101100_0;
      patterns[9227] = 25'b00100100_00001001_00101101_0;
      patterns[9228] = 25'b00100100_00001010_00101110_0;
      patterns[9229] = 25'b00100100_00001011_00101111_0;
      patterns[9230] = 25'b00100100_00001100_00110000_0;
      patterns[9231] = 25'b00100100_00001101_00110001_0;
      patterns[9232] = 25'b00100100_00001110_00110010_0;
      patterns[9233] = 25'b00100100_00001111_00110011_0;
      patterns[9234] = 25'b00100100_00010000_00110100_0;
      patterns[9235] = 25'b00100100_00010001_00110101_0;
      patterns[9236] = 25'b00100100_00010010_00110110_0;
      patterns[9237] = 25'b00100100_00010011_00110111_0;
      patterns[9238] = 25'b00100100_00010100_00111000_0;
      patterns[9239] = 25'b00100100_00010101_00111001_0;
      patterns[9240] = 25'b00100100_00010110_00111010_0;
      patterns[9241] = 25'b00100100_00010111_00111011_0;
      patterns[9242] = 25'b00100100_00011000_00111100_0;
      patterns[9243] = 25'b00100100_00011001_00111101_0;
      patterns[9244] = 25'b00100100_00011010_00111110_0;
      patterns[9245] = 25'b00100100_00011011_00111111_0;
      patterns[9246] = 25'b00100100_00011100_01000000_0;
      patterns[9247] = 25'b00100100_00011101_01000001_0;
      patterns[9248] = 25'b00100100_00011110_01000010_0;
      patterns[9249] = 25'b00100100_00011111_01000011_0;
      patterns[9250] = 25'b00100100_00100000_01000100_0;
      patterns[9251] = 25'b00100100_00100001_01000101_0;
      patterns[9252] = 25'b00100100_00100010_01000110_0;
      patterns[9253] = 25'b00100100_00100011_01000111_0;
      patterns[9254] = 25'b00100100_00100100_01001000_0;
      patterns[9255] = 25'b00100100_00100101_01001001_0;
      patterns[9256] = 25'b00100100_00100110_01001010_0;
      patterns[9257] = 25'b00100100_00100111_01001011_0;
      patterns[9258] = 25'b00100100_00101000_01001100_0;
      patterns[9259] = 25'b00100100_00101001_01001101_0;
      patterns[9260] = 25'b00100100_00101010_01001110_0;
      patterns[9261] = 25'b00100100_00101011_01001111_0;
      patterns[9262] = 25'b00100100_00101100_01010000_0;
      patterns[9263] = 25'b00100100_00101101_01010001_0;
      patterns[9264] = 25'b00100100_00101110_01010010_0;
      patterns[9265] = 25'b00100100_00101111_01010011_0;
      patterns[9266] = 25'b00100100_00110000_01010100_0;
      patterns[9267] = 25'b00100100_00110001_01010101_0;
      patterns[9268] = 25'b00100100_00110010_01010110_0;
      patterns[9269] = 25'b00100100_00110011_01010111_0;
      patterns[9270] = 25'b00100100_00110100_01011000_0;
      patterns[9271] = 25'b00100100_00110101_01011001_0;
      patterns[9272] = 25'b00100100_00110110_01011010_0;
      patterns[9273] = 25'b00100100_00110111_01011011_0;
      patterns[9274] = 25'b00100100_00111000_01011100_0;
      patterns[9275] = 25'b00100100_00111001_01011101_0;
      patterns[9276] = 25'b00100100_00111010_01011110_0;
      patterns[9277] = 25'b00100100_00111011_01011111_0;
      patterns[9278] = 25'b00100100_00111100_01100000_0;
      patterns[9279] = 25'b00100100_00111101_01100001_0;
      patterns[9280] = 25'b00100100_00111110_01100010_0;
      patterns[9281] = 25'b00100100_00111111_01100011_0;
      patterns[9282] = 25'b00100100_01000000_01100100_0;
      patterns[9283] = 25'b00100100_01000001_01100101_0;
      patterns[9284] = 25'b00100100_01000010_01100110_0;
      patterns[9285] = 25'b00100100_01000011_01100111_0;
      patterns[9286] = 25'b00100100_01000100_01101000_0;
      patterns[9287] = 25'b00100100_01000101_01101001_0;
      patterns[9288] = 25'b00100100_01000110_01101010_0;
      patterns[9289] = 25'b00100100_01000111_01101011_0;
      patterns[9290] = 25'b00100100_01001000_01101100_0;
      patterns[9291] = 25'b00100100_01001001_01101101_0;
      patterns[9292] = 25'b00100100_01001010_01101110_0;
      patterns[9293] = 25'b00100100_01001011_01101111_0;
      patterns[9294] = 25'b00100100_01001100_01110000_0;
      patterns[9295] = 25'b00100100_01001101_01110001_0;
      patterns[9296] = 25'b00100100_01001110_01110010_0;
      patterns[9297] = 25'b00100100_01001111_01110011_0;
      patterns[9298] = 25'b00100100_01010000_01110100_0;
      patterns[9299] = 25'b00100100_01010001_01110101_0;
      patterns[9300] = 25'b00100100_01010010_01110110_0;
      patterns[9301] = 25'b00100100_01010011_01110111_0;
      patterns[9302] = 25'b00100100_01010100_01111000_0;
      patterns[9303] = 25'b00100100_01010101_01111001_0;
      patterns[9304] = 25'b00100100_01010110_01111010_0;
      patterns[9305] = 25'b00100100_01010111_01111011_0;
      patterns[9306] = 25'b00100100_01011000_01111100_0;
      patterns[9307] = 25'b00100100_01011001_01111101_0;
      patterns[9308] = 25'b00100100_01011010_01111110_0;
      patterns[9309] = 25'b00100100_01011011_01111111_0;
      patterns[9310] = 25'b00100100_01011100_10000000_0;
      patterns[9311] = 25'b00100100_01011101_10000001_0;
      patterns[9312] = 25'b00100100_01011110_10000010_0;
      patterns[9313] = 25'b00100100_01011111_10000011_0;
      patterns[9314] = 25'b00100100_01100000_10000100_0;
      patterns[9315] = 25'b00100100_01100001_10000101_0;
      patterns[9316] = 25'b00100100_01100010_10000110_0;
      patterns[9317] = 25'b00100100_01100011_10000111_0;
      patterns[9318] = 25'b00100100_01100100_10001000_0;
      patterns[9319] = 25'b00100100_01100101_10001001_0;
      patterns[9320] = 25'b00100100_01100110_10001010_0;
      patterns[9321] = 25'b00100100_01100111_10001011_0;
      patterns[9322] = 25'b00100100_01101000_10001100_0;
      patterns[9323] = 25'b00100100_01101001_10001101_0;
      patterns[9324] = 25'b00100100_01101010_10001110_0;
      patterns[9325] = 25'b00100100_01101011_10001111_0;
      patterns[9326] = 25'b00100100_01101100_10010000_0;
      patterns[9327] = 25'b00100100_01101101_10010001_0;
      patterns[9328] = 25'b00100100_01101110_10010010_0;
      patterns[9329] = 25'b00100100_01101111_10010011_0;
      patterns[9330] = 25'b00100100_01110000_10010100_0;
      patterns[9331] = 25'b00100100_01110001_10010101_0;
      patterns[9332] = 25'b00100100_01110010_10010110_0;
      patterns[9333] = 25'b00100100_01110011_10010111_0;
      patterns[9334] = 25'b00100100_01110100_10011000_0;
      patterns[9335] = 25'b00100100_01110101_10011001_0;
      patterns[9336] = 25'b00100100_01110110_10011010_0;
      patterns[9337] = 25'b00100100_01110111_10011011_0;
      patterns[9338] = 25'b00100100_01111000_10011100_0;
      patterns[9339] = 25'b00100100_01111001_10011101_0;
      patterns[9340] = 25'b00100100_01111010_10011110_0;
      patterns[9341] = 25'b00100100_01111011_10011111_0;
      patterns[9342] = 25'b00100100_01111100_10100000_0;
      patterns[9343] = 25'b00100100_01111101_10100001_0;
      patterns[9344] = 25'b00100100_01111110_10100010_0;
      patterns[9345] = 25'b00100100_01111111_10100011_0;
      patterns[9346] = 25'b00100100_10000000_10100100_0;
      patterns[9347] = 25'b00100100_10000001_10100101_0;
      patterns[9348] = 25'b00100100_10000010_10100110_0;
      patterns[9349] = 25'b00100100_10000011_10100111_0;
      patterns[9350] = 25'b00100100_10000100_10101000_0;
      patterns[9351] = 25'b00100100_10000101_10101001_0;
      patterns[9352] = 25'b00100100_10000110_10101010_0;
      patterns[9353] = 25'b00100100_10000111_10101011_0;
      patterns[9354] = 25'b00100100_10001000_10101100_0;
      patterns[9355] = 25'b00100100_10001001_10101101_0;
      patterns[9356] = 25'b00100100_10001010_10101110_0;
      patterns[9357] = 25'b00100100_10001011_10101111_0;
      patterns[9358] = 25'b00100100_10001100_10110000_0;
      patterns[9359] = 25'b00100100_10001101_10110001_0;
      patterns[9360] = 25'b00100100_10001110_10110010_0;
      patterns[9361] = 25'b00100100_10001111_10110011_0;
      patterns[9362] = 25'b00100100_10010000_10110100_0;
      patterns[9363] = 25'b00100100_10010001_10110101_0;
      patterns[9364] = 25'b00100100_10010010_10110110_0;
      patterns[9365] = 25'b00100100_10010011_10110111_0;
      patterns[9366] = 25'b00100100_10010100_10111000_0;
      patterns[9367] = 25'b00100100_10010101_10111001_0;
      patterns[9368] = 25'b00100100_10010110_10111010_0;
      patterns[9369] = 25'b00100100_10010111_10111011_0;
      patterns[9370] = 25'b00100100_10011000_10111100_0;
      patterns[9371] = 25'b00100100_10011001_10111101_0;
      patterns[9372] = 25'b00100100_10011010_10111110_0;
      patterns[9373] = 25'b00100100_10011011_10111111_0;
      patterns[9374] = 25'b00100100_10011100_11000000_0;
      patterns[9375] = 25'b00100100_10011101_11000001_0;
      patterns[9376] = 25'b00100100_10011110_11000010_0;
      patterns[9377] = 25'b00100100_10011111_11000011_0;
      patterns[9378] = 25'b00100100_10100000_11000100_0;
      patterns[9379] = 25'b00100100_10100001_11000101_0;
      patterns[9380] = 25'b00100100_10100010_11000110_0;
      patterns[9381] = 25'b00100100_10100011_11000111_0;
      patterns[9382] = 25'b00100100_10100100_11001000_0;
      patterns[9383] = 25'b00100100_10100101_11001001_0;
      patterns[9384] = 25'b00100100_10100110_11001010_0;
      patterns[9385] = 25'b00100100_10100111_11001011_0;
      patterns[9386] = 25'b00100100_10101000_11001100_0;
      patterns[9387] = 25'b00100100_10101001_11001101_0;
      patterns[9388] = 25'b00100100_10101010_11001110_0;
      patterns[9389] = 25'b00100100_10101011_11001111_0;
      patterns[9390] = 25'b00100100_10101100_11010000_0;
      patterns[9391] = 25'b00100100_10101101_11010001_0;
      patterns[9392] = 25'b00100100_10101110_11010010_0;
      patterns[9393] = 25'b00100100_10101111_11010011_0;
      patterns[9394] = 25'b00100100_10110000_11010100_0;
      patterns[9395] = 25'b00100100_10110001_11010101_0;
      patterns[9396] = 25'b00100100_10110010_11010110_0;
      patterns[9397] = 25'b00100100_10110011_11010111_0;
      patterns[9398] = 25'b00100100_10110100_11011000_0;
      patterns[9399] = 25'b00100100_10110101_11011001_0;
      patterns[9400] = 25'b00100100_10110110_11011010_0;
      patterns[9401] = 25'b00100100_10110111_11011011_0;
      patterns[9402] = 25'b00100100_10111000_11011100_0;
      patterns[9403] = 25'b00100100_10111001_11011101_0;
      patterns[9404] = 25'b00100100_10111010_11011110_0;
      patterns[9405] = 25'b00100100_10111011_11011111_0;
      patterns[9406] = 25'b00100100_10111100_11100000_0;
      patterns[9407] = 25'b00100100_10111101_11100001_0;
      patterns[9408] = 25'b00100100_10111110_11100010_0;
      patterns[9409] = 25'b00100100_10111111_11100011_0;
      patterns[9410] = 25'b00100100_11000000_11100100_0;
      patterns[9411] = 25'b00100100_11000001_11100101_0;
      patterns[9412] = 25'b00100100_11000010_11100110_0;
      patterns[9413] = 25'b00100100_11000011_11100111_0;
      patterns[9414] = 25'b00100100_11000100_11101000_0;
      patterns[9415] = 25'b00100100_11000101_11101001_0;
      patterns[9416] = 25'b00100100_11000110_11101010_0;
      patterns[9417] = 25'b00100100_11000111_11101011_0;
      patterns[9418] = 25'b00100100_11001000_11101100_0;
      patterns[9419] = 25'b00100100_11001001_11101101_0;
      patterns[9420] = 25'b00100100_11001010_11101110_0;
      patterns[9421] = 25'b00100100_11001011_11101111_0;
      patterns[9422] = 25'b00100100_11001100_11110000_0;
      patterns[9423] = 25'b00100100_11001101_11110001_0;
      patterns[9424] = 25'b00100100_11001110_11110010_0;
      patterns[9425] = 25'b00100100_11001111_11110011_0;
      patterns[9426] = 25'b00100100_11010000_11110100_0;
      patterns[9427] = 25'b00100100_11010001_11110101_0;
      patterns[9428] = 25'b00100100_11010010_11110110_0;
      patterns[9429] = 25'b00100100_11010011_11110111_0;
      patterns[9430] = 25'b00100100_11010100_11111000_0;
      patterns[9431] = 25'b00100100_11010101_11111001_0;
      patterns[9432] = 25'b00100100_11010110_11111010_0;
      patterns[9433] = 25'b00100100_11010111_11111011_0;
      patterns[9434] = 25'b00100100_11011000_11111100_0;
      patterns[9435] = 25'b00100100_11011001_11111101_0;
      patterns[9436] = 25'b00100100_11011010_11111110_0;
      patterns[9437] = 25'b00100100_11011011_11111111_0;
      patterns[9438] = 25'b00100100_11011100_00000000_1;
      patterns[9439] = 25'b00100100_11011101_00000001_1;
      patterns[9440] = 25'b00100100_11011110_00000010_1;
      patterns[9441] = 25'b00100100_11011111_00000011_1;
      patterns[9442] = 25'b00100100_11100000_00000100_1;
      patterns[9443] = 25'b00100100_11100001_00000101_1;
      patterns[9444] = 25'b00100100_11100010_00000110_1;
      patterns[9445] = 25'b00100100_11100011_00000111_1;
      patterns[9446] = 25'b00100100_11100100_00001000_1;
      patterns[9447] = 25'b00100100_11100101_00001001_1;
      patterns[9448] = 25'b00100100_11100110_00001010_1;
      patterns[9449] = 25'b00100100_11100111_00001011_1;
      patterns[9450] = 25'b00100100_11101000_00001100_1;
      patterns[9451] = 25'b00100100_11101001_00001101_1;
      patterns[9452] = 25'b00100100_11101010_00001110_1;
      patterns[9453] = 25'b00100100_11101011_00001111_1;
      patterns[9454] = 25'b00100100_11101100_00010000_1;
      patterns[9455] = 25'b00100100_11101101_00010001_1;
      patterns[9456] = 25'b00100100_11101110_00010010_1;
      patterns[9457] = 25'b00100100_11101111_00010011_1;
      patterns[9458] = 25'b00100100_11110000_00010100_1;
      patterns[9459] = 25'b00100100_11110001_00010101_1;
      patterns[9460] = 25'b00100100_11110010_00010110_1;
      patterns[9461] = 25'b00100100_11110011_00010111_1;
      patterns[9462] = 25'b00100100_11110100_00011000_1;
      patterns[9463] = 25'b00100100_11110101_00011001_1;
      patterns[9464] = 25'b00100100_11110110_00011010_1;
      patterns[9465] = 25'b00100100_11110111_00011011_1;
      patterns[9466] = 25'b00100100_11111000_00011100_1;
      patterns[9467] = 25'b00100100_11111001_00011101_1;
      patterns[9468] = 25'b00100100_11111010_00011110_1;
      patterns[9469] = 25'b00100100_11111011_00011111_1;
      patterns[9470] = 25'b00100100_11111100_00100000_1;
      patterns[9471] = 25'b00100100_11111101_00100001_1;
      patterns[9472] = 25'b00100100_11111110_00100010_1;
      patterns[9473] = 25'b00100100_11111111_00100011_1;
      patterns[9474] = 25'b00100101_00000000_00100101_0;
      patterns[9475] = 25'b00100101_00000001_00100110_0;
      patterns[9476] = 25'b00100101_00000010_00100111_0;
      patterns[9477] = 25'b00100101_00000011_00101000_0;
      patterns[9478] = 25'b00100101_00000100_00101001_0;
      patterns[9479] = 25'b00100101_00000101_00101010_0;
      patterns[9480] = 25'b00100101_00000110_00101011_0;
      patterns[9481] = 25'b00100101_00000111_00101100_0;
      patterns[9482] = 25'b00100101_00001000_00101101_0;
      patterns[9483] = 25'b00100101_00001001_00101110_0;
      patterns[9484] = 25'b00100101_00001010_00101111_0;
      patterns[9485] = 25'b00100101_00001011_00110000_0;
      patterns[9486] = 25'b00100101_00001100_00110001_0;
      patterns[9487] = 25'b00100101_00001101_00110010_0;
      patterns[9488] = 25'b00100101_00001110_00110011_0;
      patterns[9489] = 25'b00100101_00001111_00110100_0;
      patterns[9490] = 25'b00100101_00010000_00110101_0;
      patterns[9491] = 25'b00100101_00010001_00110110_0;
      patterns[9492] = 25'b00100101_00010010_00110111_0;
      patterns[9493] = 25'b00100101_00010011_00111000_0;
      patterns[9494] = 25'b00100101_00010100_00111001_0;
      patterns[9495] = 25'b00100101_00010101_00111010_0;
      patterns[9496] = 25'b00100101_00010110_00111011_0;
      patterns[9497] = 25'b00100101_00010111_00111100_0;
      patterns[9498] = 25'b00100101_00011000_00111101_0;
      patterns[9499] = 25'b00100101_00011001_00111110_0;
      patterns[9500] = 25'b00100101_00011010_00111111_0;
      patterns[9501] = 25'b00100101_00011011_01000000_0;
      patterns[9502] = 25'b00100101_00011100_01000001_0;
      patterns[9503] = 25'b00100101_00011101_01000010_0;
      patterns[9504] = 25'b00100101_00011110_01000011_0;
      patterns[9505] = 25'b00100101_00011111_01000100_0;
      patterns[9506] = 25'b00100101_00100000_01000101_0;
      patterns[9507] = 25'b00100101_00100001_01000110_0;
      patterns[9508] = 25'b00100101_00100010_01000111_0;
      patterns[9509] = 25'b00100101_00100011_01001000_0;
      patterns[9510] = 25'b00100101_00100100_01001001_0;
      patterns[9511] = 25'b00100101_00100101_01001010_0;
      patterns[9512] = 25'b00100101_00100110_01001011_0;
      patterns[9513] = 25'b00100101_00100111_01001100_0;
      patterns[9514] = 25'b00100101_00101000_01001101_0;
      patterns[9515] = 25'b00100101_00101001_01001110_0;
      patterns[9516] = 25'b00100101_00101010_01001111_0;
      patterns[9517] = 25'b00100101_00101011_01010000_0;
      patterns[9518] = 25'b00100101_00101100_01010001_0;
      patterns[9519] = 25'b00100101_00101101_01010010_0;
      patterns[9520] = 25'b00100101_00101110_01010011_0;
      patterns[9521] = 25'b00100101_00101111_01010100_0;
      patterns[9522] = 25'b00100101_00110000_01010101_0;
      patterns[9523] = 25'b00100101_00110001_01010110_0;
      patterns[9524] = 25'b00100101_00110010_01010111_0;
      patterns[9525] = 25'b00100101_00110011_01011000_0;
      patterns[9526] = 25'b00100101_00110100_01011001_0;
      patterns[9527] = 25'b00100101_00110101_01011010_0;
      patterns[9528] = 25'b00100101_00110110_01011011_0;
      patterns[9529] = 25'b00100101_00110111_01011100_0;
      patterns[9530] = 25'b00100101_00111000_01011101_0;
      patterns[9531] = 25'b00100101_00111001_01011110_0;
      patterns[9532] = 25'b00100101_00111010_01011111_0;
      patterns[9533] = 25'b00100101_00111011_01100000_0;
      patterns[9534] = 25'b00100101_00111100_01100001_0;
      patterns[9535] = 25'b00100101_00111101_01100010_0;
      patterns[9536] = 25'b00100101_00111110_01100011_0;
      patterns[9537] = 25'b00100101_00111111_01100100_0;
      patterns[9538] = 25'b00100101_01000000_01100101_0;
      patterns[9539] = 25'b00100101_01000001_01100110_0;
      patterns[9540] = 25'b00100101_01000010_01100111_0;
      patterns[9541] = 25'b00100101_01000011_01101000_0;
      patterns[9542] = 25'b00100101_01000100_01101001_0;
      patterns[9543] = 25'b00100101_01000101_01101010_0;
      patterns[9544] = 25'b00100101_01000110_01101011_0;
      patterns[9545] = 25'b00100101_01000111_01101100_0;
      patterns[9546] = 25'b00100101_01001000_01101101_0;
      patterns[9547] = 25'b00100101_01001001_01101110_0;
      patterns[9548] = 25'b00100101_01001010_01101111_0;
      patterns[9549] = 25'b00100101_01001011_01110000_0;
      patterns[9550] = 25'b00100101_01001100_01110001_0;
      patterns[9551] = 25'b00100101_01001101_01110010_0;
      patterns[9552] = 25'b00100101_01001110_01110011_0;
      patterns[9553] = 25'b00100101_01001111_01110100_0;
      patterns[9554] = 25'b00100101_01010000_01110101_0;
      patterns[9555] = 25'b00100101_01010001_01110110_0;
      patterns[9556] = 25'b00100101_01010010_01110111_0;
      patterns[9557] = 25'b00100101_01010011_01111000_0;
      patterns[9558] = 25'b00100101_01010100_01111001_0;
      patterns[9559] = 25'b00100101_01010101_01111010_0;
      patterns[9560] = 25'b00100101_01010110_01111011_0;
      patterns[9561] = 25'b00100101_01010111_01111100_0;
      patterns[9562] = 25'b00100101_01011000_01111101_0;
      patterns[9563] = 25'b00100101_01011001_01111110_0;
      patterns[9564] = 25'b00100101_01011010_01111111_0;
      patterns[9565] = 25'b00100101_01011011_10000000_0;
      patterns[9566] = 25'b00100101_01011100_10000001_0;
      patterns[9567] = 25'b00100101_01011101_10000010_0;
      patterns[9568] = 25'b00100101_01011110_10000011_0;
      patterns[9569] = 25'b00100101_01011111_10000100_0;
      patterns[9570] = 25'b00100101_01100000_10000101_0;
      patterns[9571] = 25'b00100101_01100001_10000110_0;
      patterns[9572] = 25'b00100101_01100010_10000111_0;
      patterns[9573] = 25'b00100101_01100011_10001000_0;
      patterns[9574] = 25'b00100101_01100100_10001001_0;
      patterns[9575] = 25'b00100101_01100101_10001010_0;
      patterns[9576] = 25'b00100101_01100110_10001011_0;
      patterns[9577] = 25'b00100101_01100111_10001100_0;
      patterns[9578] = 25'b00100101_01101000_10001101_0;
      patterns[9579] = 25'b00100101_01101001_10001110_0;
      patterns[9580] = 25'b00100101_01101010_10001111_0;
      patterns[9581] = 25'b00100101_01101011_10010000_0;
      patterns[9582] = 25'b00100101_01101100_10010001_0;
      patterns[9583] = 25'b00100101_01101101_10010010_0;
      patterns[9584] = 25'b00100101_01101110_10010011_0;
      patterns[9585] = 25'b00100101_01101111_10010100_0;
      patterns[9586] = 25'b00100101_01110000_10010101_0;
      patterns[9587] = 25'b00100101_01110001_10010110_0;
      patterns[9588] = 25'b00100101_01110010_10010111_0;
      patterns[9589] = 25'b00100101_01110011_10011000_0;
      patterns[9590] = 25'b00100101_01110100_10011001_0;
      patterns[9591] = 25'b00100101_01110101_10011010_0;
      patterns[9592] = 25'b00100101_01110110_10011011_0;
      patterns[9593] = 25'b00100101_01110111_10011100_0;
      patterns[9594] = 25'b00100101_01111000_10011101_0;
      patterns[9595] = 25'b00100101_01111001_10011110_0;
      patterns[9596] = 25'b00100101_01111010_10011111_0;
      patterns[9597] = 25'b00100101_01111011_10100000_0;
      patterns[9598] = 25'b00100101_01111100_10100001_0;
      patterns[9599] = 25'b00100101_01111101_10100010_0;
      patterns[9600] = 25'b00100101_01111110_10100011_0;
      patterns[9601] = 25'b00100101_01111111_10100100_0;
      patterns[9602] = 25'b00100101_10000000_10100101_0;
      patterns[9603] = 25'b00100101_10000001_10100110_0;
      patterns[9604] = 25'b00100101_10000010_10100111_0;
      patterns[9605] = 25'b00100101_10000011_10101000_0;
      patterns[9606] = 25'b00100101_10000100_10101001_0;
      patterns[9607] = 25'b00100101_10000101_10101010_0;
      patterns[9608] = 25'b00100101_10000110_10101011_0;
      patterns[9609] = 25'b00100101_10000111_10101100_0;
      patterns[9610] = 25'b00100101_10001000_10101101_0;
      patterns[9611] = 25'b00100101_10001001_10101110_0;
      patterns[9612] = 25'b00100101_10001010_10101111_0;
      patterns[9613] = 25'b00100101_10001011_10110000_0;
      patterns[9614] = 25'b00100101_10001100_10110001_0;
      patterns[9615] = 25'b00100101_10001101_10110010_0;
      patterns[9616] = 25'b00100101_10001110_10110011_0;
      patterns[9617] = 25'b00100101_10001111_10110100_0;
      patterns[9618] = 25'b00100101_10010000_10110101_0;
      patterns[9619] = 25'b00100101_10010001_10110110_0;
      patterns[9620] = 25'b00100101_10010010_10110111_0;
      patterns[9621] = 25'b00100101_10010011_10111000_0;
      patterns[9622] = 25'b00100101_10010100_10111001_0;
      patterns[9623] = 25'b00100101_10010101_10111010_0;
      patterns[9624] = 25'b00100101_10010110_10111011_0;
      patterns[9625] = 25'b00100101_10010111_10111100_0;
      patterns[9626] = 25'b00100101_10011000_10111101_0;
      patterns[9627] = 25'b00100101_10011001_10111110_0;
      patterns[9628] = 25'b00100101_10011010_10111111_0;
      patterns[9629] = 25'b00100101_10011011_11000000_0;
      patterns[9630] = 25'b00100101_10011100_11000001_0;
      patterns[9631] = 25'b00100101_10011101_11000010_0;
      patterns[9632] = 25'b00100101_10011110_11000011_0;
      patterns[9633] = 25'b00100101_10011111_11000100_0;
      patterns[9634] = 25'b00100101_10100000_11000101_0;
      patterns[9635] = 25'b00100101_10100001_11000110_0;
      patterns[9636] = 25'b00100101_10100010_11000111_0;
      patterns[9637] = 25'b00100101_10100011_11001000_0;
      patterns[9638] = 25'b00100101_10100100_11001001_0;
      patterns[9639] = 25'b00100101_10100101_11001010_0;
      patterns[9640] = 25'b00100101_10100110_11001011_0;
      patterns[9641] = 25'b00100101_10100111_11001100_0;
      patterns[9642] = 25'b00100101_10101000_11001101_0;
      patterns[9643] = 25'b00100101_10101001_11001110_0;
      patterns[9644] = 25'b00100101_10101010_11001111_0;
      patterns[9645] = 25'b00100101_10101011_11010000_0;
      patterns[9646] = 25'b00100101_10101100_11010001_0;
      patterns[9647] = 25'b00100101_10101101_11010010_0;
      patterns[9648] = 25'b00100101_10101110_11010011_0;
      patterns[9649] = 25'b00100101_10101111_11010100_0;
      patterns[9650] = 25'b00100101_10110000_11010101_0;
      patterns[9651] = 25'b00100101_10110001_11010110_0;
      patterns[9652] = 25'b00100101_10110010_11010111_0;
      patterns[9653] = 25'b00100101_10110011_11011000_0;
      patterns[9654] = 25'b00100101_10110100_11011001_0;
      patterns[9655] = 25'b00100101_10110101_11011010_0;
      patterns[9656] = 25'b00100101_10110110_11011011_0;
      patterns[9657] = 25'b00100101_10110111_11011100_0;
      patterns[9658] = 25'b00100101_10111000_11011101_0;
      patterns[9659] = 25'b00100101_10111001_11011110_0;
      patterns[9660] = 25'b00100101_10111010_11011111_0;
      patterns[9661] = 25'b00100101_10111011_11100000_0;
      patterns[9662] = 25'b00100101_10111100_11100001_0;
      patterns[9663] = 25'b00100101_10111101_11100010_0;
      patterns[9664] = 25'b00100101_10111110_11100011_0;
      patterns[9665] = 25'b00100101_10111111_11100100_0;
      patterns[9666] = 25'b00100101_11000000_11100101_0;
      patterns[9667] = 25'b00100101_11000001_11100110_0;
      patterns[9668] = 25'b00100101_11000010_11100111_0;
      patterns[9669] = 25'b00100101_11000011_11101000_0;
      patterns[9670] = 25'b00100101_11000100_11101001_0;
      patterns[9671] = 25'b00100101_11000101_11101010_0;
      patterns[9672] = 25'b00100101_11000110_11101011_0;
      patterns[9673] = 25'b00100101_11000111_11101100_0;
      patterns[9674] = 25'b00100101_11001000_11101101_0;
      patterns[9675] = 25'b00100101_11001001_11101110_0;
      patterns[9676] = 25'b00100101_11001010_11101111_0;
      patterns[9677] = 25'b00100101_11001011_11110000_0;
      patterns[9678] = 25'b00100101_11001100_11110001_0;
      patterns[9679] = 25'b00100101_11001101_11110010_0;
      patterns[9680] = 25'b00100101_11001110_11110011_0;
      patterns[9681] = 25'b00100101_11001111_11110100_0;
      patterns[9682] = 25'b00100101_11010000_11110101_0;
      patterns[9683] = 25'b00100101_11010001_11110110_0;
      patterns[9684] = 25'b00100101_11010010_11110111_0;
      patterns[9685] = 25'b00100101_11010011_11111000_0;
      patterns[9686] = 25'b00100101_11010100_11111001_0;
      patterns[9687] = 25'b00100101_11010101_11111010_0;
      patterns[9688] = 25'b00100101_11010110_11111011_0;
      patterns[9689] = 25'b00100101_11010111_11111100_0;
      patterns[9690] = 25'b00100101_11011000_11111101_0;
      patterns[9691] = 25'b00100101_11011001_11111110_0;
      patterns[9692] = 25'b00100101_11011010_11111111_0;
      patterns[9693] = 25'b00100101_11011011_00000000_1;
      patterns[9694] = 25'b00100101_11011100_00000001_1;
      patterns[9695] = 25'b00100101_11011101_00000010_1;
      patterns[9696] = 25'b00100101_11011110_00000011_1;
      patterns[9697] = 25'b00100101_11011111_00000100_1;
      patterns[9698] = 25'b00100101_11100000_00000101_1;
      patterns[9699] = 25'b00100101_11100001_00000110_1;
      patterns[9700] = 25'b00100101_11100010_00000111_1;
      patterns[9701] = 25'b00100101_11100011_00001000_1;
      patterns[9702] = 25'b00100101_11100100_00001001_1;
      patterns[9703] = 25'b00100101_11100101_00001010_1;
      patterns[9704] = 25'b00100101_11100110_00001011_1;
      patterns[9705] = 25'b00100101_11100111_00001100_1;
      patterns[9706] = 25'b00100101_11101000_00001101_1;
      patterns[9707] = 25'b00100101_11101001_00001110_1;
      patterns[9708] = 25'b00100101_11101010_00001111_1;
      patterns[9709] = 25'b00100101_11101011_00010000_1;
      patterns[9710] = 25'b00100101_11101100_00010001_1;
      patterns[9711] = 25'b00100101_11101101_00010010_1;
      patterns[9712] = 25'b00100101_11101110_00010011_1;
      patterns[9713] = 25'b00100101_11101111_00010100_1;
      patterns[9714] = 25'b00100101_11110000_00010101_1;
      patterns[9715] = 25'b00100101_11110001_00010110_1;
      patterns[9716] = 25'b00100101_11110010_00010111_1;
      patterns[9717] = 25'b00100101_11110011_00011000_1;
      patterns[9718] = 25'b00100101_11110100_00011001_1;
      patterns[9719] = 25'b00100101_11110101_00011010_1;
      patterns[9720] = 25'b00100101_11110110_00011011_1;
      patterns[9721] = 25'b00100101_11110111_00011100_1;
      patterns[9722] = 25'b00100101_11111000_00011101_1;
      patterns[9723] = 25'b00100101_11111001_00011110_1;
      patterns[9724] = 25'b00100101_11111010_00011111_1;
      patterns[9725] = 25'b00100101_11111011_00100000_1;
      patterns[9726] = 25'b00100101_11111100_00100001_1;
      patterns[9727] = 25'b00100101_11111101_00100010_1;
      patterns[9728] = 25'b00100101_11111110_00100011_1;
      patterns[9729] = 25'b00100101_11111111_00100100_1;
      patterns[9730] = 25'b00100110_00000000_00100110_0;
      patterns[9731] = 25'b00100110_00000001_00100111_0;
      patterns[9732] = 25'b00100110_00000010_00101000_0;
      patterns[9733] = 25'b00100110_00000011_00101001_0;
      patterns[9734] = 25'b00100110_00000100_00101010_0;
      patterns[9735] = 25'b00100110_00000101_00101011_0;
      patterns[9736] = 25'b00100110_00000110_00101100_0;
      patterns[9737] = 25'b00100110_00000111_00101101_0;
      patterns[9738] = 25'b00100110_00001000_00101110_0;
      patterns[9739] = 25'b00100110_00001001_00101111_0;
      patterns[9740] = 25'b00100110_00001010_00110000_0;
      patterns[9741] = 25'b00100110_00001011_00110001_0;
      patterns[9742] = 25'b00100110_00001100_00110010_0;
      patterns[9743] = 25'b00100110_00001101_00110011_0;
      patterns[9744] = 25'b00100110_00001110_00110100_0;
      patterns[9745] = 25'b00100110_00001111_00110101_0;
      patterns[9746] = 25'b00100110_00010000_00110110_0;
      patterns[9747] = 25'b00100110_00010001_00110111_0;
      patterns[9748] = 25'b00100110_00010010_00111000_0;
      patterns[9749] = 25'b00100110_00010011_00111001_0;
      patterns[9750] = 25'b00100110_00010100_00111010_0;
      patterns[9751] = 25'b00100110_00010101_00111011_0;
      patterns[9752] = 25'b00100110_00010110_00111100_0;
      patterns[9753] = 25'b00100110_00010111_00111101_0;
      patterns[9754] = 25'b00100110_00011000_00111110_0;
      patterns[9755] = 25'b00100110_00011001_00111111_0;
      patterns[9756] = 25'b00100110_00011010_01000000_0;
      patterns[9757] = 25'b00100110_00011011_01000001_0;
      patterns[9758] = 25'b00100110_00011100_01000010_0;
      patterns[9759] = 25'b00100110_00011101_01000011_0;
      patterns[9760] = 25'b00100110_00011110_01000100_0;
      patterns[9761] = 25'b00100110_00011111_01000101_0;
      patterns[9762] = 25'b00100110_00100000_01000110_0;
      patterns[9763] = 25'b00100110_00100001_01000111_0;
      patterns[9764] = 25'b00100110_00100010_01001000_0;
      patterns[9765] = 25'b00100110_00100011_01001001_0;
      patterns[9766] = 25'b00100110_00100100_01001010_0;
      patterns[9767] = 25'b00100110_00100101_01001011_0;
      patterns[9768] = 25'b00100110_00100110_01001100_0;
      patterns[9769] = 25'b00100110_00100111_01001101_0;
      patterns[9770] = 25'b00100110_00101000_01001110_0;
      patterns[9771] = 25'b00100110_00101001_01001111_0;
      patterns[9772] = 25'b00100110_00101010_01010000_0;
      patterns[9773] = 25'b00100110_00101011_01010001_0;
      patterns[9774] = 25'b00100110_00101100_01010010_0;
      patterns[9775] = 25'b00100110_00101101_01010011_0;
      patterns[9776] = 25'b00100110_00101110_01010100_0;
      patterns[9777] = 25'b00100110_00101111_01010101_0;
      patterns[9778] = 25'b00100110_00110000_01010110_0;
      patterns[9779] = 25'b00100110_00110001_01010111_0;
      patterns[9780] = 25'b00100110_00110010_01011000_0;
      patterns[9781] = 25'b00100110_00110011_01011001_0;
      patterns[9782] = 25'b00100110_00110100_01011010_0;
      patterns[9783] = 25'b00100110_00110101_01011011_0;
      patterns[9784] = 25'b00100110_00110110_01011100_0;
      patterns[9785] = 25'b00100110_00110111_01011101_0;
      patterns[9786] = 25'b00100110_00111000_01011110_0;
      patterns[9787] = 25'b00100110_00111001_01011111_0;
      patterns[9788] = 25'b00100110_00111010_01100000_0;
      patterns[9789] = 25'b00100110_00111011_01100001_0;
      patterns[9790] = 25'b00100110_00111100_01100010_0;
      patterns[9791] = 25'b00100110_00111101_01100011_0;
      patterns[9792] = 25'b00100110_00111110_01100100_0;
      patterns[9793] = 25'b00100110_00111111_01100101_0;
      patterns[9794] = 25'b00100110_01000000_01100110_0;
      patterns[9795] = 25'b00100110_01000001_01100111_0;
      patterns[9796] = 25'b00100110_01000010_01101000_0;
      patterns[9797] = 25'b00100110_01000011_01101001_0;
      patterns[9798] = 25'b00100110_01000100_01101010_0;
      patterns[9799] = 25'b00100110_01000101_01101011_0;
      patterns[9800] = 25'b00100110_01000110_01101100_0;
      patterns[9801] = 25'b00100110_01000111_01101101_0;
      patterns[9802] = 25'b00100110_01001000_01101110_0;
      patterns[9803] = 25'b00100110_01001001_01101111_0;
      patterns[9804] = 25'b00100110_01001010_01110000_0;
      patterns[9805] = 25'b00100110_01001011_01110001_0;
      patterns[9806] = 25'b00100110_01001100_01110010_0;
      patterns[9807] = 25'b00100110_01001101_01110011_0;
      patterns[9808] = 25'b00100110_01001110_01110100_0;
      patterns[9809] = 25'b00100110_01001111_01110101_0;
      patterns[9810] = 25'b00100110_01010000_01110110_0;
      patterns[9811] = 25'b00100110_01010001_01110111_0;
      patterns[9812] = 25'b00100110_01010010_01111000_0;
      patterns[9813] = 25'b00100110_01010011_01111001_0;
      patterns[9814] = 25'b00100110_01010100_01111010_0;
      patterns[9815] = 25'b00100110_01010101_01111011_0;
      patterns[9816] = 25'b00100110_01010110_01111100_0;
      patterns[9817] = 25'b00100110_01010111_01111101_0;
      patterns[9818] = 25'b00100110_01011000_01111110_0;
      patterns[9819] = 25'b00100110_01011001_01111111_0;
      patterns[9820] = 25'b00100110_01011010_10000000_0;
      patterns[9821] = 25'b00100110_01011011_10000001_0;
      patterns[9822] = 25'b00100110_01011100_10000010_0;
      patterns[9823] = 25'b00100110_01011101_10000011_0;
      patterns[9824] = 25'b00100110_01011110_10000100_0;
      patterns[9825] = 25'b00100110_01011111_10000101_0;
      patterns[9826] = 25'b00100110_01100000_10000110_0;
      patterns[9827] = 25'b00100110_01100001_10000111_0;
      patterns[9828] = 25'b00100110_01100010_10001000_0;
      patterns[9829] = 25'b00100110_01100011_10001001_0;
      patterns[9830] = 25'b00100110_01100100_10001010_0;
      patterns[9831] = 25'b00100110_01100101_10001011_0;
      patterns[9832] = 25'b00100110_01100110_10001100_0;
      patterns[9833] = 25'b00100110_01100111_10001101_0;
      patterns[9834] = 25'b00100110_01101000_10001110_0;
      patterns[9835] = 25'b00100110_01101001_10001111_0;
      patterns[9836] = 25'b00100110_01101010_10010000_0;
      patterns[9837] = 25'b00100110_01101011_10010001_0;
      patterns[9838] = 25'b00100110_01101100_10010010_0;
      patterns[9839] = 25'b00100110_01101101_10010011_0;
      patterns[9840] = 25'b00100110_01101110_10010100_0;
      patterns[9841] = 25'b00100110_01101111_10010101_0;
      patterns[9842] = 25'b00100110_01110000_10010110_0;
      patterns[9843] = 25'b00100110_01110001_10010111_0;
      patterns[9844] = 25'b00100110_01110010_10011000_0;
      patterns[9845] = 25'b00100110_01110011_10011001_0;
      patterns[9846] = 25'b00100110_01110100_10011010_0;
      patterns[9847] = 25'b00100110_01110101_10011011_0;
      patterns[9848] = 25'b00100110_01110110_10011100_0;
      patterns[9849] = 25'b00100110_01110111_10011101_0;
      patterns[9850] = 25'b00100110_01111000_10011110_0;
      patterns[9851] = 25'b00100110_01111001_10011111_0;
      patterns[9852] = 25'b00100110_01111010_10100000_0;
      patterns[9853] = 25'b00100110_01111011_10100001_0;
      patterns[9854] = 25'b00100110_01111100_10100010_0;
      patterns[9855] = 25'b00100110_01111101_10100011_0;
      patterns[9856] = 25'b00100110_01111110_10100100_0;
      patterns[9857] = 25'b00100110_01111111_10100101_0;
      patterns[9858] = 25'b00100110_10000000_10100110_0;
      patterns[9859] = 25'b00100110_10000001_10100111_0;
      patterns[9860] = 25'b00100110_10000010_10101000_0;
      patterns[9861] = 25'b00100110_10000011_10101001_0;
      patterns[9862] = 25'b00100110_10000100_10101010_0;
      patterns[9863] = 25'b00100110_10000101_10101011_0;
      patterns[9864] = 25'b00100110_10000110_10101100_0;
      patterns[9865] = 25'b00100110_10000111_10101101_0;
      patterns[9866] = 25'b00100110_10001000_10101110_0;
      patterns[9867] = 25'b00100110_10001001_10101111_0;
      patterns[9868] = 25'b00100110_10001010_10110000_0;
      patterns[9869] = 25'b00100110_10001011_10110001_0;
      patterns[9870] = 25'b00100110_10001100_10110010_0;
      patterns[9871] = 25'b00100110_10001101_10110011_0;
      patterns[9872] = 25'b00100110_10001110_10110100_0;
      patterns[9873] = 25'b00100110_10001111_10110101_0;
      patterns[9874] = 25'b00100110_10010000_10110110_0;
      patterns[9875] = 25'b00100110_10010001_10110111_0;
      patterns[9876] = 25'b00100110_10010010_10111000_0;
      patterns[9877] = 25'b00100110_10010011_10111001_0;
      patterns[9878] = 25'b00100110_10010100_10111010_0;
      patterns[9879] = 25'b00100110_10010101_10111011_0;
      patterns[9880] = 25'b00100110_10010110_10111100_0;
      patterns[9881] = 25'b00100110_10010111_10111101_0;
      patterns[9882] = 25'b00100110_10011000_10111110_0;
      patterns[9883] = 25'b00100110_10011001_10111111_0;
      patterns[9884] = 25'b00100110_10011010_11000000_0;
      patterns[9885] = 25'b00100110_10011011_11000001_0;
      patterns[9886] = 25'b00100110_10011100_11000010_0;
      patterns[9887] = 25'b00100110_10011101_11000011_0;
      patterns[9888] = 25'b00100110_10011110_11000100_0;
      patterns[9889] = 25'b00100110_10011111_11000101_0;
      patterns[9890] = 25'b00100110_10100000_11000110_0;
      patterns[9891] = 25'b00100110_10100001_11000111_0;
      patterns[9892] = 25'b00100110_10100010_11001000_0;
      patterns[9893] = 25'b00100110_10100011_11001001_0;
      patterns[9894] = 25'b00100110_10100100_11001010_0;
      patterns[9895] = 25'b00100110_10100101_11001011_0;
      patterns[9896] = 25'b00100110_10100110_11001100_0;
      patterns[9897] = 25'b00100110_10100111_11001101_0;
      patterns[9898] = 25'b00100110_10101000_11001110_0;
      patterns[9899] = 25'b00100110_10101001_11001111_0;
      patterns[9900] = 25'b00100110_10101010_11010000_0;
      patterns[9901] = 25'b00100110_10101011_11010001_0;
      patterns[9902] = 25'b00100110_10101100_11010010_0;
      patterns[9903] = 25'b00100110_10101101_11010011_0;
      patterns[9904] = 25'b00100110_10101110_11010100_0;
      patterns[9905] = 25'b00100110_10101111_11010101_0;
      patterns[9906] = 25'b00100110_10110000_11010110_0;
      patterns[9907] = 25'b00100110_10110001_11010111_0;
      patterns[9908] = 25'b00100110_10110010_11011000_0;
      patterns[9909] = 25'b00100110_10110011_11011001_0;
      patterns[9910] = 25'b00100110_10110100_11011010_0;
      patterns[9911] = 25'b00100110_10110101_11011011_0;
      patterns[9912] = 25'b00100110_10110110_11011100_0;
      patterns[9913] = 25'b00100110_10110111_11011101_0;
      patterns[9914] = 25'b00100110_10111000_11011110_0;
      patterns[9915] = 25'b00100110_10111001_11011111_0;
      patterns[9916] = 25'b00100110_10111010_11100000_0;
      patterns[9917] = 25'b00100110_10111011_11100001_0;
      patterns[9918] = 25'b00100110_10111100_11100010_0;
      patterns[9919] = 25'b00100110_10111101_11100011_0;
      patterns[9920] = 25'b00100110_10111110_11100100_0;
      patterns[9921] = 25'b00100110_10111111_11100101_0;
      patterns[9922] = 25'b00100110_11000000_11100110_0;
      patterns[9923] = 25'b00100110_11000001_11100111_0;
      patterns[9924] = 25'b00100110_11000010_11101000_0;
      patterns[9925] = 25'b00100110_11000011_11101001_0;
      patterns[9926] = 25'b00100110_11000100_11101010_0;
      patterns[9927] = 25'b00100110_11000101_11101011_0;
      patterns[9928] = 25'b00100110_11000110_11101100_0;
      patterns[9929] = 25'b00100110_11000111_11101101_0;
      patterns[9930] = 25'b00100110_11001000_11101110_0;
      patterns[9931] = 25'b00100110_11001001_11101111_0;
      patterns[9932] = 25'b00100110_11001010_11110000_0;
      patterns[9933] = 25'b00100110_11001011_11110001_0;
      patterns[9934] = 25'b00100110_11001100_11110010_0;
      patterns[9935] = 25'b00100110_11001101_11110011_0;
      patterns[9936] = 25'b00100110_11001110_11110100_0;
      patterns[9937] = 25'b00100110_11001111_11110101_0;
      patterns[9938] = 25'b00100110_11010000_11110110_0;
      patterns[9939] = 25'b00100110_11010001_11110111_0;
      patterns[9940] = 25'b00100110_11010010_11111000_0;
      patterns[9941] = 25'b00100110_11010011_11111001_0;
      patterns[9942] = 25'b00100110_11010100_11111010_0;
      patterns[9943] = 25'b00100110_11010101_11111011_0;
      patterns[9944] = 25'b00100110_11010110_11111100_0;
      patterns[9945] = 25'b00100110_11010111_11111101_0;
      patterns[9946] = 25'b00100110_11011000_11111110_0;
      patterns[9947] = 25'b00100110_11011001_11111111_0;
      patterns[9948] = 25'b00100110_11011010_00000000_1;
      patterns[9949] = 25'b00100110_11011011_00000001_1;
      patterns[9950] = 25'b00100110_11011100_00000010_1;
      patterns[9951] = 25'b00100110_11011101_00000011_1;
      patterns[9952] = 25'b00100110_11011110_00000100_1;
      patterns[9953] = 25'b00100110_11011111_00000101_1;
      patterns[9954] = 25'b00100110_11100000_00000110_1;
      patterns[9955] = 25'b00100110_11100001_00000111_1;
      patterns[9956] = 25'b00100110_11100010_00001000_1;
      patterns[9957] = 25'b00100110_11100011_00001001_1;
      patterns[9958] = 25'b00100110_11100100_00001010_1;
      patterns[9959] = 25'b00100110_11100101_00001011_1;
      patterns[9960] = 25'b00100110_11100110_00001100_1;
      patterns[9961] = 25'b00100110_11100111_00001101_1;
      patterns[9962] = 25'b00100110_11101000_00001110_1;
      patterns[9963] = 25'b00100110_11101001_00001111_1;
      patterns[9964] = 25'b00100110_11101010_00010000_1;
      patterns[9965] = 25'b00100110_11101011_00010001_1;
      patterns[9966] = 25'b00100110_11101100_00010010_1;
      patterns[9967] = 25'b00100110_11101101_00010011_1;
      patterns[9968] = 25'b00100110_11101110_00010100_1;
      patterns[9969] = 25'b00100110_11101111_00010101_1;
      patterns[9970] = 25'b00100110_11110000_00010110_1;
      patterns[9971] = 25'b00100110_11110001_00010111_1;
      patterns[9972] = 25'b00100110_11110010_00011000_1;
      patterns[9973] = 25'b00100110_11110011_00011001_1;
      patterns[9974] = 25'b00100110_11110100_00011010_1;
      patterns[9975] = 25'b00100110_11110101_00011011_1;
      patterns[9976] = 25'b00100110_11110110_00011100_1;
      patterns[9977] = 25'b00100110_11110111_00011101_1;
      patterns[9978] = 25'b00100110_11111000_00011110_1;
      patterns[9979] = 25'b00100110_11111001_00011111_1;
      patterns[9980] = 25'b00100110_11111010_00100000_1;
      patterns[9981] = 25'b00100110_11111011_00100001_1;
      patterns[9982] = 25'b00100110_11111100_00100010_1;
      patterns[9983] = 25'b00100110_11111101_00100011_1;
      patterns[9984] = 25'b00100110_11111110_00100100_1;
      patterns[9985] = 25'b00100110_11111111_00100101_1;
      patterns[9986] = 25'b00100111_00000000_00100111_0;
      patterns[9987] = 25'b00100111_00000001_00101000_0;
      patterns[9988] = 25'b00100111_00000010_00101001_0;
      patterns[9989] = 25'b00100111_00000011_00101010_0;
      patterns[9990] = 25'b00100111_00000100_00101011_0;
      patterns[9991] = 25'b00100111_00000101_00101100_0;
      patterns[9992] = 25'b00100111_00000110_00101101_0;
      patterns[9993] = 25'b00100111_00000111_00101110_0;
      patterns[9994] = 25'b00100111_00001000_00101111_0;
      patterns[9995] = 25'b00100111_00001001_00110000_0;
      patterns[9996] = 25'b00100111_00001010_00110001_0;
      patterns[9997] = 25'b00100111_00001011_00110010_0;
      patterns[9998] = 25'b00100111_00001100_00110011_0;
      patterns[9999] = 25'b00100111_00001101_00110100_0;
      patterns[10000] = 25'b00100111_00001110_00110101_0;
      patterns[10001] = 25'b00100111_00001111_00110110_0;
      patterns[10002] = 25'b00100111_00010000_00110111_0;
      patterns[10003] = 25'b00100111_00010001_00111000_0;
      patterns[10004] = 25'b00100111_00010010_00111001_0;
      patterns[10005] = 25'b00100111_00010011_00111010_0;
      patterns[10006] = 25'b00100111_00010100_00111011_0;
      patterns[10007] = 25'b00100111_00010101_00111100_0;
      patterns[10008] = 25'b00100111_00010110_00111101_0;
      patterns[10009] = 25'b00100111_00010111_00111110_0;
      patterns[10010] = 25'b00100111_00011000_00111111_0;
      patterns[10011] = 25'b00100111_00011001_01000000_0;
      patterns[10012] = 25'b00100111_00011010_01000001_0;
      patterns[10013] = 25'b00100111_00011011_01000010_0;
      patterns[10014] = 25'b00100111_00011100_01000011_0;
      patterns[10015] = 25'b00100111_00011101_01000100_0;
      patterns[10016] = 25'b00100111_00011110_01000101_0;
      patterns[10017] = 25'b00100111_00011111_01000110_0;
      patterns[10018] = 25'b00100111_00100000_01000111_0;
      patterns[10019] = 25'b00100111_00100001_01001000_0;
      patterns[10020] = 25'b00100111_00100010_01001001_0;
      patterns[10021] = 25'b00100111_00100011_01001010_0;
      patterns[10022] = 25'b00100111_00100100_01001011_0;
      patterns[10023] = 25'b00100111_00100101_01001100_0;
      patterns[10024] = 25'b00100111_00100110_01001101_0;
      patterns[10025] = 25'b00100111_00100111_01001110_0;
      patterns[10026] = 25'b00100111_00101000_01001111_0;
      patterns[10027] = 25'b00100111_00101001_01010000_0;
      patterns[10028] = 25'b00100111_00101010_01010001_0;
      patterns[10029] = 25'b00100111_00101011_01010010_0;
      patterns[10030] = 25'b00100111_00101100_01010011_0;
      patterns[10031] = 25'b00100111_00101101_01010100_0;
      patterns[10032] = 25'b00100111_00101110_01010101_0;
      patterns[10033] = 25'b00100111_00101111_01010110_0;
      patterns[10034] = 25'b00100111_00110000_01010111_0;
      patterns[10035] = 25'b00100111_00110001_01011000_0;
      patterns[10036] = 25'b00100111_00110010_01011001_0;
      patterns[10037] = 25'b00100111_00110011_01011010_0;
      patterns[10038] = 25'b00100111_00110100_01011011_0;
      patterns[10039] = 25'b00100111_00110101_01011100_0;
      patterns[10040] = 25'b00100111_00110110_01011101_0;
      patterns[10041] = 25'b00100111_00110111_01011110_0;
      patterns[10042] = 25'b00100111_00111000_01011111_0;
      patterns[10043] = 25'b00100111_00111001_01100000_0;
      patterns[10044] = 25'b00100111_00111010_01100001_0;
      patterns[10045] = 25'b00100111_00111011_01100010_0;
      patterns[10046] = 25'b00100111_00111100_01100011_0;
      patterns[10047] = 25'b00100111_00111101_01100100_0;
      patterns[10048] = 25'b00100111_00111110_01100101_0;
      patterns[10049] = 25'b00100111_00111111_01100110_0;
      patterns[10050] = 25'b00100111_01000000_01100111_0;
      patterns[10051] = 25'b00100111_01000001_01101000_0;
      patterns[10052] = 25'b00100111_01000010_01101001_0;
      patterns[10053] = 25'b00100111_01000011_01101010_0;
      patterns[10054] = 25'b00100111_01000100_01101011_0;
      patterns[10055] = 25'b00100111_01000101_01101100_0;
      patterns[10056] = 25'b00100111_01000110_01101101_0;
      patterns[10057] = 25'b00100111_01000111_01101110_0;
      patterns[10058] = 25'b00100111_01001000_01101111_0;
      patterns[10059] = 25'b00100111_01001001_01110000_0;
      patterns[10060] = 25'b00100111_01001010_01110001_0;
      patterns[10061] = 25'b00100111_01001011_01110010_0;
      patterns[10062] = 25'b00100111_01001100_01110011_0;
      patterns[10063] = 25'b00100111_01001101_01110100_0;
      patterns[10064] = 25'b00100111_01001110_01110101_0;
      patterns[10065] = 25'b00100111_01001111_01110110_0;
      patterns[10066] = 25'b00100111_01010000_01110111_0;
      patterns[10067] = 25'b00100111_01010001_01111000_0;
      patterns[10068] = 25'b00100111_01010010_01111001_0;
      patterns[10069] = 25'b00100111_01010011_01111010_0;
      patterns[10070] = 25'b00100111_01010100_01111011_0;
      patterns[10071] = 25'b00100111_01010101_01111100_0;
      patterns[10072] = 25'b00100111_01010110_01111101_0;
      patterns[10073] = 25'b00100111_01010111_01111110_0;
      patterns[10074] = 25'b00100111_01011000_01111111_0;
      patterns[10075] = 25'b00100111_01011001_10000000_0;
      patterns[10076] = 25'b00100111_01011010_10000001_0;
      patterns[10077] = 25'b00100111_01011011_10000010_0;
      patterns[10078] = 25'b00100111_01011100_10000011_0;
      patterns[10079] = 25'b00100111_01011101_10000100_0;
      patterns[10080] = 25'b00100111_01011110_10000101_0;
      patterns[10081] = 25'b00100111_01011111_10000110_0;
      patterns[10082] = 25'b00100111_01100000_10000111_0;
      patterns[10083] = 25'b00100111_01100001_10001000_0;
      patterns[10084] = 25'b00100111_01100010_10001001_0;
      patterns[10085] = 25'b00100111_01100011_10001010_0;
      patterns[10086] = 25'b00100111_01100100_10001011_0;
      patterns[10087] = 25'b00100111_01100101_10001100_0;
      patterns[10088] = 25'b00100111_01100110_10001101_0;
      patterns[10089] = 25'b00100111_01100111_10001110_0;
      patterns[10090] = 25'b00100111_01101000_10001111_0;
      patterns[10091] = 25'b00100111_01101001_10010000_0;
      patterns[10092] = 25'b00100111_01101010_10010001_0;
      patterns[10093] = 25'b00100111_01101011_10010010_0;
      patterns[10094] = 25'b00100111_01101100_10010011_0;
      patterns[10095] = 25'b00100111_01101101_10010100_0;
      patterns[10096] = 25'b00100111_01101110_10010101_0;
      patterns[10097] = 25'b00100111_01101111_10010110_0;
      patterns[10098] = 25'b00100111_01110000_10010111_0;
      patterns[10099] = 25'b00100111_01110001_10011000_0;
      patterns[10100] = 25'b00100111_01110010_10011001_0;
      patterns[10101] = 25'b00100111_01110011_10011010_0;
      patterns[10102] = 25'b00100111_01110100_10011011_0;
      patterns[10103] = 25'b00100111_01110101_10011100_0;
      patterns[10104] = 25'b00100111_01110110_10011101_0;
      patterns[10105] = 25'b00100111_01110111_10011110_0;
      patterns[10106] = 25'b00100111_01111000_10011111_0;
      patterns[10107] = 25'b00100111_01111001_10100000_0;
      patterns[10108] = 25'b00100111_01111010_10100001_0;
      patterns[10109] = 25'b00100111_01111011_10100010_0;
      patterns[10110] = 25'b00100111_01111100_10100011_0;
      patterns[10111] = 25'b00100111_01111101_10100100_0;
      patterns[10112] = 25'b00100111_01111110_10100101_0;
      patterns[10113] = 25'b00100111_01111111_10100110_0;
      patterns[10114] = 25'b00100111_10000000_10100111_0;
      patterns[10115] = 25'b00100111_10000001_10101000_0;
      patterns[10116] = 25'b00100111_10000010_10101001_0;
      patterns[10117] = 25'b00100111_10000011_10101010_0;
      patterns[10118] = 25'b00100111_10000100_10101011_0;
      patterns[10119] = 25'b00100111_10000101_10101100_0;
      patterns[10120] = 25'b00100111_10000110_10101101_0;
      patterns[10121] = 25'b00100111_10000111_10101110_0;
      patterns[10122] = 25'b00100111_10001000_10101111_0;
      patterns[10123] = 25'b00100111_10001001_10110000_0;
      patterns[10124] = 25'b00100111_10001010_10110001_0;
      patterns[10125] = 25'b00100111_10001011_10110010_0;
      patterns[10126] = 25'b00100111_10001100_10110011_0;
      patterns[10127] = 25'b00100111_10001101_10110100_0;
      patterns[10128] = 25'b00100111_10001110_10110101_0;
      patterns[10129] = 25'b00100111_10001111_10110110_0;
      patterns[10130] = 25'b00100111_10010000_10110111_0;
      patterns[10131] = 25'b00100111_10010001_10111000_0;
      patterns[10132] = 25'b00100111_10010010_10111001_0;
      patterns[10133] = 25'b00100111_10010011_10111010_0;
      patterns[10134] = 25'b00100111_10010100_10111011_0;
      patterns[10135] = 25'b00100111_10010101_10111100_0;
      patterns[10136] = 25'b00100111_10010110_10111101_0;
      patterns[10137] = 25'b00100111_10010111_10111110_0;
      patterns[10138] = 25'b00100111_10011000_10111111_0;
      patterns[10139] = 25'b00100111_10011001_11000000_0;
      patterns[10140] = 25'b00100111_10011010_11000001_0;
      patterns[10141] = 25'b00100111_10011011_11000010_0;
      patterns[10142] = 25'b00100111_10011100_11000011_0;
      patterns[10143] = 25'b00100111_10011101_11000100_0;
      patterns[10144] = 25'b00100111_10011110_11000101_0;
      patterns[10145] = 25'b00100111_10011111_11000110_0;
      patterns[10146] = 25'b00100111_10100000_11000111_0;
      patterns[10147] = 25'b00100111_10100001_11001000_0;
      patterns[10148] = 25'b00100111_10100010_11001001_0;
      patterns[10149] = 25'b00100111_10100011_11001010_0;
      patterns[10150] = 25'b00100111_10100100_11001011_0;
      patterns[10151] = 25'b00100111_10100101_11001100_0;
      patterns[10152] = 25'b00100111_10100110_11001101_0;
      patterns[10153] = 25'b00100111_10100111_11001110_0;
      patterns[10154] = 25'b00100111_10101000_11001111_0;
      patterns[10155] = 25'b00100111_10101001_11010000_0;
      patterns[10156] = 25'b00100111_10101010_11010001_0;
      patterns[10157] = 25'b00100111_10101011_11010010_0;
      patterns[10158] = 25'b00100111_10101100_11010011_0;
      patterns[10159] = 25'b00100111_10101101_11010100_0;
      patterns[10160] = 25'b00100111_10101110_11010101_0;
      patterns[10161] = 25'b00100111_10101111_11010110_0;
      patterns[10162] = 25'b00100111_10110000_11010111_0;
      patterns[10163] = 25'b00100111_10110001_11011000_0;
      patterns[10164] = 25'b00100111_10110010_11011001_0;
      patterns[10165] = 25'b00100111_10110011_11011010_0;
      patterns[10166] = 25'b00100111_10110100_11011011_0;
      patterns[10167] = 25'b00100111_10110101_11011100_0;
      patterns[10168] = 25'b00100111_10110110_11011101_0;
      patterns[10169] = 25'b00100111_10110111_11011110_0;
      patterns[10170] = 25'b00100111_10111000_11011111_0;
      patterns[10171] = 25'b00100111_10111001_11100000_0;
      patterns[10172] = 25'b00100111_10111010_11100001_0;
      patterns[10173] = 25'b00100111_10111011_11100010_0;
      patterns[10174] = 25'b00100111_10111100_11100011_0;
      patterns[10175] = 25'b00100111_10111101_11100100_0;
      patterns[10176] = 25'b00100111_10111110_11100101_0;
      patterns[10177] = 25'b00100111_10111111_11100110_0;
      patterns[10178] = 25'b00100111_11000000_11100111_0;
      patterns[10179] = 25'b00100111_11000001_11101000_0;
      patterns[10180] = 25'b00100111_11000010_11101001_0;
      patterns[10181] = 25'b00100111_11000011_11101010_0;
      patterns[10182] = 25'b00100111_11000100_11101011_0;
      patterns[10183] = 25'b00100111_11000101_11101100_0;
      patterns[10184] = 25'b00100111_11000110_11101101_0;
      patterns[10185] = 25'b00100111_11000111_11101110_0;
      patterns[10186] = 25'b00100111_11001000_11101111_0;
      patterns[10187] = 25'b00100111_11001001_11110000_0;
      patterns[10188] = 25'b00100111_11001010_11110001_0;
      patterns[10189] = 25'b00100111_11001011_11110010_0;
      patterns[10190] = 25'b00100111_11001100_11110011_0;
      patterns[10191] = 25'b00100111_11001101_11110100_0;
      patterns[10192] = 25'b00100111_11001110_11110101_0;
      patterns[10193] = 25'b00100111_11001111_11110110_0;
      patterns[10194] = 25'b00100111_11010000_11110111_0;
      patterns[10195] = 25'b00100111_11010001_11111000_0;
      patterns[10196] = 25'b00100111_11010010_11111001_0;
      patterns[10197] = 25'b00100111_11010011_11111010_0;
      patterns[10198] = 25'b00100111_11010100_11111011_0;
      patterns[10199] = 25'b00100111_11010101_11111100_0;
      patterns[10200] = 25'b00100111_11010110_11111101_0;
      patterns[10201] = 25'b00100111_11010111_11111110_0;
      patterns[10202] = 25'b00100111_11011000_11111111_0;
      patterns[10203] = 25'b00100111_11011001_00000000_1;
      patterns[10204] = 25'b00100111_11011010_00000001_1;
      patterns[10205] = 25'b00100111_11011011_00000010_1;
      patterns[10206] = 25'b00100111_11011100_00000011_1;
      patterns[10207] = 25'b00100111_11011101_00000100_1;
      patterns[10208] = 25'b00100111_11011110_00000101_1;
      patterns[10209] = 25'b00100111_11011111_00000110_1;
      patterns[10210] = 25'b00100111_11100000_00000111_1;
      patterns[10211] = 25'b00100111_11100001_00001000_1;
      patterns[10212] = 25'b00100111_11100010_00001001_1;
      patterns[10213] = 25'b00100111_11100011_00001010_1;
      patterns[10214] = 25'b00100111_11100100_00001011_1;
      patterns[10215] = 25'b00100111_11100101_00001100_1;
      patterns[10216] = 25'b00100111_11100110_00001101_1;
      patterns[10217] = 25'b00100111_11100111_00001110_1;
      patterns[10218] = 25'b00100111_11101000_00001111_1;
      patterns[10219] = 25'b00100111_11101001_00010000_1;
      patterns[10220] = 25'b00100111_11101010_00010001_1;
      patterns[10221] = 25'b00100111_11101011_00010010_1;
      patterns[10222] = 25'b00100111_11101100_00010011_1;
      patterns[10223] = 25'b00100111_11101101_00010100_1;
      patterns[10224] = 25'b00100111_11101110_00010101_1;
      patterns[10225] = 25'b00100111_11101111_00010110_1;
      patterns[10226] = 25'b00100111_11110000_00010111_1;
      patterns[10227] = 25'b00100111_11110001_00011000_1;
      patterns[10228] = 25'b00100111_11110010_00011001_1;
      patterns[10229] = 25'b00100111_11110011_00011010_1;
      patterns[10230] = 25'b00100111_11110100_00011011_1;
      patterns[10231] = 25'b00100111_11110101_00011100_1;
      patterns[10232] = 25'b00100111_11110110_00011101_1;
      patterns[10233] = 25'b00100111_11110111_00011110_1;
      patterns[10234] = 25'b00100111_11111000_00011111_1;
      patterns[10235] = 25'b00100111_11111001_00100000_1;
      patterns[10236] = 25'b00100111_11111010_00100001_1;
      patterns[10237] = 25'b00100111_11111011_00100010_1;
      patterns[10238] = 25'b00100111_11111100_00100011_1;
      patterns[10239] = 25'b00100111_11111101_00100100_1;
      patterns[10240] = 25'b00100111_11111110_00100101_1;
      patterns[10241] = 25'b00100111_11111111_00100110_1;
      patterns[10242] = 25'b00101000_00000000_00101000_0;
      patterns[10243] = 25'b00101000_00000001_00101001_0;
      patterns[10244] = 25'b00101000_00000010_00101010_0;
      patterns[10245] = 25'b00101000_00000011_00101011_0;
      patterns[10246] = 25'b00101000_00000100_00101100_0;
      patterns[10247] = 25'b00101000_00000101_00101101_0;
      patterns[10248] = 25'b00101000_00000110_00101110_0;
      patterns[10249] = 25'b00101000_00000111_00101111_0;
      patterns[10250] = 25'b00101000_00001000_00110000_0;
      patterns[10251] = 25'b00101000_00001001_00110001_0;
      patterns[10252] = 25'b00101000_00001010_00110010_0;
      patterns[10253] = 25'b00101000_00001011_00110011_0;
      patterns[10254] = 25'b00101000_00001100_00110100_0;
      patterns[10255] = 25'b00101000_00001101_00110101_0;
      patterns[10256] = 25'b00101000_00001110_00110110_0;
      patterns[10257] = 25'b00101000_00001111_00110111_0;
      patterns[10258] = 25'b00101000_00010000_00111000_0;
      patterns[10259] = 25'b00101000_00010001_00111001_0;
      patterns[10260] = 25'b00101000_00010010_00111010_0;
      patterns[10261] = 25'b00101000_00010011_00111011_0;
      patterns[10262] = 25'b00101000_00010100_00111100_0;
      patterns[10263] = 25'b00101000_00010101_00111101_0;
      patterns[10264] = 25'b00101000_00010110_00111110_0;
      patterns[10265] = 25'b00101000_00010111_00111111_0;
      patterns[10266] = 25'b00101000_00011000_01000000_0;
      patterns[10267] = 25'b00101000_00011001_01000001_0;
      patterns[10268] = 25'b00101000_00011010_01000010_0;
      patterns[10269] = 25'b00101000_00011011_01000011_0;
      patterns[10270] = 25'b00101000_00011100_01000100_0;
      patterns[10271] = 25'b00101000_00011101_01000101_0;
      patterns[10272] = 25'b00101000_00011110_01000110_0;
      patterns[10273] = 25'b00101000_00011111_01000111_0;
      patterns[10274] = 25'b00101000_00100000_01001000_0;
      patterns[10275] = 25'b00101000_00100001_01001001_0;
      patterns[10276] = 25'b00101000_00100010_01001010_0;
      patterns[10277] = 25'b00101000_00100011_01001011_0;
      patterns[10278] = 25'b00101000_00100100_01001100_0;
      patterns[10279] = 25'b00101000_00100101_01001101_0;
      patterns[10280] = 25'b00101000_00100110_01001110_0;
      patterns[10281] = 25'b00101000_00100111_01001111_0;
      patterns[10282] = 25'b00101000_00101000_01010000_0;
      patterns[10283] = 25'b00101000_00101001_01010001_0;
      patterns[10284] = 25'b00101000_00101010_01010010_0;
      patterns[10285] = 25'b00101000_00101011_01010011_0;
      patterns[10286] = 25'b00101000_00101100_01010100_0;
      patterns[10287] = 25'b00101000_00101101_01010101_0;
      patterns[10288] = 25'b00101000_00101110_01010110_0;
      patterns[10289] = 25'b00101000_00101111_01010111_0;
      patterns[10290] = 25'b00101000_00110000_01011000_0;
      patterns[10291] = 25'b00101000_00110001_01011001_0;
      patterns[10292] = 25'b00101000_00110010_01011010_0;
      patterns[10293] = 25'b00101000_00110011_01011011_0;
      patterns[10294] = 25'b00101000_00110100_01011100_0;
      patterns[10295] = 25'b00101000_00110101_01011101_0;
      patterns[10296] = 25'b00101000_00110110_01011110_0;
      patterns[10297] = 25'b00101000_00110111_01011111_0;
      patterns[10298] = 25'b00101000_00111000_01100000_0;
      patterns[10299] = 25'b00101000_00111001_01100001_0;
      patterns[10300] = 25'b00101000_00111010_01100010_0;
      patterns[10301] = 25'b00101000_00111011_01100011_0;
      patterns[10302] = 25'b00101000_00111100_01100100_0;
      patterns[10303] = 25'b00101000_00111101_01100101_0;
      patterns[10304] = 25'b00101000_00111110_01100110_0;
      patterns[10305] = 25'b00101000_00111111_01100111_0;
      patterns[10306] = 25'b00101000_01000000_01101000_0;
      patterns[10307] = 25'b00101000_01000001_01101001_0;
      patterns[10308] = 25'b00101000_01000010_01101010_0;
      patterns[10309] = 25'b00101000_01000011_01101011_0;
      patterns[10310] = 25'b00101000_01000100_01101100_0;
      patterns[10311] = 25'b00101000_01000101_01101101_0;
      patterns[10312] = 25'b00101000_01000110_01101110_0;
      patterns[10313] = 25'b00101000_01000111_01101111_0;
      patterns[10314] = 25'b00101000_01001000_01110000_0;
      patterns[10315] = 25'b00101000_01001001_01110001_0;
      patterns[10316] = 25'b00101000_01001010_01110010_0;
      patterns[10317] = 25'b00101000_01001011_01110011_0;
      patterns[10318] = 25'b00101000_01001100_01110100_0;
      patterns[10319] = 25'b00101000_01001101_01110101_0;
      patterns[10320] = 25'b00101000_01001110_01110110_0;
      patterns[10321] = 25'b00101000_01001111_01110111_0;
      patterns[10322] = 25'b00101000_01010000_01111000_0;
      patterns[10323] = 25'b00101000_01010001_01111001_0;
      patterns[10324] = 25'b00101000_01010010_01111010_0;
      patterns[10325] = 25'b00101000_01010011_01111011_0;
      patterns[10326] = 25'b00101000_01010100_01111100_0;
      patterns[10327] = 25'b00101000_01010101_01111101_0;
      patterns[10328] = 25'b00101000_01010110_01111110_0;
      patterns[10329] = 25'b00101000_01010111_01111111_0;
      patterns[10330] = 25'b00101000_01011000_10000000_0;
      patterns[10331] = 25'b00101000_01011001_10000001_0;
      patterns[10332] = 25'b00101000_01011010_10000010_0;
      patterns[10333] = 25'b00101000_01011011_10000011_0;
      patterns[10334] = 25'b00101000_01011100_10000100_0;
      patterns[10335] = 25'b00101000_01011101_10000101_0;
      patterns[10336] = 25'b00101000_01011110_10000110_0;
      patterns[10337] = 25'b00101000_01011111_10000111_0;
      patterns[10338] = 25'b00101000_01100000_10001000_0;
      patterns[10339] = 25'b00101000_01100001_10001001_0;
      patterns[10340] = 25'b00101000_01100010_10001010_0;
      patterns[10341] = 25'b00101000_01100011_10001011_0;
      patterns[10342] = 25'b00101000_01100100_10001100_0;
      patterns[10343] = 25'b00101000_01100101_10001101_0;
      patterns[10344] = 25'b00101000_01100110_10001110_0;
      patterns[10345] = 25'b00101000_01100111_10001111_0;
      patterns[10346] = 25'b00101000_01101000_10010000_0;
      patterns[10347] = 25'b00101000_01101001_10010001_0;
      patterns[10348] = 25'b00101000_01101010_10010010_0;
      patterns[10349] = 25'b00101000_01101011_10010011_0;
      patterns[10350] = 25'b00101000_01101100_10010100_0;
      patterns[10351] = 25'b00101000_01101101_10010101_0;
      patterns[10352] = 25'b00101000_01101110_10010110_0;
      patterns[10353] = 25'b00101000_01101111_10010111_0;
      patterns[10354] = 25'b00101000_01110000_10011000_0;
      patterns[10355] = 25'b00101000_01110001_10011001_0;
      patterns[10356] = 25'b00101000_01110010_10011010_0;
      patterns[10357] = 25'b00101000_01110011_10011011_0;
      patterns[10358] = 25'b00101000_01110100_10011100_0;
      patterns[10359] = 25'b00101000_01110101_10011101_0;
      patterns[10360] = 25'b00101000_01110110_10011110_0;
      patterns[10361] = 25'b00101000_01110111_10011111_0;
      patterns[10362] = 25'b00101000_01111000_10100000_0;
      patterns[10363] = 25'b00101000_01111001_10100001_0;
      patterns[10364] = 25'b00101000_01111010_10100010_0;
      patterns[10365] = 25'b00101000_01111011_10100011_0;
      patterns[10366] = 25'b00101000_01111100_10100100_0;
      patterns[10367] = 25'b00101000_01111101_10100101_0;
      patterns[10368] = 25'b00101000_01111110_10100110_0;
      patterns[10369] = 25'b00101000_01111111_10100111_0;
      patterns[10370] = 25'b00101000_10000000_10101000_0;
      patterns[10371] = 25'b00101000_10000001_10101001_0;
      patterns[10372] = 25'b00101000_10000010_10101010_0;
      patterns[10373] = 25'b00101000_10000011_10101011_0;
      patterns[10374] = 25'b00101000_10000100_10101100_0;
      patterns[10375] = 25'b00101000_10000101_10101101_0;
      patterns[10376] = 25'b00101000_10000110_10101110_0;
      patterns[10377] = 25'b00101000_10000111_10101111_0;
      patterns[10378] = 25'b00101000_10001000_10110000_0;
      patterns[10379] = 25'b00101000_10001001_10110001_0;
      patterns[10380] = 25'b00101000_10001010_10110010_0;
      patterns[10381] = 25'b00101000_10001011_10110011_0;
      patterns[10382] = 25'b00101000_10001100_10110100_0;
      patterns[10383] = 25'b00101000_10001101_10110101_0;
      patterns[10384] = 25'b00101000_10001110_10110110_0;
      patterns[10385] = 25'b00101000_10001111_10110111_0;
      patterns[10386] = 25'b00101000_10010000_10111000_0;
      patterns[10387] = 25'b00101000_10010001_10111001_0;
      patterns[10388] = 25'b00101000_10010010_10111010_0;
      patterns[10389] = 25'b00101000_10010011_10111011_0;
      patterns[10390] = 25'b00101000_10010100_10111100_0;
      patterns[10391] = 25'b00101000_10010101_10111101_0;
      patterns[10392] = 25'b00101000_10010110_10111110_0;
      patterns[10393] = 25'b00101000_10010111_10111111_0;
      patterns[10394] = 25'b00101000_10011000_11000000_0;
      patterns[10395] = 25'b00101000_10011001_11000001_0;
      patterns[10396] = 25'b00101000_10011010_11000010_0;
      patterns[10397] = 25'b00101000_10011011_11000011_0;
      patterns[10398] = 25'b00101000_10011100_11000100_0;
      patterns[10399] = 25'b00101000_10011101_11000101_0;
      patterns[10400] = 25'b00101000_10011110_11000110_0;
      patterns[10401] = 25'b00101000_10011111_11000111_0;
      patterns[10402] = 25'b00101000_10100000_11001000_0;
      patterns[10403] = 25'b00101000_10100001_11001001_0;
      patterns[10404] = 25'b00101000_10100010_11001010_0;
      patterns[10405] = 25'b00101000_10100011_11001011_0;
      patterns[10406] = 25'b00101000_10100100_11001100_0;
      patterns[10407] = 25'b00101000_10100101_11001101_0;
      patterns[10408] = 25'b00101000_10100110_11001110_0;
      patterns[10409] = 25'b00101000_10100111_11001111_0;
      patterns[10410] = 25'b00101000_10101000_11010000_0;
      patterns[10411] = 25'b00101000_10101001_11010001_0;
      patterns[10412] = 25'b00101000_10101010_11010010_0;
      patterns[10413] = 25'b00101000_10101011_11010011_0;
      patterns[10414] = 25'b00101000_10101100_11010100_0;
      patterns[10415] = 25'b00101000_10101101_11010101_0;
      patterns[10416] = 25'b00101000_10101110_11010110_0;
      patterns[10417] = 25'b00101000_10101111_11010111_0;
      patterns[10418] = 25'b00101000_10110000_11011000_0;
      patterns[10419] = 25'b00101000_10110001_11011001_0;
      patterns[10420] = 25'b00101000_10110010_11011010_0;
      patterns[10421] = 25'b00101000_10110011_11011011_0;
      patterns[10422] = 25'b00101000_10110100_11011100_0;
      patterns[10423] = 25'b00101000_10110101_11011101_0;
      patterns[10424] = 25'b00101000_10110110_11011110_0;
      patterns[10425] = 25'b00101000_10110111_11011111_0;
      patterns[10426] = 25'b00101000_10111000_11100000_0;
      patterns[10427] = 25'b00101000_10111001_11100001_0;
      patterns[10428] = 25'b00101000_10111010_11100010_0;
      patterns[10429] = 25'b00101000_10111011_11100011_0;
      patterns[10430] = 25'b00101000_10111100_11100100_0;
      patterns[10431] = 25'b00101000_10111101_11100101_0;
      patterns[10432] = 25'b00101000_10111110_11100110_0;
      patterns[10433] = 25'b00101000_10111111_11100111_0;
      patterns[10434] = 25'b00101000_11000000_11101000_0;
      patterns[10435] = 25'b00101000_11000001_11101001_0;
      patterns[10436] = 25'b00101000_11000010_11101010_0;
      patterns[10437] = 25'b00101000_11000011_11101011_0;
      patterns[10438] = 25'b00101000_11000100_11101100_0;
      patterns[10439] = 25'b00101000_11000101_11101101_0;
      patterns[10440] = 25'b00101000_11000110_11101110_0;
      patterns[10441] = 25'b00101000_11000111_11101111_0;
      patterns[10442] = 25'b00101000_11001000_11110000_0;
      patterns[10443] = 25'b00101000_11001001_11110001_0;
      patterns[10444] = 25'b00101000_11001010_11110010_0;
      patterns[10445] = 25'b00101000_11001011_11110011_0;
      patterns[10446] = 25'b00101000_11001100_11110100_0;
      patterns[10447] = 25'b00101000_11001101_11110101_0;
      patterns[10448] = 25'b00101000_11001110_11110110_0;
      patterns[10449] = 25'b00101000_11001111_11110111_0;
      patterns[10450] = 25'b00101000_11010000_11111000_0;
      patterns[10451] = 25'b00101000_11010001_11111001_0;
      patterns[10452] = 25'b00101000_11010010_11111010_0;
      patterns[10453] = 25'b00101000_11010011_11111011_0;
      patterns[10454] = 25'b00101000_11010100_11111100_0;
      patterns[10455] = 25'b00101000_11010101_11111101_0;
      patterns[10456] = 25'b00101000_11010110_11111110_0;
      patterns[10457] = 25'b00101000_11010111_11111111_0;
      patterns[10458] = 25'b00101000_11011000_00000000_1;
      patterns[10459] = 25'b00101000_11011001_00000001_1;
      patterns[10460] = 25'b00101000_11011010_00000010_1;
      patterns[10461] = 25'b00101000_11011011_00000011_1;
      patterns[10462] = 25'b00101000_11011100_00000100_1;
      patterns[10463] = 25'b00101000_11011101_00000101_1;
      patterns[10464] = 25'b00101000_11011110_00000110_1;
      patterns[10465] = 25'b00101000_11011111_00000111_1;
      patterns[10466] = 25'b00101000_11100000_00001000_1;
      patterns[10467] = 25'b00101000_11100001_00001001_1;
      patterns[10468] = 25'b00101000_11100010_00001010_1;
      patterns[10469] = 25'b00101000_11100011_00001011_1;
      patterns[10470] = 25'b00101000_11100100_00001100_1;
      patterns[10471] = 25'b00101000_11100101_00001101_1;
      patterns[10472] = 25'b00101000_11100110_00001110_1;
      patterns[10473] = 25'b00101000_11100111_00001111_1;
      patterns[10474] = 25'b00101000_11101000_00010000_1;
      patterns[10475] = 25'b00101000_11101001_00010001_1;
      patterns[10476] = 25'b00101000_11101010_00010010_1;
      patterns[10477] = 25'b00101000_11101011_00010011_1;
      patterns[10478] = 25'b00101000_11101100_00010100_1;
      patterns[10479] = 25'b00101000_11101101_00010101_1;
      patterns[10480] = 25'b00101000_11101110_00010110_1;
      patterns[10481] = 25'b00101000_11101111_00010111_1;
      patterns[10482] = 25'b00101000_11110000_00011000_1;
      patterns[10483] = 25'b00101000_11110001_00011001_1;
      patterns[10484] = 25'b00101000_11110010_00011010_1;
      patterns[10485] = 25'b00101000_11110011_00011011_1;
      patterns[10486] = 25'b00101000_11110100_00011100_1;
      patterns[10487] = 25'b00101000_11110101_00011101_1;
      patterns[10488] = 25'b00101000_11110110_00011110_1;
      patterns[10489] = 25'b00101000_11110111_00011111_1;
      patterns[10490] = 25'b00101000_11111000_00100000_1;
      patterns[10491] = 25'b00101000_11111001_00100001_1;
      patterns[10492] = 25'b00101000_11111010_00100010_1;
      patterns[10493] = 25'b00101000_11111011_00100011_1;
      patterns[10494] = 25'b00101000_11111100_00100100_1;
      patterns[10495] = 25'b00101000_11111101_00100101_1;
      patterns[10496] = 25'b00101000_11111110_00100110_1;
      patterns[10497] = 25'b00101000_11111111_00100111_1;
      patterns[10498] = 25'b00101001_00000000_00101001_0;
      patterns[10499] = 25'b00101001_00000001_00101010_0;
      patterns[10500] = 25'b00101001_00000010_00101011_0;
      patterns[10501] = 25'b00101001_00000011_00101100_0;
      patterns[10502] = 25'b00101001_00000100_00101101_0;
      patterns[10503] = 25'b00101001_00000101_00101110_0;
      patterns[10504] = 25'b00101001_00000110_00101111_0;
      patterns[10505] = 25'b00101001_00000111_00110000_0;
      patterns[10506] = 25'b00101001_00001000_00110001_0;
      patterns[10507] = 25'b00101001_00001001_00110010_0;
      patterns[10508] = 25'b00101001_00001010_00110011_0;
      patterns[10509] = 25'b00101001_00001011_00110100_0;
      patterns[10510] = 25'b00101001_00001100_00110101_0;
      patterns[10511] = 25'b00101001_00001101_00110110_0;
      patterns[10512] = 25'b00101001_00001110_00110111_0;
      patterns[10513] = 25'b00101001_00001111_00111000_0;
      patterns[10514] = 25'b00101001_00010000_00111001_0;
      patterns[10515] = 25'b00101001_00010001_00111010_0;
      patterns[10516] = 25'b00101001_00010010_00111011_0;
      patterns[10517] = 25'b00101001_00010011_00111100_0;
      patterns[10518] = 25'b00101001_00010100_00111101_0;
      patterns[10519] = 25'b00101001_00010101_00111110_0;
      patterns[10520] = 25'b00101001_00010110_00111111_0;
      patterns[10521] = 25'b00101001_00010111_01000000_0;
      patterns[10522] = 25'b00101001_00011000_01000001_0;
      patterns[10523] = 25'b00101001_00011001_01000010_0;
      patterns[10524] = 25'b00101001_00011010_01000011_0;
      patterns[10525] = 25'b00101001_00011011_01000100_0;
      patterns[10526] = 25'b00101001_00011100_01000101_0;
      patterns[10527] = 25'b00101001_00011101_01000110_0;
      patterns[10528] = 25'b00101001_00011110_01000111_0;
      patterns[10529] = 25'b00101001_00011111_01001000_0;
      patterns[10530] = 25'b00101001_00100000_01001001_0;
      patterns[10531] = 25'b00101001_00100001_01001010_0;
      patterns[10532] = 25'b00101001_00100010_01001011_0;
      patterns[10533] = 25'b00101001_00100011_01001100_0;
      patterns[10534] = 25'b00101001_00100100_01001101_0;
      patterns[10535] = 25'b00101001_00100101_01001110_0;
      patterns[10536] = 25'b00101001_00100110_01001111_0;
      patterns[10537] = 25'b00101001_00100111_01010000_0;
      patterns[10538] = 25'b00101001_00101000_01010001_0;
      patterns[10539] = 25'b00101001_00101001_01010010_0;
      patterns[10540] = 25'b00101001_00101010_01010011_0;
      patterns[10541] = 25'b00101001_00101011_01010100_0;
      patterns[10542] = 25'b00101001_00101100_01010101_0;
      patterns[10543] = 25'b00101001_00101101_01010110_0;
      patterns[10544] = 25'b00101001_00101110_01010111_0;
      patterns[10545] = 25'b00101001_00101111_01011000_0;
      patterns[10546] = 25'b00101001_00110000_01011001_0;
      patterns[10547] = 25'b00101001_00110001_01011010_0;
      patterns[10548] = 25'b00101001_00110010_01011011_0;
      patterns[10549] = 25'b00101001_00110011_01011100_0;
      patterns[10550] = 25'b00101001_00110100_01011101_0;
      patterns[10551] = 25'b00101001_00110101_01011110_0;
      patterns[10552] = 25'b00101001_00110110_01011111_0;
      patterns[10553] = 25'b00101001_00110111_01100000_0;
      patterns[10554] = 25'b00101001_00111000_01100001_0;
      patterns[10555] = 25'b00101001_00111001_01100010_0;
      patterns[10556] = 25'b00101001_00111010_01100011_0;
      patterns[10557] = 25'b00101001_00111011_01100100_0;
      patterns[10558] = 25'b00101001_00111100_01100101_0;
      patterns[10559] = 25'b00101001_00111101_01100110_0;
      patterns[10560] = 25'b00101001_00111110_01100111_0;
      patterns[10561] = 25'b00101001_00111111_01101000_0;
      patterns[10562] = 25'b00101001_01000000_01101001_0;
      patterns[10563] = 25'b00101001_01000001_01101010_0;
      patterns[10564] = 25'b00101001_01000010_01101011_0;
      patterns[10565] = 25'b00101001_01000011_01101100_0;
      patterns[10566] = 25'b00101001_01000100_01101101_0;
      patterns[10567] = 25'b00101001_01000101_01101110_0;
      patterns[10568] = 25'b00101001_01000110_01101111_0;
      patterns[10569] = 25'b00101001_01000111_01110000_0;
      patterns[10570] = 25'b00101001_01001000_01110001_0;
      patterns[10571] = 25'b00101001_01001001_01110010_0;
      patterns[10572] = 25'b00101001_01001010_01110011_0;
      patterns[10573] = 25'b00101001_01001011_01110100_0;
      patterns[10574] = 25'b00101001_01001100_01110101_0;
      patterns[10575] = 25'b00101001_01001101_01110110_0;
      patterns[10576] = 25'b00101001_01001110_01110111_0;
      patterns[10577] = 25'b00101001_01001111_01111000_0;
      patterns[10578] = 25'b00101001_01010000_01111001_0;
      patterns[10579] = 25'b00101001_01010001_01111010_0;
      patterns[10580] = 25'b00101001_01010010_01111011_0;
      patterns[10581] = 25'b00101001_01010011_01111100_0;
      patterns[10582] = 25'b00101001_01010100_01111101_0;
      patterns[10583] = 25'b00101001_01010101_01111110_0;
      patterns[10584] = 25'b00101001_01010110_01111111_0;
      patterns[10585] = 25'b00101001_01010111_10000000_0;
      patterns[10586] = 25'b00101001_01011000_10000001_0;
      patterns[10587] = 25'b00101001_01011001_10000010_0;
      patterns[10588] = 25'b00101001_01011010_10000011_0;
      patterns[10589] = 25'b00101001_01011011_10000100_0;
      patterns[10590] = 25'b00101001_01011100_10000101_0;
      patterns[10591] = 25'b00101001_01011101_10000110_0;
      patterns[10592] = 25'b00101001_01011110_10000111_0;
      patterns[10593] = 25'b00101001_01011111_10001000_0;
      patterns[10594] = 25'b00101001_01100000_10001001_0;
      patterns[10595] = 25'b00101001_01100001_10001010_0;
      patterns[10596] = 25'b00101001_01100010_10001011_0;
      patterns[10597] = 25'b00101001_01100011_10001100_0;
      patterns[10598] = 25'b00101001_01100100_10001101_0;
      patterns[10599] = 25'b00101001_01100101_10001110_0;
      patterns[10600] = 25'b00101001_01100110_10001111_0;
      patterns[10601] = 25'b00101001_01100111_10010000_0;
      patterns[10602] = 25'b00101001_01101000_10010001_0;
      patterns[10603] = 25'b00101001_01101001_10010010_0;
      patterns[10604] = 25'b00101001_01101010_10010011_0;
      patterns[10605] = 25'b00101001_01101011_10010100_0;
      patterns[10606] = 25'b00101001_01101100_10010101_0;
      patterns[10607] = 25'b00101001_01101101_10010110_0;
      patterns[10608] = 25'b00101001_01101110_10010111_0;
      patterns[10609] = 25'b00101001_01101111_10011000_0;
      patterns[10610] = 25'b00101001_01110000_10011001_0;
      patterns[10611] = 25'b00101001_01110001_10011010_0;
      patterns[10612] = 25'b00101001_01110010_10011011_0;
      patterns[10613] = 25'b00101001_01110011_10011100_0;
      patterns[10614] = 25'b00101001_01110100_10011101_0;
      patterns[10615] = 25'b00101001_01110101_10011110_0;
      patterns[10616] = 25'b00101001_01110110_10011111_0;
      patterns[10617] = 25'b00101001_01110111_10100000_0;
      patterns[10618] = 25'b00101001_01111000_10100001_0;
      patterns[10619] = 25'b00101001_01111001_10100010_0;
      patterns[10620] = 25'b00101001_01111010_10100011_0;
      patterns[10621] = 25'b00101001_01111011_10100100_0;
      patterns[10622] = 25'b00101001_01111100_10100101_0;
      patterns[10623] = 25'b00101001_01111101_10100110_0;
      patterns[10624] = 25'b00101001_01111110_10100111_0;
      patterns[10625] = 25'b00101001_01111111_10101000_0;
      patterns[10626] = 25'b00101001_10000000_10101001_0;
      patterns[10627] = 25'b00101001_10000001_10101010_0;
      patterns[10628] = 25'b00101001_10000010_10101011_0;
      patterns[10629] = 25'b00101001_10000011_10101100_0;
      patterns[10630] = 25'b00101001_10000100_10101101_0;
      patterns[10631] = 25'b00101001_10000101_10101110_0;
      patterns[10632] = 25'b00101001_10000110_10101111_0;
      patterns[10633] = 25'b00101001_10000111_10110000_0;
      patterns[10634] = 25'b00101001_10001000_10110001_0;
      patterns[10635] = 25'b00101001_10001001_10110010_0;
      patterns[10636] = 25'b00101001_10001010_10110011_0;
      patterns[10637] = 25'b00101001_10001011_10110100_0;
      patterns[10638] = 25'b00101001_10001100_10110101_0;
      patterns[10639] = 25'b00101001_10001101_10110110_0;
      patterns[10640] = 25'b00101001_10001110_10110111_0;
      patterns[10641] = 25'b00101001_10001111_10111000_0;
      patterns[10642] = 25'b00101001_10010000_10111001_0;
      patterns[10643] = 25'b00101001_10010001_10111010_0;
      patterns[10644] = 25'b00101001_10010010_10111011_0;
      patterns[10645] = 25'b00101001_10010011_10111100_0;
      patterns[10646] = 25'b00101001_10010100_10111101_0;
      patterns[10647] = 25'b00101001_10010101_10111110_0;
      patterns[10648] = 25'b00101001_10010110_10111111_0;
      patterns[10649] = 25'b00101001_10010111_11000000_0;
      patterns[10650] = 25'b00101001_10011000_11000001_0;
      patterns[10651] = 25'b00101001_10011001_11000010_0;
      patterns[10652] = 25'b00101001_10011010_11000011_0;
      patterns[10653] = 25'b00101001_10011011_11000100_0;
      patterns[10654] = 25'b00101001_10011100_11000101_0;
      patterns[10655] = 25'b00101001_10011101_11000110_0;
      patterns[10656] = 25'b00101001_10011110_11000111_0;
      patterns[10657] = 25'b00101001_10011111_11001000_0;
      patterns[10658] = 25'b00101001_10100000_11001001_0;
      patterns[10659] = 25'b00101001_10100001_11001010_0;
      patterns[10660] = 25'b00101001_10100010_11001011_0;
      patterns[10661] = 25'b00101001_10100011_11001100_0;
      patterns[10662] = 25'b00101001_10100100_11001101_0;
      patterns[10663] = 25'b00101001_10100101_11001110_0;
      patterns[10664] = 25'b00101001_10100110_11001111_0;
      patterns[10665] = 25'b00101001_10100111_11010000_0;
      patterns[10666] = 25'b00101001_10101000_11010001_0;
      patterns[10667] = 25'b00101001_10101001_11010010_0;
      patterns[10668] = 25'b00101001_10101010_11010011_0;
      patterns[10669] = 25'b00101001_10101011_11010100_0;
      patterns[10670] = 25'b00101001_10101100_11010101_0;
      patterns[10671] = 25'b00101001_10101101_11010110_0;
      patterns[10672] = 25'b00101001_10101110_11010111_0;
      patterns[10673] = 25'b00101001_10101111_11011000_0;
      patterns[10674] = 25'b00101001_10110000_11011001_0;
      patterns[10675] = 25'b00101001_10110001_11011010_0;
      patterns[10676] = 25'b00101001_10110010_11011011_0;
      patterns[10677] = 25'b00101001_10110011_11011100_0;
      patterns[10678] = 25'b00101001_10110100_11011101_0;
      patterns[10679] = 25'b00101001_10110101_11011110_0;
      patterns[10680] = 25'b00101001_10110110_11011111_0;
      patterns[10681] = 25'b00101001_10110111_11100000_0;
      patterns[10682] = 25'b00101001_10111000_11100001_0;
      patterns[10683] = 25'b00101001_10111001_11100010_0;
      patterns[10684] = 25'b00101001_10111010_11100011_0;
      patterns[10685] = 25'b00101001_10111011_11100100_0;
      patterns[10686] = 25'b00101001_10111100_11100101_0;
      patterns[10687] = 25'b00101001_10111101_11100110_0;
      patterns[10688] = 25'b00101001_10111110_11100111_0;
      patterns[10689] = 25'b00101001_10111111_11101000_0;
      patterns[10690] = 25'b00101001_11000000_11101001_0;
      patterns[10691] = 25'b00101001_11000001_11101010_0;
      patterns[10692] = 25'b00101001_11000010_11101011_0;
      patterns[10693] = 25'b00101001_11000011_11101100_0;
      patterns[10694] = 25'b00101001_11000100_11101101_0;
      patterns[10695] = 25'b00101001_11000101_11101110_0;
      patterns[10696] = 25'b00101001_11000110_11101111_0;
      patterns[10697] = 25'b00101001_11000111_11110000_0;
      patterns[10698] = 25'b00101001_11001000_11110001_0;
      patterns[10699] = 25'b00101001_11001001_11110010_0;
      patterns[10700] = 25'b00101001_11001010_11110011_0;
      patterns[10701] = 25'b00101001_11001011_11110100_0;
      patterns[10702] = 25'b00101001_11001100_11110101_0;
      patterns[10703] = 25'b00101001_11001101_11110110_0;
      patterns[10704] = 25'b00101001_11001110_11110111_0;
      patterns[10705] = 25'b00101001_11001111_11111000_0;
      patterns[10706] = 25'b00101001_11010000_11111001_0;
      patterns[10707] = 25'b00101001_11010001_11111010_0;
      patterns[10708] = 25'b00101001_11010010_11111011_0;
      patterns[10709] = 25'b00101001_11010011_11111100_0;
      patterns[10710] = 25'b00101001_11010100_11111101_0;
      patterns[10711] = 25'b00101001_11010101_11111110_0;
      patterns[10712] = 25'b00101001_11010110_11111111_0;
      patterns[10713] = 25'b00101001_11010111_00000000_1;
      patterns[10714] = 25'b00101001_11011000_00000001_1;
      patterns[10715] = 25'b00101001_11011001_00000010_1;
      patterns[10716] = 25'b00101001_11011010_00000011_1;
      patterns[10717] = 25'b00101001_11011011_00000100_1;
      patterns[10718] = 25'b00101001_11011100_00000101_1;
      patterns[10719] = 25'b00101001_11011101_00000110_1;
      patterns[10720] = 25'b00101001_11011110_00000111_1;
      patterns[10721] = 25'b00101001_11011111_00001000_1;
      patterns[10722] = 25'b00101001_11100000_00001001_1;
      patterns[10723] = 25'b00101001_11100001_00001010_1;
      patterns[10724] = 25'b00101001_11100010_00001011_1;
      patterns[10725] = 25'b00101001_11100011_00001100_1;
      patterns[10726] = 25'b00101001_11100100_00001101_1;
      patterns[10727] = 25'b00101001_11100101_00001110_1;
      patterns[10728] = 25'b00101001_11100110_00001111_1;
      patterns[10729] = 25'b00101001_11100111_00010000_1;
      patterns[10730] = 25'b00101001_11101000_00010001_1;
      patterns[10731] = 25'b00101001_11101001_00010010_1;
      patterns[10732] = 25'b00101001_11101010_00010011_1;
      patterns[10733] = 25'b00101001_11101011_00010100_1;
      patterns[10734] = 25'b00101001_11101100_00010101_1;
      patterns[10735] = 25'b00101001_11101101_00010110_1;
      patterns[10736] = 25'b00101001_11101110_00010111_1;
      patterns[10737] = 25'b00101001_11101111_00011000_1;
      patterns[10738] = 25'b00101001_11110000_00011001_1;
      patterns[10739] = 25'b00101001_11110001_00011010_1;
      patterns[10740] = 25'b00101001_11110010_00011011_1;
      patterns[10741] = 25'b00101001_11110011_00011100_1;
      patterns[10742] = 25'b00101001_11110100_00011101_1;
      patterns[10743] = 25'b00101001_11110101_00011110_1;
      patterns[10744] = 25'b00101001_11110110_00011111_1;
      patterns[10745] = 25'b00101001_11110111_00100000_1;
      patterns[10746] = 25'b00101001_11111000_00100001_1;
      patterns[10747] = 25'b00101001_11111001_00100010_1;
      patterns[10748] = 25'b00101001_11111010_00100011_1;
      patterns[10749] = 25'b00101001_11111011_00100100_1;
      patterns[10750] = 25'b00101001_11111100_00100101_1;
      patterns[10751] = 25'b00101001_11111101_00100110_1;
      patterns[10752] = 25'b00101001_11111110_00100111_1;
      patterns[10753] = 25'b00101001_11111111_00101000_1;
      patterns[10754] = 25'b00101010_00000000_00101010_0;
      patterns[10755] = 25'b00101010_00000001_00101011_0;
      patterns[10756] = 25'b00101010_00000010_00101100_0;
      patterns[10757] = 25'b00101010_00000011_00101101_0;
      patterns[10758] = 25'b00101010_00000100_00101110_0;
      patterns[10759] = 25'b00101010_00000101_00101111_0;
      patterns[10760] = 25'b00101010_00000110_00110000_0;
      patterns[10761] = 25'b00101010_00000111_00110001_0;
      patterns[10762] = 25'b00101010_00001000_00110010_0;
      patterns[10763] = 25'b00101010_00001001_00110011_0;
      patterns[10764] = 25'b00101010_00001010_00110100_0;
      patterns[10765] = 25'b00101010_00001011_00110101_0;
      patterns[10766] = 25'b00101010_00001100_00110110_0;
      patterns[10767] = 25'b00101010_00001101_00110111_0;
      patterns[10768] = 25'b00101010_00001110_00111000_0;
      patterns[10769] = 25'b00101010_00001111_00111001_0;
      patterns[10770] = 25'b00101010_00010000_00111010_0;
      patterns[10771] = 25'b00101010_00010001_00111011_0;
      patterns[10772] = 25'b00101010_00010010_00111100_0;
      patterns[10773] = 25'b00101010_00010011_00111101_0;
      patterns[10774] = 25'b00101010_00010100_00111110_0;
      patterns[10775] = 25'b00101010_00010101_00111111_0;
      patterns[10776] = 25'b00101010_00010110_01000000_0;
      patterns[10777] = 25'b00101010_00010111_01000001_0;
      patterns[10778] = 25'b00101010_00011000_01000010_0;
      patterns[10779] = 25'b00101010_00011001_01000011_0;
      patterns[10780] = 25'b00101010_00011010_01000100_0;
      patterns[10781] = 25'b00101010_00011011_01000101_0;
      patterns[10782] = 25'b00101010_00011100_01000110_0;
      patterns[10783] = 25'b00101010_00011101_01000111_0;
      patterns[10784] = 25'b00101010_00011110_01001000_0;
      patterns[10785] = 25'b00101010_00011111_01001001_0;
      patterns[10786] = 25'b00101010_00100000_01001010_0;
      patterns[10787] = 25'b00101010_00100001_01001011_0;
      patterns[10788] = 25'b00101010_00100010_01001100_0;
      patterns[10789] = 25'b00101010_00100011_01001101_0;
      patterns[10790] = 25'b00101010_00100100_01001110_0;
      patterns[10791] = 25'b00101010_00100101_01001111_0;
      patterns[10792] = 25'b00101010_00100110_01010000_0;
      patterns[10793] = 25'b00101010_00100111_01010001_0;
      patterns[10794] = 25'b00101010_00101000_01010010_0;
      patterns[10795] = 25'b00101010_00101001_01010011_0;
      patterns[10796] = 25'b00101010_00101010_01010100_0;
      patterns[10797] = 25'b00101010_00101011_01010101_0;
      patterns[10798] = 25'b00101010_00101100_01010110_0;
      patterns[10799] = 25'b00101010_00101101_01010111_0;
      patterns[10800] = 25'b00101010_00101110_01011000_0;
      patterns[10801] = 25'b00101010_00101111_01011001_0;
      patterns[10802] = 25'b00101010_00110000_01011010_0;
      patterns[10803] = 25'b00101010_00110001_01011011_0;
      patterns[10804] = 25'b00101010_00110010_01011100_0;
      patterns[10805] = 25'b00101010_00110011_01011101_0;
      patterns[10806] = 25'b00101010_00110100_01011110_0;
      patterns[10807] = 25'b00101010_00110101_01011111_0;
      patterns[10808] = 25'b00101010_00110110_01100000_0;
      patterns[10809] = 25'b00101010_00110111_01100001_0;
      patterns[10810] = 25'b00101010_00111000_01100010_0;
      patterns[10811] = 25'b00101010_00111001_01100011_0;
      patterns[10812] = 25'b00101010_00111010_01100100_0;
      patterns[10813] = 25'b00101010_00111011_01100101_0;
      patterns[10814] = 25'b00101010_00111100_01100110_0;
      patterns[10815] = 25'b00101010_00111101_01100111_0;
      patterns[10816] = 25'b00101010_00111110_01101000_0;
      patterns[10817] = 25'b00101010_00111111_01101001_0;
      patterns[10818] = 25'b00101010_01000000_01101010_0;
      patterns[10819] = 25'b00101010_01000001_01101011_0;
      patterns[10820] = 25'b00101010_01000010_01101100_0;
      patterns[10821] = 25'b00101010_01000011_01101101_0;
      patterns[10822] = 25'b00101010_01000100_01101110_0;
      patterns[10823] = 25'b00101010_01000101_01101111_0;
      patterns[10824] = 25'b00101010_01000110_01110000_0;
      patterns[10825] = 25'b00101010_01000111_01110001_0;
      patterns[10826] = 25'b00101010_01001000_01110010_0;
      patterns[10827] = 25'b00101010_01001001_01110011_0;
      patterns[10828] = 25'b00101010_01001010_01110100_0;
      patterns[10829] = 25'b00101010_01001011_01110101_0;
      patterns[10830] = 25'b00101010_01001100_01110110_0;
      patterns[10831] = 25'b00101010_01001101_01110111_0;
      patterns[10832] = 25'b00101010_01001110_01111000_0;
      patterns[10833] = 25'b00101010_01001111_01111001_0;
      patterns[10834] = 25'b00101010_01010000_01111010_0;
      patterns[10835] = 25'b00101010_01010001_01111011_0;
      patterns[10836] = 25'b00101010_01010010_01111100_0;
      patterns[10837] = 25'b00101010_01010011_01111101_0;
      patterns[10838] = 25'b00101010_01010100_01111110_0;
      patterns[10839] = 25'b00101010_01010101_01111111_0;
      patterns[10840] = 25'b00101010_01010110_10000000_0;
      patterns[10841] = 25'b00101010_01010111_10000001_0;
      patterns[10842] = 25'b00101010_01011000_10000010_0;
      patterns[10843] = 25'b00101010_01011001_10000011_0;
      patterns[10844] = 25'b00101010_01011010_10000100_0;
      patterns[10845] = 25'b00101010_01011011_10000101_0;
      patterns[10846] = 25'b00101010_01011100_10000110_0;
      patterns[10847] = 25'b00101010_01011101_10000111_0;
      patterns[10848] = 25'b00101010_01011110_10001000_0;
      patterns[10849] = 25'b00101010_01011111_10001001_0;
      patterns[10850] = 25'b00101010_01100000_10001010_0;
      patterns[10851] = 25'b00101010_01100001_10001011_0;
      patterns[10852] = 25'b00101010_01100010_10001100_0;
      patterns[10853] = 25'b00101010_01100011_10001101_0;
      patterns[10854] = 25'b00101010_01100100_10001110_0;
      patterns[10855] = 25'b00101010_01100101_10001111_0;
      patterns[10856] = 25'b00101010_01100110_10010000_0;
      patterns[10857] = 25'b00101010_01100111_10010001_0;
      patterns[10858] = 25'b00101010_01101000_10010010_0;
      patterns[10859] = 25'b00101010_01101001_10010011_0;
      patterns[10860] = 25'b00101010_01101010_10010100_0;
      patterns[10861] = 25'b00101010_01101011_10010101_0;
      patterns[10862] = 25'b00101010_01101100_10010110_0;
      patterns[10863] = 25'b00101010_01101101_10010111_0;
      patterns[10864] = 25'b00101010_01101110_10011000_0;
      patterns[10865] = 25'b00101010_01101111_10011001_0;
      patterns[10866] = 25'b00101010_01110000_10011010_0;
      patterns[10867] = 25'b00101010_01110001_10011011_0;
      patterns[10868] = 25'b00101010_01110010_10011100_0;
      patterns[10869] = 25'b00101010_01110011_10011101_0;
      patterns[10870] = 25'b00101010_01110100_10011110_0;
      patterns[10871] = 25'b00101010_01110101_10011111_0;
      patterns[10872] = 25'b00101010_01110110_10100000_0;
      patterns[10873] = 25'b00101010_01110111_10100001_0;
      patterns[10874] = 25'b00101010_01111000_10100010_0;
      patterns[10875] = 25'b00101010_01111001_10100011_0;
      patterns[10876] = 25'b00101010_01111010_10100100_0;
      patterns[10877] = 25'b00101010_01111011_10100101_0;
      patterns[10878] = 25'b00101010_01111100_10100110_0;
      patterns[10879] = 25'b00101010_01111101_10100111_0;
      patterns[10880] = 25'b00101010_01111110_10101000_0;
      patterns[10881] = 25'b00101010_01111111_10101001_0;
      patterns[10882] = 25'b00101010_10000000_10101010_0;
      patterns[10883] = 25'b00101010_10000001_10101011_0;
      patterns[10884] = 25'b00101010_10000010_10101100_0;
      patterns[10885] = 25'b00101010_10000011_10101101_0;
      patterns[10886] = 25'b00101010_10000100_10101110_0;
      patterns[10887] = 25'b00101010_10000101_10101111_0;
      patterns[10888] = 25'b00101010_10000110_10110000_0;
      patterns[10889] = 25'b00101010_10000111_10110001_0;
      patterns[10890] = 25'b00101010_10001000_10110010_0;
      patterns[10891] = 25'b00101010_10001001_10110011_0;
      patterns[10892] = 25'b00101010_10001010_10110100_0;
      patterns[10893] = 25'b00101010_10001011_10110101_0;
      patterns[10894] = 25'b00101010_10001100_10110110_0;
      patterns[10895] = 25'b00101010_10001101_10110111_0;
      patterns[10896] = 25'b00101010_10001110_10111000_0;
      patterns[10897] = 25'b00101010_10001111_10111001_0;
      patterns[10898] = 25'b00101010_10010000_10111010_0;
      patterns[10899] = 25'b00101010_10010001_10111011_0;
      patterns[10900] = 25'b00101010_10010010_10111100_0;
      patterns[10901] = 25'b00101010_10010011_10111101_0;
      patterns[10902] = 25'b00101010_10010100_10111110_0;
      patterns[10903] = 25'b00101010_10010101_10111111_0;
      patterns[10904] = 25'b00101010_10010110_11000000_0;
      patterns[10905] = 25'b00101010_10010111_11000001_0;
      patterns[10906] = 25'b00101010_10011000_11000010_0;
      patterns[10907] = 25'b00101010_10011001_11000011_0;
      patterns[10908] = 25'b00101010_10011010_11000100_0;
      patterns[10909] = 25'b00101010_10011011_11000101_0;
      patterns[10910] = 25'b00101010_10011100_11000110_0;
      patterns[10911] = 25'b00101010_10011101_11000111_0;
      patterns[10912] = 25'b00101010_10011110_11001000_0;
      patterns[10913] = 25'b00101010_10011111_11001001_0;
      patterns[10914] = 25'b00101010_10100000_11001010_0;
      patterns[10915] = 25'b00101010_10100001_11001011_0;
      patterns[10916] = 25'b00101010_10100010_11001100_0;
      patterns[10917] = 25'b00101010_10100011_11001101_0;
      patterns[10918] = 25'b00101010_10100100_11001110_0;
      patterns[10919] = 25'b00101010_10100101_11001111_0;
      patterns[10920] = 25'b00101010_10100110_11010000_0;
      patterns[10921] = 25'b00101010_10100111_11010001_0;
      patterns[10922] = 25'b00101010_10101000_11010010_0;
      patterns[10923] = 25'b00101010_10101001_11010011_0;
      patterns[10924] = 25'b00101010_10101010_11010100_0;
      patterns[10925] = 25'b00101010_10101011_11010101_0;
      patterns[10926] = 25'b00101010_10101100_11010110_0;
      patterns[10927] = 25'b00101010_10101101_11010111_0;
      patterns[10928] = 25'b00101010_10101110_11011000_0;
      patterns[10929] = 25'b00101010_10101111_11011001_0;
      patterns[10930] = 25'b00101010_10110000_11011010_0;
      patterns[10931] = 25'b00101010_10110001_11011011_0;
      patterns[10932] = 25'b00101010_10110010_11011100_0;
      patterns[10933] = 25'b00101010_10110011_11011101_0;
      patterns[10934] = 25'b00101010_10110100_11011110_0;
      patterns[10935] = 25'b00101010_10110101_11011111_0;
      patterns[10936] = 25'b00101010_10110110_11100000_0;
      patterns[10937] = 25'b00101010_10110111_11100001_0;
      patterns[10938] = 25'b00101010_10111000_11100010_0;
      patterns[10939] = 25'b00101010_10111001_11100011_0;
      patterns[10940] = 25'b00101010_10111010_11100100_0;
      patterns[10941] = 25'b00101010_10111011_11100101_0;
      patterns[10942] = 25'b00101010_10111100_11100110_0;
      patterns[10943] = 25'b00101010_10111101_11100111_0;
      patterns[10944] = 25'b00101010_10111110_11101000_0;
      patterns[10945] = 25'b00101010_10111111_11101001_0;
      patterns[10946] = 25'b00101010_11000000_11101010_0;
      patterns[10947] = 25'b00101010_11000001_11101011_0;
      patterns[10948] = 25'b00101010_11000010_11101100_0;
      patterns[10949] = 25'b00101010_11000011_11101101_0;
      patterns[10950] = 25'b00101010_11000100_11101110_0;
      patterns[10951] = 25'b00101010_11000101_11101111_0;
      patterns[10952] = 25'b00101010_11000110_11110000_0;
      patterns[10953] = 25'b00101010_11000111_11110001_0;
      patterns[10954] = 25'b00101010_11001000_11110010_0;
      patterns[10955] = 25'b00101010_11001001_11110011_0;
      patterns[10956] = 25'b00101010_11001010_11110100_0;
      patterns[10957] = 25'b00101010_11001011_11110101_0;
      patterns[10958] = 25'b00101010_11001100_11110110_0;
      patterns[10959] = 25'b00101010_11001101_11110111_0;
      patterns[10960] = 25'b00101010_11001110_11111000_0;
      patterns[10961] = 25'b00101010_11001111_11111001_0;
      patterns[10962] = 25'b00101010_11010000_11111010_0;
      patterns[10963] = 25'b00101010_11010001_11111011_0;
      patterns[10964] = 25'b00101010_11010010_11111100_0;
      patterns[10965] = 25'b00101010_11010011_11111101_0;
      patterns[10966] = 25'b00101010_11010100_11111110_0;
      patterns[10967] = 25'b00101010_11010101_11111111_0;
      patterns[10968] = 25'b00101010_11010110_00000000_1;
      patterns[10969] = 25'b00101010_11010111_00000001_1;
      patterns[10970] = 25'b00101010_11011000_00000010_1;
      patterns[10971] = 25'b00101010_11011001_00000011_1;
      patterns[10972] = 25'b00101010_11011010_00000100_1;
      patterns[10973] = 25'b00101010_11011011_00000101_1;
      patterns[10974] = 25'b00101010_11011100_00000110_1;
      patterns[10975] = 25'b00101010_11011101_00000111_1;
      patterns[10976] = 25'b00101010_11011110_00001000_1;
      patterns[10977] = 25'b00101010_11011111_00001001_1;
      patterns[10978] = 25'b00101010_11100000_00001010_1;
      patterns[10979] = 25'b00101010_11100001_00001011_1;
      patterns[10980] = 25'b00101010_11100010_00001100_1;
      patterns[10981] = 25'b00101010_11100011_00001101_1;
      patterns[10982] = 25'b00101010_11100100_00001110_1;
      patterns[10983] = 25'b00101010_11100101_00001111_1;
      patterns[10984] = 25'b00101010_11100110_00010000_1;
      patterns[10985] = 25'b00101010_11100111_00010001_1;
      patterns[10986] = 25'b00101010_11101000_00010010_1;
      patterns[10987] = 25'b00101010_11101001_00010011_1;
      patterns[10988] = 25'b00101010_11101010_00010100_1;
      patterns[10989] = 25'b00101010_11101011_00010101_1;
      patterns[10990] = 25'b00101010_11101100_00010110_1;
      patterns[10991] = 25'b00101010_11101101_00010111_1;
      patterns[10992] = 25'b00101010_11101110_00011000_1;
      patterns[10993] = 25'b00101010_11101111_00011001_1;
      patterns[10994] = 25'b00101010_11110000_00011010_1;
      patterns[10995] = 25'b00101010_11110001_00011011_1;
      patterns[10996] = 25'b00101010_11110010_00011100_1;
      patterns[10997] = 25'b00101010_11110011_00011101_1;
      patterns[10998] = 25'b00101010_11110100_00011110_1;
      patterns[10999] = 25'b00101010_11110101_00011111_1;
      patterns[11000] = 25'b00101010_11110110_00100000_1;
      patterns[11001] = 25'b00101010_11110111_00100001_1;
      patterns[11002] = 25'b00101010_11111000_00100010_1;
      patterns[11003] = 25'b00101010_11111001_00100011_1;
      patterns[11004] = 25'b00101010_11111010_00100100_1;
      patterns[11005] = 25'b00101010_11111011_00100101_1;
      patterns[11006] = 25'b00101010_11111100_00100110_1;
      patterns[11007] = 25'b00101010_11111101_00100111_1;
      patterns[11008] = 25'b00101010_11111110_00101000_1;
      patterns[11009] = 25'b00101010_11111111_00101001_1;
      patterns[11010] = 25'b00101011_00000000_00101011_0;
      patterns[11011] = 25'b00101011_00000001_00101100_0;
      patterns[11012] = 25'b00101011_00000010_00101101_0;
      patterns[11013] = 25'b00101011_00000011_00101110_0;
      patterns[11014] = 25'b00101011_00000100_00101111_0;
      patterns[11015] = 25'b00101011_00000101_00110000_0;
      patterns[11016] = 25'b00101011_00000110_00110001_0;
      patterns[11017] = 25'b00101011_00000111_00110010_0;
      patterns[11018] = 25'b00101011_00001000_00110011_0;
      patterns[11019] = 25'b00101011_00001001_00110100_0;
      patterns[11020] = 25'b00101011_00001010_00110101_0;
      patterns[11021] = 25'b00101011_00001011_00110110_0;
      patterns[11022] = 25'b00101011_00001100_00110111_0;
      patterns[11023] = 25'b00101011_00001101_00111000_0;
      patterns[11024] = 25'b00101011_00001110_00111001_0;
      patterns[11025] = 25'b00101011_00001111_00111010_0;
      patterns[11026] = 25'b00101011_00010000_00111011_0;
      patterns[11027] = 25'b00101011_00010001_00111100_0;
      patterns[11028] = 25'b00101011_00010010_00111101_0;
      patterns[11029] = 25'b00101011_00010011_00111110_0;
      patterns[11030] = 25'b00101011_00010100_00111111_0;
      patterns[11031] = 25'b00101011_00010101_01000000_0;
      patterns[11032] = 25'b00101011_00010110_01000001_0;
      patterns[11033] = 25'b00101011_00010111_01000010_0;
      patterns[11034] = 25'b00101011_00011000_01000011_0;
      patterns[11035] = 25'b00101011_00011001_01000100_0;
      patterns[11036] = 25'b00101011_00011010_01000101_0;
      patterns[11037] = 25'b00101011_00011011_01000110_0;
      patterns[11038] = 25'b00101011_00011100_01000111_0;
      patterns[11039] = 25'b00101011_00011101_01001000_0;
      patterns[11040] = 25'b00101011_00011110_01001001_0;
      patterns[11041] = 25'b00101011_00011111_01001010_0;
      patterns[11042] = 25'b00101011_00100000_01001011_0;
      patterns[11043] = 25'b00101011_00100001_01001100_0;
      patterns[11044] = 25'b00101011_00100010_01001101_0;
      patterns[11045] = 25'b00101011_00100011_01001110_0;
      patterns[11046] = 25'b00101011_00100100_01001111_0;
      patterns[11047] = 25'b00101011_00100101_01010000_0;
      patterns[11048] = 25'b00101011_00100110_01010001_0;
      patterns[11049] = 25'b00101011_00100111_01010010_0;
      patterns[11050] = 25'b00101011_00101000_01010011_0;
      patterns[11051] = 25'b00101011_00101001_01010100_0;
      patterns[11052] = 25'b00101011_00101010_01010101_0;
      patterns[11053] = 25'b00101011_00101011_01010110_0;
      patterns[11054] = 25'b00101011_00101100_01010111_0;
      patterns[11055] = 25'b00101011_00101101_01011000_0;
      patterns[11056] = 25'b00101011_00101110_01011001_0;
      patterns[11057] = 25'b00101011_00101111_01011010_0;
      patterns[11058] = 25'b00101011_00110000_01011011_0;
      patterns[11059] = 25'b00101011_00110001_01011100_0;
      patterns[11060] = 25'b00101011_00110010_01011101_0;
      patterns[11061] = 25'b00101011_00110011_01011110_0;
      patterns[11062] = 25'b00101011_00110100_01011111_0;
      patterns[11063] = 25'b00101011_00110101_01100000_0;
      patterns[11064] = 25'b00101011_00110110_01100001_0;
      patterns[11065] = 25'b00101011_00110111_01100010_0;
      patterns[11066] = 25'b00101011_00111000_01100011_0;
      patterns[11067] = 25'b00101011_00111001_01100100_0;
      patterns[11068] = 25'b00101011_00111010_01100101_0;
      patterns[11069] = 25'b00101011_00111011_01100110_0;
      patterns[11070] = 25'b00101011_00111100_01100111_0;
      patterns[11071] = 25'b00101011_00111101_01101000_0;
      patterns[11072] = 25'b00101011_00111110_01101001_0;
      patterns[11073] = 25'b00101011_00111111_01101010_0;
      patterns[11074] = 25'b00101011_01000000_01101011_0;
      patterns[11075] = 25'b00101011_01000001_01101100_0;
      patterns[11076] = 25'b00101011_01000010_01101101_0;
      patterns[11077] = 25'b00101011_01000011_01101110_0;
      patterns[11078] = 25'b00101011_01000100_01101111_0;
      patterns[11079] = 25'b00101011_01000101_01110000_0;
      patterns[11080] = 25'b00101011_01000110_01110001_0;
      patterns[11081] = 25'b00101011_01000111_01110010_0;
      patterns[11082] = 25'b00101011_01001000_01110011_0;
      patterns[11083] = 25'b00101011_01001001_01110100_0;
      patterns[11084] = 25'b00101011_01001010_01110101_0;
      patterns[11085] = 25'b00101011_01001011_01110110_0;
      patterns[11086] = 25'b00101011_01001100_01110111_0;
      patterns[11087] = 25'b00101011_01001101_01111000_0;
      patterns[11088] = 25'b00101011_01001110_01111001_0;
      patterns[11089] = 25'b00101011_01001111_01111010_0;
      patterns[11090] = 25'b00101011_01010000_01111011_0;
      patterns[11091] = 25'b00101011_01010001_01111100_0;
      patterns[11092] = 25'b00101011_01010010_01111101_0;
      patterns[11093] = 25'b00101011_01010011_01111110_0;
      patterns[11094] = 25'b00101011_01010100_01111111_0;
      patterns[11095] = 25'b00101011_01010101_10000000_0;
      patterns[11096] = 25'b00101011_01010110_10000001_0;
      patterns[11097] = 25'b00101011_01010111_10000010_0;
      patterns[11098] = 25'b00101011_01011000_10000011_0;
      patterns[11099] = 25'b00101011_01011001_10000100_0;
      patterns[11100] = 25'b00101011_01011010_10000101_0;
      patterns[11101] = 25'b00101011_01011011_10000110_0;
      patterns[11102] = 25'b00101011_01011100_10000111_0;
      patterns[11103] = 25'b00101011_01011101_10001000_0;
      patterns[11104] = 25'b00101011_01011110_10001001_0;
      patterns[11105] = 25'b00101011_01011111_10001010_0;
      patterns[11106] = 25'b00101011_01100000_10001011_0;
      patterns[11107] = 25'b00101011_01100001_10001100_0;
      patterns[11108] = 25'b00101011_01100010_10001101_0;
      patterns[11109] = 25'b00101011_01100011_10001110_0;
      patterns[11110] = 25'b00101011_01100100_10001111_0;
      patterns[11111] = 25'b00101011_01100101_10010000_0;
      patterns[11112] = 25'b00101011_01100110_10010001_0;
      patterns[11113] = 25'b00101011_01100111_10010010_0;
      patterns[11114] = 25'b00101011_01101000_10010011_0;
      patterns[11115] = 25'b00101011_01101001_10010100_0;
      patterns[11116] = 25'b00101011_01101010_10010101_0;
      patterns[11117] = 25'b00101011_01101011_10010110_0;
      patterns[11118] = 25'b00101011_01101100_10010111_0;
      patterns[11119] = 25'b00101011_01101101_10011000_0;
      patterns[11120] = 25'b00101011_01101110_10011001_0;
      patterns[11121] = 25'b00101011_01101111_10011010_0;
      patterns[11122] = 25'b00101011_01110000_10011011_0;
      patterns[11123] = 25'b00101011_01110001_10011100_0;
      patterns[11124] = 25'b00101011_01110010_10011101_0;
      patterns[11125] = 25'b00101011_01110011_10011110_0;
      patterns[11126] = 25'b00101011_01110100_10011111_0;
      patterns[11127] = 25'b00101011_01110101_10100000_0;
      patterns[11128] = 25'b00101011_01110110_10100001_0;
      patterns[11129] = 25'b00101011_01110111_10100010_0;
      patterns[11130] = 25'b00101011_01111000_10100011_0;
      patterns[11131] = 25'b00101011_01111001_10100100_0;
      patterns[11132] = 25'b00101011_01111010_10100101_0;
      patterns[11133] = 25'b00101011_01111011_10100110_0;
      patterns[11134] = 25'b00101011_01111100_10100111_0;
      patterns[11135] = 25'b00101011_01111101_10101000_0;
      patterns[11136] = 25'b00101011_01111110_10101001_0;
      patterns[11137] = 25'b00101011_01111111_10101010_0;
      patterns[11138] = 25'b00101011_10000000_10101011_0;
      patterns[11139] = 25'b00101011_10000001_10101100_0;
      patterns[11140] = 25'b00101011_10000010_10101101_0;
      patterns[11141] = 25'b00101011_10000011_10101110_0;
      patterns[11142] = 25'b00101011_10000100_10101111_0;
      patterns[11143] = 25'b00101011_10000101_10110000_0;
      patterns[11144] = 25'b00101011_10000110_10110001_0;
      patterns[11145] = 25'b00101011_10000111_10110010_0;
      patterns[11146] = 25'b00101011_10001000_10110011_0;
      patterns[11147] = 25'b00101011_10001001_10110100_0;
      patterns[11148] = 25'b00101011_10001010_10110101_0;
      patterns[11149] = 25'b00101011_10001011_10110110_0;
      patterns[11150] = 25'b00101011_10001100_10110111_0;
      patterns[11151] = 25'b00101011_10001101_10111000_0;
      patterns[11152] = 25'b00101011_10001110_10111001_0;
      patterns[11153] = 25'b00101011_10001111_10111010_0;
      patterns[11154] = 25'b00101011_10010000_10111011_0;
      patterns[11155] = 25'b00101011_10010001_10111100_0;
      patterns[11156] = 25'b00101011_10010010_10111101_0;
      patterns[11157] = 25'b00101011_10010011_10111110_0;
      patterns[11158] = 25'b00101011_10010100_10111111_0;
      patterns[11159] = 25'b00101011_10010101_11000000_0;
      patterns[11160] = 25'b00101011_10010110_11000001_0;
      patterns[11161] = 25'b00101011_10010111_11000010_0;
      patterns[11162] = 25'b00101011_10011000_11000011_0;
      patterns[11163] = 25'b00101011_10011001_11000100_0;
      patterns[11164] = 25'b00101011_10011010_11000101_0;
      patterns[11165] = 25'b00101011_10011011_11000110_0;
      patterns[11166] = 25'b00101011_10011100_11000111_0;
      patterns[11167] = 25'b00101011_10011101_11001000_0;
      patterns[11168] = 25'b00101011_10011110_11001001_0;
      patterns[11169] = 25'b00101011_10011111_11001010_0;
      patterns[11170] = 25'b00101011_10100000_11001011_0;
      patterns[11171] = 25'b00101011_10100001_11001100_0;
      patterns[11172] = 25'b00101011_10100010_11001101_0;
      patterns[11173] = 25'b00101011_10100011_11001110_0;
      patterns[11174] = 25'b00101011_10100100_11001111_0;
      patterns[11175] = 25'b00101011_10100101_11010000_0;
      patterns[11176] = 25'b00101011_10100110_11010001_0;
      patterns[11177] = 25'b00101011_10100111_11010010_0;
      patterns[11178] = 25'b00101011_10101000_11010011_0;
      patterns[11179] = 25'b00101011_10101001_11010100_0;
      patterns[11180] = 25'b00101011_10101010_11010101_0;
      patterns[11181] = 25'b00101011_10101011_11010110_0;
      patterns[11182] = 25'b00101011_10101100_11010111_0;
      patterns[11183] = 25'b00101011_10101101_11011000_0;
      patterns[11184] = 25'b00101011_10101110_11011001_0;
      patterns[11185] = 25'b00101011_10101111_11011010_0;
      patterns[11186] = 25'b00101011_10110000_11011011_0;
      patterns[11187] = 25'b00101011_10110001_11011100_0;
      patterns[11188] = 25'b00101011_10110010_11011101_0;
      patterns[11189] = 25'b00101011_10110011_11011110_0;
      patterns[11190] = 25'b00101011_10110100_11011111_0;
      patterns[11191] = 25'b00101011_10110101_11100000_0;
      patterns[11192] = 25'b00101011_10110110_11100001_0;
      patterns[11193] = 25'b00101011_10110111_11100010_0;
      patterns[11194] = 25'b00101011_10111000_11100011_0;
      patterns[11195] = 25'b00101011_10111001_11100100_0;
      patterns[11196] = 25'b00101011_10111010_11100101_0;
      patterns[11197] = 25'b00101011_10111011_11100110_0;
      patterns[11198] = 25'b00101011_10111100_11100111_0;
      patterns[11199] = 25'b00101011_10111101_11101000_0;
      patterns[11200] = 25'b00101011_10111110_11101001_0;
      patterns[11201] = 25'b00101011_10111111_11101010_0;
      patterns[11202] = 25'b00101011_11000000_11101011_0;
      patterns[11203] = 25'b00101011_11000001_11101100_0;
      patterns[11204] = 25'b00101011_11000010_11101101_0;
      patterns[11205] = 25'b00101011_11000011_11101110_0;
      patterns[11206] = 25'b00101011_11000100_11101111_0;
      patterns[11207] = 25'b00101011_11000101_11110000_0;
      patterns[11208] = 25'b00101011_11000110_11110001_0;
      patterns[11209] = 25'b00101011_11000111_11110010_0;
      patterns[11210] = 25'b00101011_11001000_11110011_0;
      patterns[11211] = 25'b00101011_11001001_11110100_0;
      patterns[11212] = 25'b00101011_11001010_11110101_0;
      patterns[11213] = 25'b00101011_11001011_11110110_0;
      patterns[11214] = 25'b00101011_11001100_11110111_0;
      patterns[11215] = 25'b00101011_11001101_11111000_0;
      patterns[11216] = 25'b00101011_11001110_11111001_0;
      patterns[11217] = 25'b00101011_11001111_11111010_0;
      patterns[11218] = 25'b00101011_11010000_11111011_0;
      patterns[11219] = 25'b00101011_11010001_11111100_0;
      patterns[11220] = 25'b00101011_11010010_11111101_0;
      patterns[11221] = 25'b00101011_11010011_11111110_0;
      patterns[11222] = 25'b00101011_11010100_11111111_0;
      patterns[11223] = 25'b00101011_11010101_00000000_1;
      patterns[11224] = 25'b00101011_11010110_00000001_1;
      patterns[11225] = 25'b00101011_11010111_00000010_1;
      patterns[11226] = 25'b00101011_11011000_00000011_1;
      patterns[11227] = 25'b00101011_11011001_00000100_1;
      patterns[11228] = 25'b00101011_11011010_00000101_1;
      patterns[11229] = 25'b00101011_11011011_00000110_1;
      patterns[11230] = 25'b00101011_11011100_00000111_1;
      patterns[11231] = 25'b00101011_11011101_00001000_1;
      patterns[11232] = 25'b00101011_11011110_00001001_1;
      patterns[11233] = 25'b00101011_11011111_00001010_1;
      patterns[11234] = 25'b00101011_11100000_00001011_1;
      patterns[11235] = 25'b00101011_11100001_00001100_1;
      patterns[11236] = 25'b00101011_11100010_00001101_1;
      patterns[11237] = 25'b00101011_11100011_00001110_1;
      patterns[11238] = 25'b00101011_11100100_00001111_1;
      patterns[11239] = 25'b00101011_11100101_00010000_1;
      patterns[11240] = 25'b00101011_11100110_00010001_1;
      patterns[11241] = 25'b00101011_11100111_00010010_1;
      patterns[11242] = 25'b00101011_11101000_00010011_1;
      patterns[11243] = 25'b00101011_11101001_00010100_1;
      patterns[11244] = 25'b00101011_11101010_00010101_1;
      patterns[11245] = 25'b00101011_11101011_00010110_1;
      patterns[11246] = 25'b00101011_11101100_00010111_1;
      patterns[11247] = 25'b00101011_11101101_00011000_1;
      patterns[11248] = 25'b00101011_11101110_00011001_1;
      patterns[11249] = 25'b00101011_11101111_00011010_1;
      patterns[11250] = 25'b00101011_11110000_00011011_1;
      patterns[11251] = 25'b00101011_11110001_00011100_1;
      patterns[11252] = 25'b00101011_11110010_00011101_1;
      patterns[11253] = 25'b00101011_11110011_00011110_1;
      patterns[11254] = 25'b00101011_11110100_00011111_1;
      patterns[11255] = 25'b00101011_11110101_00100000_1;
      patterns[11256] = 25'b00101011_11110110_00100001_1;
      patterns[11257] = 25'b00101011_11110111_00100010_1;
      patterns[11258] = 25'b00101011_11111000_00100011_1;
      patterns[11259] = 25'b00101011_11111001_00100100_1;
      patterns[11260] = 25'b00101011_11111010_00100101_1;
      patterns[11261] = 25'b00101011_11111011_00100110_1;
      patterns[11262] = 25'b00101011_11111100_00100111_1;
      patterns[11263] = 25'b00101011_11111101_00101000_1;
      patterns[11264] = 25'b00101011_11111110_00101001_1;
      patterns[11265] = 25'b00101011_11111111_00101010_1;
      patterns[11266] = 25'b00101100_00000000_00101100_0;
      patterns[11267] = 25'b00101100_00000001_00101101_0;
      patterns[11268] = 25'b00101100_00000010_00101110_0;
      patterns[11269] = 25'b00101100_00000011_00101111_0;
      patterns[11270] = 25'b00101100_00000100_00110000_0;
      patterns[11271] = 25'b00101100_00000101_00110001_0;
      patterns[11272] = 25'b00101100_00000110_00110010_0;
      patterns[11273] = 25'b00101100_00000111_00110011_0;
      patterns[11274] = 25'b00101100_00001000_00110100_0;
      patterns[11275] = 25'b00101100_00001001_00110101_0;
      patterns[11276] = 25'b00101100_00001010_00110110_0;
      patterns[11277] = 25'b00101100_00001011_00110111_0;
      patterns[11278] = 25'b00101100_00001100_00111000_0;
      patterns[11279] = 25'b00101100_00001101_00111001_0;
      patterns[11280] = 25'b00101100_00001110_00111010_0;
      patterns[11281] = 25'b00101100_00001111_00111011_0;
      patterns[11282] = 25'b00101100_00010000_00111100_0;
      patterns[11283] = 25'b00101100_00010001_00111101_0;
      patterns[11284] = 25'b00101100_00010010_00111110_0;
      patterns[11285] = 25'b00101100_00010011_00111111_0;
      patterns[11286] = 25'b00101100_00010100_01000000_0;
      patterns[11287] = 25'b00101100_00010101_01000001_0;
      patterns[11288] = 25'b00101100_00010110_01000010_0;
      patterns[11289] = 25'b00101100_00010111_01000011_0;
      patterns[11290] = 25'b00101100_00011000_01000100_0;
      patterns[11291] = 25'b00101100_00011001_01000101_0;
      patterns[11292] = 25'b00101100_00011010_01000110_0;
      patterns[11293] = 25'b00101100_00011011_01000111_0;
      patterns[11294] = 25'b00101100_00011100_01001000_0;
      patterns[11295] = 25'b00101100_00011101_01001001_0;
      patterns[11296] = 25'b00101100_00011110_01001010_0;
      patterns[11297] = 25'b00101100_00011111_01001011_0;
      patterns[11298] = 25'b00101100_00100000_01001100_0;
      patterns[11299] = 25'b00101100_00100001_01001101_0;
      patterns[11300] = 25'b00101100_00100010_01001110_0;
      patterns[11301] = 25'b00101100_00100011_01001111_0;
      patterns[11302] = 25'b00101100_00100100_01010000_0;
      patterns[11303] = 25'b00101100_00100101_01010001_0;
      patterns[11304] = 25'b00101100_00100110_01010010_0;
      patterns[11305] = 25'b00101100_00100111_01010011_0;
      patterns[11306] = 25'b00101100_00101000_01010100_0;
      patterns[11307] = 25'b00101100_00101001_01010101_0;
      patterns[11308] = 25'b00101100_00101010_01010110_0;
      patterns[11309] = 25'b00101100_00101011_01010111_0;
      patterns[11310] = 25'b00101100_00101100_01011000_0;
      patterns[11311] = 25'b00101100_00101101_01011001_0;
      patterns[11312] = 25'b00101100_00101110_01011010_0;
      patterns[11313] = 25'b00101100_00101111_01011011_0;
      patterns[11314] = 25'b00101100_00110000_01011100_0;
      patterns[11315] = 25'b00101100_00110001_01011101_0;
      patterns[11316] = 25'b00101100_00110010_01011110_0;
      patterns[11317] = 25'b00101100_00110011_01011111_0;
      patterns[11318] = 25'b00101100_00110100_01100000_0;
      patterns[11319] = 25'b00101100_00110101_01100001_0;
      patterns[11320] = 25'b00101100_00110110_01100010_0;
      patterns[11321] = 25'b00101100_00110111_01100011_0;
      patterns[11322] = 25'b00101100_00111000_01100100_0;
      patterns[11323] = 25'b00101100_00111001_01100101_0;
      patterns[11324] = 25'b00101100_00111010_01100110_0;
      patterns[11325] = 25'b00101100_00111011_01100111_0;
      patterns[11326] = 25'b00101100_00111100_01101000_0;
      patterns[11327] = 25'b00101100_00111101_01101001_0;
      patterns[11328] = 25'b00101100_00111110_01101010_0;
      patterns[11329] = 25'b00101100_00111111_01101011_0;
      patterns[11330] = 25'b00101100_01000000_01101100_0;
      patterns[11331] = 25'b00101100_01000001_01101101_0;
      patterns[11332] = 25'b00101100_01000010_01101110_0;
      patterns[11333] = 25'b00101100_01000011_01101111_0;
      patterns[11334] = 25'b00101100_01000100_01110000_0;
      patterns[11335] = 25'b00101100_01000101_01110001_0;
      patterns[11336] = 25'b00101100_01000110_01110010_0;
      patterns[11337] = 25'b00101100_01000111_01110011_0;
      patterns[11338] = 25'b00101100_01001000_01110100_0;
      patterns[11339] = 25'b00101100_01001001_01110101_0;
      patterns[11340] = 25'b00101100_01001010_01110110_0;
      patterns[11341] = 25'b00101100_01001011_01110111_0;
      patterns[11342] = 25'b00101100_01001100_01111000_0;
      patterns[11343] = 25'b00101100_01001101_01111001_0;
      patterns[11344] = 25'b00101100_01001110_01111010_0;
      patterns[11345] = 25'b00101100_01001111_01111011_0;
      patterns[11346] = 25'b00101100_01010000_01111100_0;
      patterns[11347] = 25'b00101100_01010001_01111101_0;
      patterns[11348] = 25'b00101100_01010010_01111110_0;
      patterns[11349] = 25'b00101100_01010011_01111111_0;
      patterns[11350] = 25'b00101100_01010100_10000000_0;
      patterns[11351] = 25'b00101100_01010101_10000001_0;
      patterns[11352] = 25'b00101100_01010110_10000010_0;
      patterns[11353] = 25'b00101100_01010111_10000011_0;
      patterns[11354] = 25'b00101100_01011000_10000100_0;
      patterns[11355] = 25'b00101100_01011001_10000101_0;
      patterns[11356] = 25'b00101100_01011010_10000110_0;
      patterns[11357] = 25'b00101100_01011011_10000111_0;
      patterns[11358] = 25'b00101100_01011100_10001000_0;
      patterns[11359] = 25'b00101100_01011101_10001001_0;
      patterns[11360] = 25'b00101100_01011110_10001010_0;
      patterns[11361] = 25'b00101100_01011111_10001011_0;
      patterns[11362] = 25'b00101100_01100000_10001100_0;
      patterns[11363] = 25'b00101100_01100001_10001101_0;
      patterns[11364] = 25'b00101100_01100010_10001110_0;
      patterns[11365] = 25'b00101100_01100011_10001111_0;
      patterns[11366] = 25'b00101100_01100100_10010000_0;
      patterns[11367] = 25'b00101100_01100101_10010001_0;
      patterns[11368] = 25'b00101100_01100110_10010010_0;
      patterns[11369] = 25'b00101100_01100111_10010011_0;
      patterns[11370] = 25'b00101100_01101000_10010100_0;
      patterns[11371] = 25'b00101100_01101001_10010101_0;
      patterns[11372] = 25'b00101100_01101010_10010110_0;
      patterns[11373] = 25'b00101100_01101011_10010111_0;
      patterns[11374] = 25'b00101100_01101100_10011000_0;
      patterns[11375] = 25'b00101100_01101101_10011001_0;
      patterns[11376] = 25'b00101100_01101110_10011010_0;
      patterns[11377] = 25'b00101100_01101111_10011011_0;
      patterns[11378] = 25'b00101100_01110000_10011100_0;
      patterns[11379] = 25'b00101100_01110001_10011101_0;
      patterns[11380] = 25'b00101100_01110010_10011110_0;
      patterns[11381] = 25'b00101100_01110011_10011111_0;
      patterns[11382] = 25'b00101100_01110100_10100000_0;
      patterns[11383] = 25'b00101100_01110101_10100001_0;
      patterns[11384] = 25'b00101100_01110110_10100010_0;
      patterns[11385] = 25'b00101100_01110111_10100011_0;
      patterns[11386] = 25'b00101100_01111000_10100100_0;
      patterns[11387] = 25'b00101100_01111001_10100101_0;
      patterns[11388] = 25'b00101100_01111010_10100110_0;
      patterns[11389] = 25'b00101100_01111011_10100111_0;
      patterns[11390] = 25'b00101100_01111100_10101000_0;
      patterns[11391] = 25'b00101100_01111101_10101001_0;
      patterns[11392] = 25'b00101100_01111110_10101010_0;
      patterns[11393] = 25'b00101100_01111111_10101011_0;
      patterns[11394] = 25'b00101100_10000000_10101100_0;
      patterns[11395] = 25'b00101100_10000001_10101101_0;
      patterns[11396] = 25'b00101100_10000010_10101110_0;
      patterns[11397] = 25'b00101100_10000011_10101111_0;
      patterns[11398] = 25'b00101100_10000100_10110000_0;
      patterns[11399] = 25'b00101100_10000101_10110001_0;
      patterns[11400] = 25'b00101100_10000110_10110010_0;
      patterns[11401] = 25'b00101100_10000111_10110011_0;
      patterns[11402] = 25'b00101100_10001000_10110100_0;
      patterns[11403] = 25'b00101100_10001001_10110101_0;
      patterns[11404] = 25'b00101100_10001010_10110110_0;
      patterns[11405] = 25'b00101100_10001011_10110111_0;
      patterns[11406] = 25'b00101100_10001100_10111000_0;
      patterns[11407] = 25'b00101100_10001101_10111001_0;
      patterns[11408] = 25'b00101100_10001110_10111010_0;
      patterns[11409] = 25'b00101100_10001111_10111011_0;
      patterns[11410] = 25'b00101100_10010000_10111100_0;
      patterns[11411] = 25'b00101100_10010001_10111101_0;
      patterns[11412] = 25'b00101100_10010010_10111110_0;
      patterns[11413] = 25'b00101100_10010011_10111111_0;
      patterns[11414] = 25'b00101100_10010100_11000000_0;
      patterns[11415] = 25'b00101100_10010101_11000001_0;
      patterns[11416] = 25'b00101100_10010110_11000010_0;
      patterns[11417] = 25'b00101100_10010111_11000011_0;
      patterns[11418] = 25'b00101100_10011000_11000100_0;
      patterns[11419] = 25'b00101100_10011001_11000101_0;
      patterns[11420] = 25'b00101100_10011010_11000110_0;
      patterns[11421] = 25'b00101100_10011011_11000111_0;
      patterns[11422] = 25'b00101100_10011100_11001000_0;
      patterns[11423] = 25'b00101100_10011101_11001001_0;
      patterns[11424] = 25'b00101100_10011110_11001010_0;
      patterns[11425] = 25'b00101100_10011111_11001011_0;
      patterns[11426] = 25'b00101100_10100000_11001100_0;
      patterns[11427] = 25'b00101100_10100001_11001101_0;
      patterns[11428] = 25'b00101100_10100010_11001110_0;
      patterns[11429] = 25'b00101100_10100011_11001111_0;
      patterns[11430] = 25'b00101100_10100100_11010000_0;
      patterns[11431] = 25'b00101100_10100101_11010001_0;
      patterns[11432] = 25'b00101100_10100110_11010010_0;
      patterns[11433] = 25'b00101100_10100111_11010011_0;
      patterns[11434] = 25'b00101100_10101000_11010100_0;
      patterns[11435] = 25'b00101100_10101001_11010101_0;
      patterns[11436] = 25'b00101100_10101010_11010110_0;
      patterns[11437] = 25'b00101100_10101011_11010111_0;
      patterns[11438] = 25'b00101100_10101100_11011000_0;
      patterns[11439] = 25'b00101100_10101101_11011001_0;
      patterns[11440] = 25'b00101100_10101110_11011010_0;
      patterns[11441] = 25'b00101100_10101111_11011011_0;
      patterns[11442] = 25'b00101100_10110000_11011100_0;
      patterns[11443] = 25'b00101100_10110001_11011101_0;
      patterns[11444] = 25'b00101100_10110010_11011110_0;
      patterns[11445] = 25'b00101100_10110011_11011111_0;
      patterns[11446] = 25'b00101100_10110100_11100000_0;
      patterns[11447] = 25'b00101100_10110101_11100001_0;
      patterns[11448] = 25'b00101100_10110110_11100010_0;
      patterns[11449] = 25'b00101100_10110111_11100011_0;
      patterns[11450] = 25'b00101100_10111000_11100100_0;
      patterns[11451] = 25'b00101100_10111001_11100101_0;
      patterns[11452] = 25'b00101100_10111010_11100110_0;
      patterns[11453] = 25'b00101100_10111011_11100111_0;
      patterns[11454] = 25'b00101100_10111100_11101000_0;
      patterns[11455] = 25'b00101100_10111101_11101001_0;
      patterns[11456] = 25'b00101100_10111110_11101010_0;
      patterns[11457] = 25'b00101100_10111111_11101011_0;
      patterns[11458] = 25'b00101100_11000000_11101100_0;
      patterns[11459] = 25'b00101100_11000001_11101101_0;
      patterns[11460] = 25'b00101100_11000010_11101110_0;
      patterns[11461] = 25'b00101100_11000011_11101111_0;
      patterns[11462] = 25'b00101100_11000100_11110000_0;
      patterns[11463] = 25'b00101100_11000101_11110001_0;
      patterns[11464] = 25'b00101100_11000110_11110010_0;
      patterns[11465] = 25'b00101100_11000111_11110011_0;
      patterns[11466] = 25'b00101100_11001000_11110100_0;
      patterns[11467] = 25'b00101100_11001001_11110101_0;
      patterns[11468] = 25'b00101100_11001010_11110110_0;
      patterns[11469] = 25'b00101100_11001011_11110111_0;
      patterns[11470] = 25'b00101100_11001100_11111000_0;
      patterns[11471] = 25'b00101100_11001101_11111001_0;
      patterns[11472] = 25'b00101100_11001110_11111010_0;
      patterns[11473] = 25'b00101100_11001111_11111011_0;
      patterns[11474] = 25'b00101100_11010000_11111100_0;
      patterns[11475] = 25'b00101100_11010001_11111101_0;
      patterns[11476] = 25'b00101100_11010010_11111110_0;
      patterns[11477] = 25'b00101100_11010011_11111111_0;
      patterns[11478] = 25'b00101100_11010100_00000000_1;
      patterns[11479] = 25'b00101100_11010101_00000001_1;
      patterns[11480] = 25'b00101100_11010110_00000010_1;
      patterns[11481] = 25'b00101100_11010111_00000011_1;
      patterns[11482] = 25'b00101100_11011000_00000100_1;
      patterns[11483] = 25'b00101100_11011001_00000101_1;
      patterns[11484] = 25'b00101100_11011010_00000110_1;
      patterns[11485] = 25'b00101100_11011011_00000111_1;
      patterns[11486] = 25'b00101100_11011100_00001000_1;
      patterns[11487] = 25'b00101100_11011101_00001001_1;
      patterns[11488] = 25'b00101100_11011110_00001010_1;
      patterns[11489] = 25'b00101100_11011111_00001011_1;
      patterns[11490] = 25'b00101100_11100000_00001100_1;
      patterns[11491] = 25'b00101100_11100001_00001101_1;
      patterns[11492] = 25'b00101100_11100010_00001110_1;
      patterns[11493] = 25'b00101100_11100011_00001111_1;
      patterns[11494] = 25'b00101100_11100100_00010000_1;
      patterns[11495] = 25'b00101100_11100101_00010001_1;
      patterns[11496] = 25'b00101100_11100110_00010010_1;
      patterns[11497] = 25'b00101100_11100111_00010011_1;
      patterns[11498] = 25'b00101100_11101000_00010100_1;
      patterns[11499] = 25'b00101100_11101001_00010101_1;
      patterns[11500] = 25'b00101100_11101010_00010110_1;
      patterns[11501] = 25'b00101100_11101011_00010111_1;
      patterns[11502] = 25'b00101100_11101100_00011000_1;
      patterns[11503] = 25'b00101100_11101101_00011001_1;
      patterns[11504] = 25'b00101100_11101110_00011010_1;
      patterns[11505] = 25'b00101100_11101111_00011011_1;
      patterns[11506] = 25'b00101100_11110000_00011100_1;
      patterns[11507] = 25'b00101100_11110001_00011101_1;
      patterns[11508] = 25'b00101100_11110010_00011110_1;
      patterns[11509] = 25'b00101100_11110011_00011111_1;
      patterns[11510] = 25'b00101100_11110100_00100000_1;
      patterns[11511] = 25'b00101100_11110101_00100001_1;
      patterns[11512] = 25'b00101100_11110110_00100010_1;
      patterns[11513] = 25'b00101100_11110111_00100011_1;
      patterns[11514] = 25'b00101100_11111000_00100100_1;
      patterns[11515] = 25'b00101100_11111001_00100101_1;
      patterns[11516] = 25'b00101100_11111010_00100110_1;
      patterns[11517] = 25'b00101100_11111011_00100111_1;
      patterns[11518] = 25'b00101100_11111100_00101000_1;
      patterns[11519] = 25'b00101100_11111101_00101001_1;
      patterns[11520] = 25'b00101100_11111110_00101010_1;
      patterns[11521] = 25'b00101100_11111111_00101011_1;
      patterns[11522] = 25'b00101101_00000000_00101101_0;
      patterns[11523] = 25'b00101101_00000001_00101110_0;
      patterns[11524] = 25'b00101101_00000010_00101111_0;
      patterns[11525] = 25'b00101101_00000011_00110000_0;
      patterns[11526] = 25'b00101101_00000100_00110001_0;
      patterns[11527] = 25'b00101101_00000101_00110010_0;
      patterns[11528] = 25'b00101101_00000110_00110011_0;
      patterns[11529] = 25'b00101101_00000111_00110100_0;
      patterns[11530] = 25'b00101101_00001000_00110101_0;
      patterns[11531] = 25'b00101101_00001001_00110110_0;
      patterns[11532] = 25'b00101101_00001010_00110111_0;
      patterns[11533] = 25'b00101101_00001011_00111000_0;
      patterns[11534] = 25'b00101101_00001100_00111001_0;
      patterns[11535] = 25'b00101101_00001101_00111010_0;
      patterns[11536] = 25'b00101101_00001110_00111011_0;
      patterns[11537] = 25'b00101101_00001111_00111100_0;
      patterns[11538] = 25'b00101101_00010000_00111101_0;
      patterns[11539] = 25'b00101101_00010001_00111110_0;
      patterns[11540] = 25'b00101101_00010010_00111111_0;
      patterns[11541] = 25'b00101101_00010011_01000000_0;
      patterns[11542] = 25'b00101101_00010100_01000001_0;
      patterns[11543] = 25'b00101101_00010101_01000010_0;
      patterns[11544] = 25'b00101101_00010110_01000011_0;
      patterns[11545] = 25'b00101101_00010111_01000100_0;
      patterns[11546] = 25'b00101101_00011000_01000101_0;
      patterns[11547] = 25'b00101101_00011001_01000110_0;
      patterns[11548] = 25'b00101101_00011010_01000111_0;
      patterns[11549] = 25'b00101101_00011011_01001000_0;
      patterns[11550] = 25'b00101101_00011100_01001001_0;
      patterns[11551] = 25'b00101101_00011101_01001010_0;
      patterns[11552] = 25'b00101101_00011110_01001011_0;
      patterns[11553] = 25'b00101101_00011111_01001100_0;
      patterns[11554] = 25'b00101101_00100000_01001101_0;
      patterns[11555] = 25'b00101101_00100001_01001110_0;
      patterns[11556] = 25'b00101101_00100010_01001111_0;
      patterns[11557] = 25'b00101101_00100011_01010000_0;
      patterns[11558] = 25'b00101101_00100100_01010001_0;
      patterns[11559] = 25'b00101101_00100101_01010010_0;
      patterns[11560] = 25'b00101101_00100110_01010011_0;
      patterns[11561] = 25'b00101101_00100111_01010100_0;
      patterns[11562] = 25'b00101101_00101000_01010101_0;
      patterns[11563] = 25'b00101101_00101001_01010110_0;
      patterns[11564] = 25'b00101101_00101010_01010111_0;
      patterns[11565] = 25'b00101101_00101011_01011000_0;
      patterns[11566] = 25'b00101101_00101100_01011001_0;
      patterns[11567] = 25'b00101101_00101101_01011010_0;
      patterns[11568] = 25'b00101101_00101110_01011011_0;
      patterns[11569] = 25'b00101101_00101111_01011100_0;
      patterns[11570] = 25'b00101101_00110000_01011101_0;
      patterns[11571] = 25'b00101101_00110001_01011110_0;
      patterns[11572] = 25'b00101101_00110010_01011111_0;
      patterns[11573] = 25'b00101101_00110011_01100000_0;
      patterns[11574] = 25'b00101101_00110100_01100001_0;
      patterns[11575] = 25'b00101101_00110101_01100010_0;
      patterns[11576] = 25'b00101101_00110110_01100011_0;
      patterns[11577] = 25'b00101101_00110111_01100100_0;
      patterns[11578] = 25'b00101101_00111000_01100101_0;
      patterns[11579] = 25'b00101101_00111001_01100110_0;
      patterns[11580] = 25'b00101101_00111010_01100111_0;
      patterns[11581] = 25'b00101101_00111011_01101000_0;
      patterns[11582] = 25'b00101101_00111100_01101001_0;
      patterns[11583] = 25'b00101101_00111101_01101010_0;
      patterns[11584] = 25'b00101101_00111110_01101011_0;
      patterns[11585] = 25'b00101101_00111111_01101100_0;
      patterns[11586] = 25'b00101101_01000000_01101101_0;
      patterns[11587] = 25'b00101101_01000001_01101110_0;
      patterns[11588] = 25'b00101101_01000010_01101111_0;
      patterns[11589] = 25'b00101101_01000011_01110000_0;
      patterns[11590] = 25'b00101101_01000100_01110001_0;
      patterns[11591] = 25'b00101101_01000101_01110010_0;
      patterns[11592] = 25'b00101101_01000110_01110011_0;
      patterns[11593] = 25'b00101101_01000111_01110100_0;
      patterns[11594] = 25'b00101101_01001000_01110101_0;
      patterns[11595] = 25'b00101101_01001001_01110110_0;
      patterns[11596] = 25'b00101101_01001010_01110111_0;
      patterns[11597] = 25'b00101101_01001011_01111000_0;
      patterns[11598] = 25'b00101101_01001100_01111001_0;
      patterns[11599] = 25'b00101101_01001101_01111010_0;
      patterns[11600] = 25'b00101101_01001110_01111011_0;
      patterns[11601] = 25'b00101101_01001111_01111100_0;
      patterns[11602] = 25'b00101101_01010000_01111101_0;
      patterns[11603] = 25'b00101101_01010001_01111110_0;
      patterns[11604] = 25'b00101101_01010010_01111111_0;
      patterns[11605] = 25'b00101101_01010011_10000000_0;
      patterns[11606] = 25'b00101101_01010100_10000001_0;
      patterns[11607] = 25'b00101101_01010101_10000010_0;
      patterns[11608] = 25'b00101101_01010110_10000011_0;
      patterns[11609] = 25'b00101101_01010111_10000100_0;
      patterns[11610] = 25'b00101101_01011000_10000101_0;
      patterns[11611] = 25'b00101101_01011001_10000110_0;
      patterns[11612] = 25'b00101101_01011010_10000111_0;
      patterns[11613] = 25'b00101101_01011011_10001000_0;
      patterns[11614] = 25'b00101101_01011100_10001001_0;
      patterns[11615] = 25'b00101101_01011101_10001010_0;
      patterns[11616] = 25'b00101101_01011110_10001011_0;
      patterns[11617] = 25'b00101101_01011111_10001100_0;
      patterns[11618] = 25'b00101101_01100000_10001101_0;
      patterns[11619] = 25'b00101101_01100001_10001110_0;
      patterns[11620] = 25'b00101101_01100010_10001111_0;
      patterns[11621] = 25'b00101101_01100011_10010000_0;
      patterns[11622] = 25'b00101101_01100100_10010001_0;
      patterns[11623] = 25'b00101101_01100101_10010010_0;
      patterns[11624] = 25'b00101101_01100110_10010011_0;
      patterns[11625] = 25'b00101101_01100111_10010100_0;
      patterns[11626] = 25'b00101101_01101000_10010101_0;
      patterns[11627] = 25'b00101101_01101001_10010110_0;
      patterns[11628] = 25'b00101101_01101010_10010111_0;
      patterns[11629] = 25'b00101101_01101011_10011000_0;
      patterns[11630] = 25'b00101101_01101100_10011001_0;
      patterns[11631] = 25'b00101101_01101101_10011010_0;
      patterns[11632] = 25'b00101101_01101110_10011011_0;
      patterns[11633] = 25'b00101101_01101111_10011100_0;
      patterns[11634] = 25'b00101101_01110000_10011101_0;
      patterns[11635] = 25'b00101101_01110001_10011110_0;
      patterns[11636] = 25'b00101101_01110010_10011111_0;
      patterns[11637] = 25'b00101101_01110011_10100000_0;
      patterns[11638] = 25'b00101101_01110100_10100001_0;
      patterns[11639] = 25'b00101101_01110101_10100010_0;
      patterns[11640] = 25'b00101101_01110110_10100011_0;
      patterns[11641] = 25'b00101101_01110111_10100100_0;
      patterns[11642] = 25'b00101101_01111000_10100101_0;
      patterns[11643] = 25'b00101101_01111001_10100110_0;
      patterns[11644] = 25'b00101101_01111010_10100111_0;
      patterns[11645] = 25'b00101101_01111011_10101000_0;
      patterns[11646] = 25'b00101101_01111100_10101001_0;
      patterns[11647] = 25'b00101101_01111101_10101010_0;
      patterns[11648] = 25'b00101101_01111110_10101011_0;
      patterns[11649] = 25'b00101101_01111111_10101100_0;
      patterns[11650] = 25'b00101101_10000000_10101101_0;
      patterns[11651] = 25'b00101101_10000001_10101110_0;
      patterns[11652] = 25'b00101101_10000010_10101111_0;
      patterns[11653] = 25'b00101101_10000011_10110000_0;
      patterns[11654] = 25'b00101101_10000100_10110001_0;
      patterns[11655] = 25'b00101101_10000101_10110010_0;
      patterns[11656] = 25'b00101101_10000110_10110011_0;
      patterns[11657] = 25'b00101101_10000111_10110100_0;
      patterns[11658] = 25'b00101101_10001000_10110101_0;
      patterns[11659] = 25'b00101101_10001001_10110110_0;
      patterns[11660] = 25'b00101101_10001010_10110111_0;
      patterns[11661] = 25'b00101101_10001011_10111000_0;
      patterns[11662] = 25'b00101101_10001100_10111001_0;
      patterns[11663] = 25'b00101101_10001101_10111010_0;
      patterns[11664] = 25'b00101101_10001110_10111011_0;
      patterns[11665] = 25'b00101101_10001111_10111100_0;
      patterns[11666] = 25'b00101101_10010000_10111101_0;
      patterns[11667] = 25'b00101101_10010001_10111110_0;
      patterns[11668] = 25'b00101101_10010010_10111111_0;
      patterns[11669] = 25'b00101101_10010011_11000000_0;
      patterns[11670] = 25'b00101101_10010100_11000001_0;
      patterns[11671] = 25'b00101101_10010101_11000010_0;
      patterns[11672] = 25'b00101101_10010110_11000011_0;
      patterns[11673] = 25'b00101101_10010111_11000100_0;
      patterns[11674] = 25'b00101101_10011000_11000101_0;
      patterns[11675] = 25'b00101101_10011001_11000110_0;
      patterns[11676] = 25'b00101101_10011010_11000111_0;
      patterns[11677] = 25'b00101101_10011011_11001000_0;
      patterns[11678] = 25'b00101101_10011100_11001001_0;
      patterns[11679] = 25'b00101101_10011101_11001010_0;
      patterns[11680] = 25'b00101101_10011110_11001011_0;
      patterns[11681] = 25'b00101101_10011111_11001100_0;
      patterns[11682] = 25'b00101101_10100000_11001101_0;
      patterns[11683] = 25'b00101101_10100001_11001110_0;
      patterns[11684] = 25'b00101101_10100010_11001111_0;
      patterns[11685] = 25'b00101101_10100011_11010000_0;
      patterns[11686] = 25'b00101101_10100100_11010001_0;
      patterns[11687] = 25'b00101101_10100101_11010010_0;
      patterns[11688] = 25'b00101101_10100110_11010011_0;
      patterns[11689] = 25'b00101101_10100111_11010100_0;
      patterns[11690] = 25'b00101101_10101000_11010101_0;
      patterns[11691] = 25'b00101101_10101001_11010110_0;
      patterns[11692] = 25'b00101101_10101010_11010111_0;
      patterns[11693] = 25'b00101101_10101011_11011000_0;
      patterns[11694] = 25'b00101101_10101100_11011001_0;
      patterns[11695] = 25'b00101101_10101101_11011010_0;
      patterns[11696] = 25'b00101101_10101110_11011011_0;
      patterns[11697] = 25'b00101101_10101111_11011100_0;
      patterns[11698] = 25'b00101101_10110000_11011101_0;
      patterns[11699] = 25'b00101101_10110001_11011110_0;
      patterns[11700] = 25'b00101101_10110010_11011111_0;
      patterns[11701] = 25'b00101101_10110011_11100000_0;
      patterns[11702] = 25'b00101101_10110100_11100001_0;
      patterns[11703] = 25'b00101101_10110101_11100010_0;
      patterns[11704] = 25'b00101101_10110110_11100011_0;
      patterns[11705] = 25'b00101101_10110111_11100100_0;
      patterns[11706] = 25'b00101101_10111000_11100101_0;
      patterns[11707] = 25'b00101101_10111001_11100110_0;
      patterns[11708] = 25'b00101101_10111010_11100111_0;
      patterns[11709] = 25'b00101101_10111011_11101000_0;
      patterns[11710] = 25'b00101101_10111100_11101001_0;
      patterns[11711] = 25'b00101101_10111101_11101010_0;
      patterns[11712] = 25'b00101101_10111110_11101011_0;
      patterns[11713] = 25'b00101101_10111111_11101100_0;
      patterns[11714] = 25'b00101101_11000000_11101101_0;
      patterns[11715] = 25'b00101101_11000001_11101110_0;
      patterns[11716] = 25'b00101101_11000010_11101111_0;
      patterns[11717] = 25'b00101101_11000011_11110000_0;
      patterns[11718] = 25'b00101101_11000100_11110001_0;
      patterns[11719] = 25'b00101101_11000101_11110010_0;
      patterns[11720] = 25'b00101101_11000110_11110011_0;
      patterns[11721] = 25'b00101101_11000111_11110100_0;
      patterns[11722] = 25'b00101101_11001000_11110101_0;
      patterns[11723] = 25'b00101101_11001001_11110110_0;
      patterns[11724] = 25'b00101101_11001010_11110111_0;
      patterns[11725] = 25'b00101101_11001011_11111000_0;
      patterns[11726] = 25'b00101101_11001100_11111001_0;
      patterns[11727] = 25'b00101101_11001101_11111010_0;
      patterns[11728] = 25'b00101101_11001110_11111011_0;
      patterns[11729] = 25'b00101101_11001111_11111100_0;
      patterns[11730] = 25'b00101101_11010000_11111101_0;
      patterns[11731] = 25'b00101101_11010001_11111110_0;
      patterns[11732] = 25'b00101101_11010010_11111111_0;
      patterns[11733] = 25'b00101101_11010011_00000000_1;
      patterns[11734] = 25'b00101101_11010100_00000001_1;
      patterns[11735] = 25'b00101101_11010101_00000010_1;
      patterns[11736] = 25'b00101101_11010110_00000011_1;
      patterns[11737] = 25'b00101101_11010111_00000100_1;
      patterns[11738] = 25'b00101101_11011000_00000101_1;
      patterns[11739] = 25'b00101101_11011001_00000110_1;
      patterns[11740] = 25'b00101101_11011010_00000111_1;
      patterns[11741] = 25'b00101101_11011011_00001000_1;
      patterns[11742] = 25'b00101101_11011100_00001001_1;
      patterns[11743] = 25'b00101101_11011101_00001010_1;
      patterns[11744] = 25'b00101101_11011110_00001011_1;
      patterns[11745] = 25'b00101101_11011111_00001100_1;
      patterns[11746] = 25'b00101101_11100000_00001101_1;
      patterns[11747] = 25'b00101101_11100001_00001110_1;
      patterns[11748] = 25'b00101101_11100010_00001111_1;
      patterns[11749] = 25'b00101101_11100011_00010000_1;
      patterns[11750] = 25'b00101101_11100100_00010001_1;
      patterns[11751] = 25'b00101101_11100101_00010010_1;
      patterns[11752] = 25'b00101101_11100110_00010011_1;
      patterns[11753] = 25'b00101101_11100111_00010100_1;
      patterns[11754] = 25'b00101101_11101000_00010101_1;
      patterns[11755] = 25'b00101101_11101001_00010110_1;
      patterns[11756] = 25'b00101101_11101010_00010111_1;
      patterns[11757] = 25'b00101101_11101011_00011000_1;
      patterns[11758] = 25'b00101101_11101100_00011001_1;
      patterns[11759] = 25'b00101101_11101101_00011010_1;
      patterns[11760] = 25'b00101101_11101110_00011011_1;
      patterns[11761] = 25'b00101101_11101111_00011100_1;
      patterns[11762] = 25'b00101101_11110000_00011101_1;
      patterns[11763] = 25'b00101101_11110001_00011110_1;
      patterns[11764] = 25'b00101101_11110010_00011111_1;
      patterns[11765] = 25'b00101101_11110011_00100000_1;
      patterns[11766] = 25'b00101101_11110100_00100001_1;
      patterns[11767] = 25'b00101101_11110101_00100010_1;
      patterns[11768] = 25'b00101101_11110110_00100011_1;
      patterns[11769] = 25'b00101101_11110111_00100100_1;
      patterns[11770] = 25'b00101101_11111000_00100101_1;
      patterns[11771] = 25'b00101101_11111001_00100110_1;
      patterns[11772] = 25'b00101101_11111010_00100111_1;
      patterns[11773] = 25'b00101101_11111011_00101000_1;
      patterns[11774] = 25'b00101101_11111100_00101001_1;
      patterns[11775] = 25'b00101101_11111101_00101010_1;
      patterns[11776] = 25'b00101101_11111110_00101011_1;
      patterns[11777] = 25'b00101101_11111111_00101100_1;
      patterns[11778] = 25'b00101110_00000000_00101110_0;
      patterns[11779] = 25'b00101110_00000001_00101111_0;
      patterns[11780] = 25'b00101110_00000010_00110000_0;
      patterns[11781] = 25'b00101110_00000011_00110001_0;
      patterns[11782] = 25'b00101110_00000100_00110010_0;
      patterns[11783] = 25'b00101110_00000101_00110011_0;
      patterns[11784] = 25'b00101110_00000110_00110100_0;
      patterns[11785] = 25'b00101110_00000111_00110101_0;
      patterns[11786] = 25'b00101110_00001000_00110110_0;
      patterns[11787] = 25'b00101110_00001001_00110111_0;
      patterns[11788] = 25'b00101110_00001010_00111000_0;
      patterns[11789] = 25'b00101110_00001011_00111001_0;
      patterns[11790] = 25'b00101110_00001100_00111010_0;
      patterns[11791] = 25'b00101110_00001101_00111011_0;
      patterns[11792] = 25'b00101110_00001110_00111100_0;
      patterns[11793] = 25'b00101110_00001111_00111101_0;
      patterns[11794] = 25'b00101110_00010000_00111110_0;
      patterns[11795] = 25'b00101110_00010001_00111111_0;
      patterns[11796] = 25'b00101110_00010010_01000000_0;
      patterns[11797] = 25'b00101110_00010011_01000001_0;
      patterns[11798] = 25'b00101110_00010100_01000010_0;
      patterns[11799] = 25'b00101110_00010101_01000011_0;
      patterns[11800] = 25'b00101110_00010110_01000100_0;
      patterns[11801] = 25'b00101110_00010111_01000101_0;
      patterns[11802] = 25'b00101110_00011000_01000110_0;
      patterns[11803] = 25'b00101110_00011001_01000111_0;
      patterns[11804] = 25'b00101110_00011010_01001000_0;
      patterns[11805] = 25'b00101110_00011011_01001001_0;
      patterns[11806] = 25'b00101110_00011100_01001010_0;
      patterns[11807] = 25'b00101110_00011101_01001011_0;
      patterns[11808] = 25'b00101110_00011110_01001100_0;
      patterns[11809] = 25'b00101110_00011111_01001101_0;
      patterns[11810] = 25'b00101110_00100000_01001110_0;
      patterns[11811] = 25'b00101110_00100001_01001111_0;
      patterns[11812] = 25'b00101110_00100010_01010000_0;
      patterns[11813] = 25'b00101110_00100011_01010001_0;
      patterns[11814] = 25'b00101110_00100100_01010010_0;
      patterns[11815] = 25'b00101110_00100101_01010011_0;
      patterns[11816] = 25'b00101110_00100110_01010100_0;
      patterns[11817] = 25'b00101110_00100111_01010101_0;
      patterns[11818] = 25'b00101110_00101000_01010110_0;
      patterns[11819] = 25'b00101110_00101001_01010111_0;
      patterns[11820] = 25'b00101110_00101010_01011000_0;
      patterns[11821] = 25'b00101110_00101011_01011001_0;
      patterns[11822] = 25'b00101110_00101100_01011010_0;
      patterns[11823] = 25'b00101110_00101101_01011011_0;
      patterns[11824] = 25'b00101110_00101110_01011100_0;
      patterns[11825] = 25'b00101110_00101111_01011101_0;
      patterns[11826] = 25'b00101110_00110000_01011110_0;
      patterns[11827] = 25'b00101110_00110001_01011111_0;
      patterns[11828] = 25'b00101110_00110010_01100000_0;
      patterns[11829] = 25'b00101110_00110011_01100001_0;
      patterns[11830] = 25'b00101110_00110100_01100010_0;
      patterns[11831] = 25'b00101110_00110101_01100011_0;
      patterns[11832] = 25'b00101110_00110110_01100100_0;
      patterns[11833] = 25'b00101110_00110111_01100101_0;
      patterns[11834] = 25'b00101110_00111000_01100110_0;
      patterns[11835] = 25'b00101110_00111001_01100111_0;
      patterns[11836] = 25'b00101110_00111010_01101000_0;
      patterns[11837] = 25'b00101110_00111011_01101001_0;
      patterns[11838] = 25'b00101110_00111100_01101010_0;
      patterns[11839] = 25'b00101110_00111101_01101011_0;
      patterns[11840] = 25'b00101110_00111110_01101100_0;
      patterns[11841] = 25'b00101110_00111111_01101101_0;
      patterns[11842] = 25'b00101110_01000000_01101110_0;
      patterns[11843] = 25'b00101110_01000001_01101111_0;
      patterns[11844] = 25'b00101110_01000010_01110000_0;
      patterns[11845] = 25'b00101110_01000011_01110001_0;
      patterns[11846] = 25'b00101110_01000100_01110010_0;
      patterns[11847] = 25'b00101110_01000101_01110011_0;
      patterns[11848] = 25'b00101110_01000110_01110100_0;
      patterns[11849] = 25'b00101110_01000111_01110101_0;
      patterns[11850] = 25'b00101110_01001000_01110110_0;
      patterns[11851] = 25'b00101110_01001001_01110111_0;
      patterns[11852] = 25'b00101110_01001010_01111000_0;
      patterns[11853] = 25'b00101110_01001011_01111001_0;
      patterns[11854] = 25'b00101110_01001100_01111010_0;
      patterns[11855] = 25'b00101110_01001101_01111011_0;
      patterns[11856] = 25'b00101110_01001110_01111100_0;
      patterns[11857] = 25'b00101110_01001111_01111101_0;
      patterns[11858] = 25'b00101110_01010000_01111110_0;
      patterns[11859] = 25'b00101110_01010001_01111111_0;
      patterns[11860] = 25'b00101110_01010010_10000000_0;
      patterns[11861] = 25'b00101110_01010011_10000001_0;
      patterns[11862] = 25'b00101110_01010100_10000010_0;
      patterns[11863] = 25'b00101110_01010101_10000011_0;
      patterns[11864] = 25'b00101110_01010110_10000100_0;
      patterns[11865] = 25'b00101110_01010111_10000101_0;
      patterns[11866] = 25'b00101110_01011000_10000110_0;
      patterns[11867] = 25'b00101110_01011001_10000111_0;
      patterns[11868] = 25'b00101110_01011010_10001000_0;
      patterns[11869] = 25'b00101110_01011011_10001001_0;
      patterns[11870] = 25'b00101110_01011100_10001010_0;
      patterns[11871] = 25'b00101110_01011101_10001011_0;
      patterns[11872] = 25'b00101110_01011110_10001100_0;
      patterns[11873] = 25'b00101110_01011111_10001101_0;
      patterns[11874] = 25'b00101110_01100000_10001110_0;
      patterns[11875] = 25'b00101110_01100001_10001111_0;
      patterns[11876] = 25'b00101110_01100010_10010000_0;
      patterns[11877] = 25'b00101110_01100011_10010001_0;
      patterns[11878] = 25'b00101110_01100100_10010010_0;
      patterns[11879] = 25'b00101110_01100101_10010011_0;
      patterns[11880] = 25'b00101110_01100110_10010100_0;
      patterns[11881] = 25'b00101110_01100111_10010101_0;
      patterns[11882] = 25'b00101110_01101000_10010110_0;
      patterns[11883] = 25'b00101110_01101001_10010111_0;
      patterns[11884] = 25'b00101110_01101010_10011000_0;
      patterns[11885] = 25'b00101110_01101011_10011001_0;
      patterns[11886] = 25'b00101110_01101100_10011010_0;
      patterns[11887] = 25'b00101110_01101101_10011011_0;
      patterns[11888] = 25'b00101110_01101110_10011100_0;
      patterns[11889] = 25'b00101110_01101111_10011101_0;
      patterns[11890] = 25'b00101110_01110000_10011110_0;
      patterns[11891] = 25'b00101110_01110001_10011111_0;
      patterns[11892] = 25'b00101110_01110010_10100000_0;
      patterns[11893] = 25'b00101110_01110011_10100001_0;
      patterns[11894] = 25'b00101110_01110100_10100010_0;
      patterns[11895] = 25'b00101110_01110101_10100011_0;
      patterns[11896] = 25'b00101110_01110110_10100100_0;
      patterns[11897] = 25'b00101110_01110111_10100101_0;
      patterns[11898] = 25'b00101110_01111000_10100110_0;
      patterns[11899] = 25'b00101110_01111001_10100111_0;
      patterns[11900] = 25'b00101110_01111010_10101000_0;
      patterns[11901] = 25'b00101110_01111011_10101001_0;
      patterns[11902] = 25'b00101110_01111100_10101010_0;
      patterns[11903] = 25'b00101110_01111101_10101011_0;
      patterns[11904] = 25'b00101110_01111110_10101100_0;
      patterns[11905] = 25'b00101110_01111111_10101101_0;
      patterns[11906] = 25'b00101110_10000000_10101110_0;
      patterns[11907] = 25'b00101110_10000001_10101111_0;
      patterns[11908] = 25'b00101110_10000010_10110000_0;
      patterns[11909] = 25'b00101110_10000011_10110001_0;
      patterns[11910] = 25'b00101110_10000100_10110010_0;
      patterns[11911] = 25'b00101110_10000101_10110011_0;
      patterns[11912] = 25'b00101110_10000110_10110100_0;
      patterns[11913] = 25'b00101110_10000111_10110101_0;
      patterns[11914] = 25'b00101110_10001000_10110110_0;
      patterns[11915] = 25'b00101110_10001001_10110111_0;
      patterns[11916] = 25'b00101110_10001010_10111000_0;
      patterns[11917] = 25'b00101110_10001011_10111001_0;
      patterns[11918] = 25'b00101110_10001100_10111010_0;
      patterns[11919] = 25'b00101110_10001101_10111011_0;
      patterns[11920] = 25'b00101110_10001110_10111100_0;
      patterns[11921] = 25'b00101110_10001111_10111101_0;
      patterns[11922] = 25'b00101110_10010000_10111110_0;
      patterns[11923] = 25'b00101110_10010001_10111111_0;
      patterns[11924] = 25'b00101110_10010010_11000000_0;
      patterns[11925] = 25'b00101110_10010011_11000001_0;
      patterns[11926] = 25'b00101110_10010100_11000010_0;
      patterns[11927] = 25'b00101110_10010101_11000011_0;
      patterns[11928] = 25'b00101110_10010110_11000100_0;
      patterns[11929] = 25'b00101110_10010111_11000101_0;
      patterns[11930] = 25'b00101110_10011000_11000110_0;
      patterns[11931] = 25'b00101110_10011001_11000111_0;
      patterns[11932] = 25'b00101110_10011010_11001000_0;
      patterns[11933] = 25'b00101110_10011011_11001001_0;
      patterns[11934] = 25'b00101110_10011100_11001010_0;
      patterns[11935] = 25'b00101110_10011101_11001011_0;
      patterns[11936] = 25'b00101110_10011110_11001100_0;
      patterns[11937] = 25'b00101110_10011111_11001101_0;
      patterns[11938] = 25'b00101110_10100000_11001110_0;
      patterns[11939] = 25'b00101110_10100001_11001111_0;
      patterns[11940] = 25'b00101110_10100010_11010000_0;
      patterns[11941] = 25'b00101110_10100011_11010001_0;
      patterns[11942] = 25'b00101110_10100100_11010010_0;
      patterns[11943] = 25'b00101110_10100101_11010011_0;
      patterns[11944] = 25'b00101110_10100110_11010100_0;
      patterns[11945] = 25'b00101110_10100111_11010101_0;
      patterns[11946] = 25'b00101110_10101000_11010110_0;
      patterns[11947] = 25'b00101110_10101001_11010111_0;
      patterns[11948] = 25'b00101110_10101010_11011000_0;
      patterns[11949] = 25'b00101110_10101011_11011001_0;
      patterns[11950] = 25'b00101110_10101100_11011010_0;
      patterns[11951] = 25'b00101110_10101101_11011011_0;
      patterns[11952] = 25'b00101110_10101110_11011100_0;
      patterns[11953] = 25'b00101110_10101111_11011101_0;
      patterns[11954] = 25'b00101110_10110000_11011110_0;
      patterns[11955] = 25'b00101110_10110001_11011111_0;
      patterns[11956] = 25'b00101110_10110010_11100000_0;
      patterns[11957] = 25'b00101110_10110011_11100001_0;
      patterns[11958] = 25'b00101110_10110100_11100010_0;
      patterns[11959] = 25'b00101110_10110101_11100011_0;
      patterns[11960] = 25'b00101110_10110110_11100100_0;
      patterns[11961] = 25'b00101110_10110111_11100101_0;
      patterns[11962] = 25'b00101110_10111000_11100110_0;
      patterns[11963] = 25'b00101110_10111001_11100111_0;
      patterns[11964] = 25'b00101110_10111010_11101000_0;
      patterns[11965] = 25'b00101110_10111011_11101001_0;
      patterns[11966] = 25'b00101110_10111100_11101010_0;
      patterns[11967] = 25'b00101110_10111101_11101011_0;
      patterns[11968] = 25'b00101110_10111110_11101100_0;
      patterns[11969] = 25'b00101110_10111111_11101101_0;
      patterns[11970] = 25'b00101110_11000000_11101110_0;
      patterns[11971] = 25'b00101110_11000001_11101111_0;
      patterns[11972] = 25'b00101110_11000010_11110000_0;
      patterns[11973] = 25'b00101110_11000011_11110001_0;
      patterns[11974] = 25'b00101110_11000100_11110010_0;
      patterns[11975] = 25'b00101110_11000101_11110011_0;
      patterns[11976] = 25'b00101110_11000110_11110100_0;
      patterns[11977] = 25'b00101110_11000111_11110101_0;
      patterns[11978] = 25'b00101110_11001000_11110110_0;
      patterns[11979] = 25'b00101110_11001001_11110111_0;
      patterns[11980] = 25'b00101110_11001010_11111000_0;
      patterns[11981] = 25'b00101110_11001011_11111001_0;
      patterns[11982] = 25'b00101110_11001100_11111010_0;
      patterns[11983] = 25'b00101110_11001101_11111011_0;
      patterns[11984] = 25'b00101110_11001110_11111100_0;
      patterns[11985] = 25'b00101110_11001111_11111101_0;
      patterns[11986] = 25'b00101110_11010000_11111110_0;
      patterns[11987] = 25'b00101110_11010001_11111111_0;
      patterns[11988] = 25'b00101110_11010010_00000000_1;
      patterns[11989] = 25'b00101110_11010011_00000001_1;
      patterns[11990] = 25'b00101110_11010100_00000010_1;
      patterns[11991] = 25'b00101110_11010101_00000011_1;
      patterns[11992] = 25'b00101110_11010110_00000100_1;
      patterns[11993] = 25'b00101110_11010111_00000101_1;
      patterns[11994] = 25'b00101110_11011000_00000110_1;
      patterns[11995] = 25'b00101110_11011001_00000111_1;
      patterns[11996] = 25'b00101110_11011010_00001000_1;
      patterns[11997] = 25'b00101110_11011011_00001001_1;
      patterns[11998] = 25'b00101110_11011100_00001010_1;
      patterns[11999] = 25'b00101110_11011101_00001011_1;
      patterns[12000] = 25'b00101110_11011110_00001100_1;
      patterns[12001] = 25'b00101110_11011111_00001101_1;
      patterns[12002] = 25'b00101110_11100000_00001110_1;
      patterns[12003] = 25'b00101110_11100001_00001111_1;
      patterns[12004] = 25'b00101110_11100010_00010000_1;
      patterns[12005] = 25'b00101110_11100011_00010001_1;
      patterns[12006] = 25'b00101110_11100100_00010010_1;
      patterns[12007] = 25'b00101110_11100101_00010011_1;
      patterns[12008] = 25'b00101110_11100110_00010100_1;
      patterns[12009] = 25'b00101110_11100111_00010101_1;
      patterns[12010] = 25'b00101110_11101000_00010110_1;
      patterns[12011] = 25'b00101110_11101001_00010111_1;
      patterns[12012] = 25'b00101110_11101010_00011000_1;
      patterns[12013] = 25'b00101110_11101011_00011001_1;
      patterns[12014] = 25'b00101110_11101100_00011010_1;
      patterns[12015] = 25'b00101110_11101101_00011011_1;
      patterns[12016] = 25'b00101110_11101110_00011100_1;
      patterns[12017] = 25'b00101110_11101111_00011101_1;
      patterns[12018] = 25'b00101110_11110000_00011110_1;
      patterns[12019] = 25'b00101110_11110001_00011111_1;
      patterns[12020] = 25'b00101110_11110010_00100000_1;
      patterns[12021] = 25'b00101110_11110011_00100001_1;
      patterns[12022] = 25'b00101110_11110100_00100010_1;
      patterns[12023] = 25'b00101110_11110101_00100011_1;
      patterns[12024] = 25'b00101110_11110110_00100100_1;
      patterns[12025] = 25'b00101110_11110111_00100101_1;
      patterns[12026] = 25'b00101110_11111000_00100110_1;
      patterns[12027] = 25'b00101110_11111001_00100111_1;
      patterns[12028] = 25'b00101110_11111010_00101000_1;
      patterns[12029] = 25'b00101110_11111011_00101001_1;
      patterns[12030] = 25'b00101110_11111100_00101010_1;
      patterns[12031] = 25'b00101110_11111101_00101011_1;
      patterns[12032] = 25'b00101110_11111110_00101100_1;
      patterns[12033] = 25'b00101110_11111111_00101101_1;
      patterns[12034] = 25'b00101111_00000000_00101111_0;
      patterns[12035] = 25'b00101111_00000001_00110000_0;
      patterns[12036] = 25'b00101111_00000010_00110001_0;
      patterns[12037] = 25'b00101111_00000011_00110010_0;
      patterns[12038] = 25'b00101111_00000100_00110011_0;
      patterns[12039] = 25'b00101111_00000101_00110100_0;
      patterns[12040] = 25'b00101111_00000110_00110101_0;
      patterns[12041] = 25'b00101111_00000111_00110110_0;
      patterns[12042] = 25'b00101111_00001000_00110111_0;
      patterns[12043] = 25'b00101111_00001001_00111000_0;
      patterns[12044] = 25'b00101111_00001010_00111001_0;
      patterns[12045] = 25'b00101111_00001011_00111010_0;
      patterns[12046] = 25'b00101111_00001100_00111011_0;
      patterns[12047] = 25'b00101111_00001101_00111100_0;
      patterns[12048] = 25'b00101111_00001110_00111101_0;
      patterns[12049] = 25'b00101111_00001111_00111110_0;
      patterns[12050] = 25'b00101111_00010000_00111111_0;
      patterns[12051] = 25'b00101111_00010001_01000000_0;
      patterns[12052] = 25'b00101111_00010010_01000001_0;
      patterns[12053] = 25'b00101111_00010011_01000010_0;
      patterns[12054] = 25'b00101111_00010100_01000011_0;
      patterns[12055] = 25'b00101111_00010101_01000100_0;
      patterns[12056] = 25'b00101111_00010110_01000101_0;
      patterns[12057] = 25'b00101111_00010111_01000110_0;
      patterns[12058] = 25'b00101111_00011000_01000111_0;
      patterns[12059] = 25'b00101111_00011001_01001000_0;
      patterns[12060] = 25'b00101111_00011010_01001001_0;
      patterns[12061] = 25'b00101111_00011011_01001010_0;
      patterns[12062] = 25'b00101111_00011100_01001011_0;
      patterns[12063] = 25'b00101111_00011101_01001100_0;
      patterns[12064] = 25'b00101111_00011110_01001101_0;
      patterns[12065] = 25'b00101111_00011111_01001110_0;
      patterns[12066] = 25'b00101111_00100000_01001111_0;
      patterns[12067] = 25'b00101111_00100001_01010000_0;
      patterns[12068] = 25'b00101111_00100010_01010001_0;
      patterns[12069] = 25'b00101111_00100011_01010010_0;
      patterns[12070] = 25'b00101111_00100100_01010011_0;
      patterns[12071] = 25'b00101111_00100101_01010100_0;
      patterns[12072] = 25'b00101111_00100110_01010101_0;
      patterns[12073] = 25'b00101111_00100111_01010110_0;
      patterns[12074] = 25'b00101111_00101000_01010111_0;
      patterns[12075] = 25'b00101111_00101001_01011000_0;
      patterns[12076] = 25'b00101111_00101010_01011001_0;
      patterns[12077] = 25'b00101111_00101011_01011010_0;
      patterns[12078] = 25'b00101111_00101100_01011011_0;
      patterns[12079] = 25'b00101111_00101101_01011100_0;
      patterns[12080] = 25'b00101111_00101110_01011101_0;
      patterns[12081] = 25'b00101111_00101111_01011110_0;
      patterns[12082] = 25'b00101111_00110000_01011111_0;
      patterns[12083] = 25'b00101111_00110001_01100000_0;
      patterns[12084] = 25'b00101111_00110010_01100001_0;
      patterns[12085] = 25'b00101111_00110011_01100010_0;
      patterns[12086] = 25'b00101111_00110100_01100011_0;
      patterns[12087] = 25'b00101111_00110101_01100100_0;
      patterns[12088] = 25'b00101111_00110110_01100101_0;
      patterns[12089] = 25'b00101111_00110111_01100110_0;
      patterns[12090] = 25'b00101111_00111000_01100111_0;
      patterns[12091] = 25'b00101111_00111001_01101000_0;
      patterns[12092] = 25'b00101111_00111010_01101001_0;
      patterns[12093] = 25'b00101111_00111011_01101010_0;
      patterns[12094] = 25'b00101111_00111100_01101011_0;
      patterns[12095] = 25'b00101111_00111101_01101100_0;
      patterns[12096] = 25'b00101111_00111110_01101101_0;
      patterns[12097] = 25'b00101111_00111111_01101110_0;
      patterns[12098] = 25'b00101111_01000000_01101111_0;
      patterns[12099] = 25'b00101111_01000001_01110000_0;
      patterns[12100] = 25'b00101111_01000010_01110001_0;
      patterns[12101] = 25'b00101111_01000011_01110010_0;
      patterns[12102] = 25'b00101111_01000100_01110011_0;
      patterns[12103] = 25'b00101111_01000101_01110100_0;
      patterns[12104] = 25'b00101111_01000110_01110101_0;
      patterns[12105] = 25'b00101111_01000111_01110110_0;
      patterns[12106] = 25'b00101111_01001000_01110111_0;
      patterns[12107] = 25'b00101111_01001001_01111000_0;
      patterns[12108] = 25'b00101111_01001010_01111001_0;
      patterns[12109] = 25'b00101111_01001011_01111010_0;
      patterns[12110] = 25'b00101111_01001100_01111011_0;
      patterns[12111] = 25'b00101111_01001101_01111100_0;
      patterns[12112] = 25'b00101111_01001110_01111101_0;
      patterns[12113] = 25'b00101111_01001111_01111110_0;
      patterns[12114] = 25'b00101111_01010000_01111111_0;
      patterns[12115] = 25'b00101111_01010001_10000000_0;
      patterns[12116] = 25'b00101111_01010010_10000001_0;
      patterns[12117] = 25'b00101111_01010011_10000010_0;
      patterns[12118] = 25'b00101111_01010100_10000011_0;
      patterns[12119] = 25'b00101111_01010101_10000100_0;
      patterns[12120] = 25'b00101111_01010110_10000101_0;
      patterns[12121] = 25'b00101111_01010111_10000110_0;
      patterns[12122] = 25'b00101111_01011000_10000111_0;
      patterns[12123] = 25'b00101111_01011001_10001000_0;
      patterns[12124] = 25'b00101111_01011010_10001001_0;
      patterns[12125] = 25'b00101111_01011011_10001010_0;
      patterns[12126] = 25'b00101111_01011100_10001011_0;
      patterns[12127] = 25'b00101111_01011101_10001100_0;
      patterns[12128] = 25'b00101111_01011110_10001101_0;
      patterns[12129] = 25'b00101111_01011111_10001110_0;
      patterns[12130] = 25'b00101111_01100000_10001111_0;
      patterns[12131] = 25'b00101111_01100001_10010000_0;
      patterns[12132] = 25'b00101111_01100010_10010001_0;
      patterns[12133] = 25'b00101111_01100011_10010010_0;
      patterns[12134] = 25'b00101111_01100100_10010011_0;
      patterns[12135] = 25'b00101111_01100101_10010100_0;
      patterns[12136] = 25'b00101111_01100110_10010101_0;
      patterns[12137] = 25'b00101111_01100111_10010110_0;
      patterns[12138] = 25'b00101111_01101000_10010111_0;
      patterns[12139] = 25'b00101111_01101001_10011000_0;
      patterns[12140] = 25'b00101111_01101010_10011001_0;
      patterns[12141] = 25'b00101111_01101011_10011010_0;
      patterns[12142] = 25'b00101111_01101100_10011011_0;
      patterns[12143] = 25'b00101111_01101101_10011100_0;
      patterns[12144] = 25'b00101111_01101110_10011101_0;
      patterns[12145] = 25'b00101111_01101111_10011110_0;
      patterns[12146] = 25'b00101111_01110000_10011111_0;
      patterns[12147] = 25'b00101111_01110001_10100000_0;
      patterns[12148] = 25'b00101111_01110010_10100001_0;
      patterns[12149] = 25'b00101111_01110011_10100010_0;
      patterns[12150] = 25'b00101111_01110100_10100011_0;
      patterns[12151] = 25'b00101111_01110101_10100100_0;
      patterns[12152] = 25'b00101111_01110110_10100101_0;
      patterns[12153] = 25'b00101111_01110111_10100110_0;
      patterns[12154] = 25'b00101111_01111000_10100111_0;
      patterns[12155] = 25'b00101111_01111001_10101000_0;
      patterns[12156] = 25'b00101111_01111010_10101001_0;
      patterns[12157] = 25'b00101111_01111011_10101010_0;
      patterns[12158] = 25'b00101111_01111100_10101011_0;
      patterns[12159] = 25'b00101111_01111101_10101100_0;
      patterns[12160] = 25'b00101111_01111110_10101101_0;
      patterns[12161] = 25'b00101111_01111111_10101110_0;
      patterns[12162] = 25'b00101111_10000000_10101111_0;
      patterns[12163] = 25'b00101111_10000001_10110000_0;
      patterns[12164] = 25'b00101111_10000010_10110001_0;
      patterns[12165] = 25'b00101111_10000011_10110010_0;
      patterns[12166] = 25'b00101111_10000100_10110011_0;
      patterns[12167] = 25'b00101111_10000101_10110100_0;
      patterns[12168] = 25'b00101111_10000110_10110101_0;
      patterns[12169] = 25'b00101111_10000111_10110110_0;
      patterns[12170] = 25'b00101111_10001000_10110111_0;
      patterns[12171] = 25'b00101111_10001001_10111000_0;
      patterns[12172] = 25'b00101111_10001010_10111001_0;
      patterns[12173] = 25'b00101111_10001011_10111010_0;
      patterns[12174] = 25'b00101111_10001100_10111011_0;
      patterns[12175] = 25'b00101111_10001101_10111100_0;
      patterns[12176] = 25'b00101111_10001110_10111101_0;
      patterns[12177] = 25'b00101111_10001111_10111110_0;
      patterns[12178] = 25'b00101111_10010000_10111111_0;
      patterns[12179] = 25'b00101111_10010001_11000000_0;
      patterns[12180] = 25'b00101111_10010010_11000001_0;
      patterns[12181] = 25'b00101111_10010011_11000010_0;
      patterns[12182] = 25'b00101111_10010100_11000011_0;
      patterns[12183] = 25'b00101111_10010101_11000100_0;
      patterns[12184] = 25'b00101111_10010110_11000101_0;
      patterns[12185] = 25'b00101111_10010111_11000110_0;
      patterns[12186] = 25'b00101111_10011000_11000111_0;
      patterns[12187] = 25'b00101111_10011001_11001000_0;
      patterns[12188] = 25'b00101111_10011010_11001001_0;
      patterns[12189] = 25'b00101111_10011011_11001010_0;
      patterns[12190] = 25'b00101111_10011100_11001011_0;
      patterns[12191] = 25'b00101111_10011101_11001100_0;
      patterns[12192] = 25'b00101111_10011110_11001101_0;
      patterns[12193] = 25'b00101111_10011111_11001110_0;
      patterns[12194] = 25'b00101111_10100000_11001111_0;
      patterns[12195] = 25'b00101111_10100001_11010000_0;
      patterns[12196] = 25'b00101111_10100010_11010001_0;
      patterns[12197] = 25'b00101111_10100011_11010010_0;
      patterns[12198] = 25'b00101111_10100100_11010011_0;
      patterns[12199] = 25'b00101111_10100101_11010100_0;
      patterns[12200] = 25'b00101111_10100110_11010101_0;
      patterns[12201] = 25'b00101111_10100111_11010110_0;
      patterns[12202] = 25'b00101111_10101000_11010111_0;
      patterns[12203] = 25'b00101111_10101001_11011000_0;
      patterns[12204] = 25'b00101111_10101010_11011001_0;
      patterns[12205] = 25'b00101111_10101011_11011010_0;
      patterns[12206] = 25'b00101111_10101100_11011011_0;
      patterns[12207] = 25'b00101111_10101101_11011100_0;
      patterns[12208] = 25'b00101111_10101110_11011101_0;
      patterns[12209] = 25'b00101111_10101111_11011110_0;
      patterns[12210] = 25'b00101111_10110000_11011111_0;
      patterns[12211] = 25'b00101111_10110001_11100000_0;
      patterns[12212] = 25'b00101111_10110010_11100001_0;
      patterns[12213] = 25'b00101111_10110011_11100010_0;
      patterns[12214] = 25'b00101111_10110100_11100011_0;
      patterns[12215] = 25'b00101111_10110101_11100100_0;
      patterns[12216] = 25'b00101111_10110110_11100101_0;
      patterns[12217] = 25'b00101111_10110111_11100110_0;
      patterns[12218] = 25'b00101111_10111000_11100111_0;
      patterns[12219] = 25'b00101111_10111001_11101000_0;
      patterns[12220] = 25'b00101111_10111010_11101001_0;
      patterns[12221] = 25'b00101111_10111011_11101010_0;
      patterns[12222] = 25'b00101111_10111100_11101011_0;
      patterns[12223] = 25'b00101111_10111101_11101100_0;
      patterns[12224] = 25'b00101111_10111110_11101101_0;
      patterns[12225] = 25'b00101111_10111111_11101110_0;
      patterns[12226] = 25'b00101111_11000000_11101111_0;
      patterns[12227] = 25'b00101111_11000001_11110000_0;
      patterns[12228] = 25'b00101111_11000010_11110001_0;
      patterns[12229] = 25'b00101111_11000011_11110010_0;
      patterns[12230] = 25'b00101111_11000100_11110011_0;
      patterns[12231] = 25'b00101111_11000101_11110100_0;
      patterns[12232] = 25'b00101111_11000110_11110101_0;
      patterns[12233] = 25'b00101111_11000111_11110110_0;
      patterns[12234] = 25'b00101111_11001000_11110111_0;
      patterns[12235] = 25'b00101111_11001001_11111000_0;
      patterns[12236] = 25'b00101111_11001010_11111001_0;
      patterns[12237] = 25'b00101111_11001011_11111010_0;
      patterns[12238] = 25'b00101111_11001100_11111011_0;
      patterns[12239] = 25'b00101111_11001101_11111100_0;
      patterns[12240] = 25'b00101111_11001110_11111101_0;
      patterns[12241] = 25'b00101111_11001111_11111110_0;
      patterns[12242] = 25'b00101111_11010000_11111111_0;
      patterns[12243] = 25'b00101111_11010001_00000000_1;
      patterns[12244] = 25'b00101111_11010010_00000001_1;
      patterns[12245] = 25'b00101111_11010011_00000010_1;
      patterns[12246] = 25'b00101111_11010100_00000011_1;
      patterns[12247] = 25'b00101111_11010101_00000100_1;
      patterns[12248] = 25'b00101111_11010110_00000101_1;
      patterns[12249] = 25'b00101111_11010111_00000110_1;
      patterns[12250] = 25'b00101111_11011000_00000111_1;
      patterns[12251] = 25'b00101111_11011001_00001000_1;
      patterns[12252] = 25'b00101111_11011010_00001001_1;
      patterns[12253] = 25'b00101111_11011011_00001010_1;
      patterns[12254] = 25'b00101111_11011100_00001011_1;
      patterns[12255] = 25'b00101111_11011101_00001100_1;
      patterns[12256] = 25'b00101111_11011110_00001101_1;
      patterns[12257] = 25'b00101111_11011111_00001110_1;
      patterns[12258] = 25'b00101111_11100000_00001111_1;
      patterns[12259] = 25'b00101111_11100001_00010000_1;
      patterns[12260] = 25'b00101111_11100010_00010001_1;
      patterns[12261] = 25'b00101111_11100011_00010010_1;
      patterns[12262] = 25'b00101111_11100100_00010011_1;
      patterns[12263] = 25'b00101111_11100101_00010100_1;
      patterns[12264] = 25'b00101111_11100110_00010101_1;
      patterns[12265] = 25'b00101111_11100111_00010110_1;
      patterns[12266] = 25'b00101111_11101000_00010111_1;
      patterns[12267] = 25'b00101111_11101001_00011000_1;
      patterns[12268] = 25'b00101111_11101010_00011001_1;
      patterns[12269] = 25'b00101111_11101011_00011010_1;
      patterns[12270] = 25'b00101111_11101100_00011011_1;
      patterns[12271] = 25'b00101111_11101101_00011100_1;
      patterns[12272] = 25'b00101111_11101110_00011101_1;
      patterns[12273] = 25'b00101111_11101111_00011110_1;
      patterns[12274] = 25'b00101111_11110000_00011111_1;
      patterns[12275] = 25'b00101111_11110001_00100000_1;
      patterns[12276] = 25'b00101111_11110010_00100001_1;
      patterns[12277] = 25'b00101111_11110011_00100010_1;
      patterns[12278] = 25'b00101111_11110100_00100011_1;
      patterns[12279] = 25'b00101111_11110101_00100100_1;
      patterns[12280] = 25'b00101111_11110110_00100101_1;
      patterns[12281] = 25'b00101111_11110111_00100110_1;
      patterns[12282] = 25'b00101111_11111000_00100111_1;
      patterns[12283] = 25'b00101111_11111001_00101000_1;
      patterns[12284] = 25'b00101111_11111010_00101001_1;
      patterns[12285] = 25'b00101111_11111011_00101010_1;
      patterns[12286] = 25'b00101111_11111100_00101011_1;
      patterns[12287] = 25'b00101111_11111101_00101100_1;
      patterns[12288] = 25'b00101111_11111110_00101101_1;
      patterns[12289] = 25'b00101111_11111111_00101110_1;
      patterns[12290] = 25'b00110000_00000000_00110000_0;
      patterns[12291] = 25'b00110000_00000001_00110001_0;
      patterns[12292] = 25'b00110000_00000010_00110010_0;
      patterns[12293] = 25'b00110000_00000011_00110011_0;
      patterns[12294] = 25'b00110000_00000100_00110100_0;
      patterns[12295] = 25'b00110000_00000101_00110101_0;
      patterns[12296] = 25'b00110000_00000110_00110110_0;
      patterns[12297] = 25'b00110000_00000111_00110111_0;
      patterns[12298] = 25'b00110000_00001000_00111000_0;
      patterns[12299] = 25'b00110000_00001001_00111001_0;
      patterns[12300] = 25'b00110000_00001010_00111010_0;
      patterns[12301] = 25'b00110000_00001011_00111011_0;
      patterns[12302] = 25'b00110000_00001100_00111100_0;
      patterns[12303] = 25'b00110000_00001101_00111101_0;
      patterns[12304] = 25'b00110000_00001110_00111110_0;
      patterns[12305] = 25'b00110000_00001111_00111111_0;
      patterns[12306] = 25'b00110000_00010000_01000000_0;
      patterns[12307] = 25'b00110000_00010001_01000001_0;
      patterns[12308] = 25'b00110000_00010010_01000010_0;
      patterns[12309] = 25'b00110000_00010011_01000011_0;
      patterns[12310] = 25'b00110000_00010100_01000100_0;
      patterns[12311] = 25'b00110000_00010101_01000101_0;
      patterns[12312] = 25'b00110000_00010110_01000110_0;
      patterns[12313] = 25'b00110000_00010111_01000111_0;
      patterns[12314] = 25'b00110000_00011000_01001000_0;
      patterns[12315] = 25'b00110000_00011001_01001001_0;
      patterns[12316] = 25'b00110000_00011010_01001010_0;
      patterns[12317] = 25'b00110000_00011011_01001011_0;
      patterns[12318] = 25'b00110000_00011100_01001100_0;
      patterns[12319] = 25'b00110000_00011101_01001101_0;
      patterns[12320] = 25'b00110000_00011110_01001110_0;
      patterns[12321] = 25'b00110000_00011111_01001111_0;
      patterns[12322] = 25'b00110000_00100000_01010000_0;
      patterns[12323] = 25'b00110000_00100001_01010001_0;
      patterns[12324] = 25'b00110000_00100010_01010010_0;
      patterns[12325] = 25'b00110000_00100011_01010011_0;
      patterns[12326] = 25'b00110000_00100100_01010100_0;
      patterns[12327] = 25'b00110000_00100101_01010101_0;
      patterns[12328] = 25'b00110000_00100110_01010110_0;
      patterns[12329] = 25'b00110000_00100111_01010111_0;
      patterns[12330] = 25'b00110000_00101000_01011000_0;
      patterns[12331] = 25'b00110000_00101001_01011001_0;
      patterns[12332] = 25'b00110000_00101010_01011010_0;
      patterns[12333] = 25'b00110000_00101011_01011011_0;
      patterns[12334] = 25'b00110000_00101100_01011100_0;
      patterns[12335] = 25'b00110000_00101101_01011101_0;
      patterns[12336] = 25'b00110000_00101110_01011110_0;
      patterns[12337] = 25'b00110000_00101111_01011111_0;
      patterns[12338] = 25'b00110000_00110000_01100000_0;
      patterns[12339] = 25'b00110000_00110001_01100001_0;
      patterns[12340] = 25'b00110000_00110010_01100010_0;
      patterns[12341] = 25'b00110000_00110011_01100011_0;
      patterns[12342] = 25'b00110000_00110100_01100100_0;
      patterns[12343] = 25'b00110000_00110101_01100101_0;
      patterns[12344] = 25'b00110000_00110110_01100110_0;
      patterns[12345] = 25'b00110000_00110111_01100111_0;
      patterns[12346] = 25'b00110000_00111000_01101000_0;
      patterns[12347] = 25'b00110000_00111001_01101001_0;
      patterns[12348] = 25'b00110000_00111010_01101010_0;
      patterns[12349] = 25'b00110000_00111011_01101011_0;
      patterns[12350] = 25'b00110000_00111100_01101100_0;
      patterns[12351] = 25'b00110000_00111101_01101101_0;
      patterns[12352] = 25'b00110000_00111110_01101110_0;
      patterns[12353] = 25'b00110000_00111111_01101111_0;
      patterns[12354] = 25'b00110000_01000000_01110000_0;
      patterns[12355] = 25'b00110000_01000001_01110001_0;
      patterns[12356] = 25'b00110000_01000010_01110010_0;
      patterns[12357] = 25'b00110000_01000011_01110011_0;
      patterns[12358] = 25'b00110000_01000100_01110100_0;
      patterns[12359] = 25'b00110000_01000101_01110101_0;
      patterns[12360] = 25'b00110000_01000110_01110110_0;
      patterns[12361] = 25'b00110000_01000111_01110111_0;
      patterns[12362] = 25'b00110000_01001000_01111000_0;
      patterns[12363] = 25'b00110000_01001001_01111001_0;
      patterns[12364] = 25'b00110000_01001010_01111010_0;
      patterns[12365] = 25'b00110000_01001011_01111011_0;
      patterns[12366] = 25'b00110000_01001100_01111100_0;
      patterns[12367] = 25'b00110000_01001101_01111101_0;
      patterns[12368] = 25'b00110000_01001110_01111110_0;
      patterns[12369] = 25'b00110000_01001111_01111111_0;
      patterns[12370] = 25'b00110000_01010000_10000000_0;
      patterns[12371] = 25'b00110000_01010001_10000001_0;
      patterns[12372] = 25'b00110000_01010010_10000010_0;
      patterns[12373] = 25'b00110000_01010011_10000011_0;
      patterns[12374] = 25'b00110000_01010100_10000100_0;
      patterns[12375] = 25'b00110000_01010101_10000101_0;
      patterns[12376] = 25'b00110000_01010110_10000110_0;
      patterns[12377] = 25'b00110000_01010111_10000111_0;
      patterns[12378] = 25'b00110000_01011000_10001000_0;
      patterns[12379] = 25'b00110000_01011001_10001001_0;
      patterns[12380] = 25'b00110000_01011010_10001010_0;
      patterns[12381] = 25'b00110000_01011011_10001011_0;
      patterns[12382] = 25'b00110000_01011100_10001100_0;
      patterns[12383] = 25'b00110000_01011101_10001101_0;
      patterns[12384] = 25'b00110000_01011110_10001110_0;
      patterns[12385] = 25'b00110000_01011111_10001111_0;
      patterns[12386] = 25'b00110000_01100000_10010000_0;
      patterns[12387] = 25'b00110000_01100001_10010001_0;
      patterns[12388] = 25'b00110000_01100010_10010010_0;
      patterns[12389] = 25'b00110000_01100011_10010011_0;
      patterns[12390] = 25'b00110000_01100100_10010100_0;
      patterns[12391] = 25'b00110000_01100101_10010101_0;
      patterns[12392] = 25'b00110000_01100110_10010110_0;
      patterns[12393] = 25'b00110000_01100111_10010111_0;
      patterns[12394] = 25'b00110000_01101000_10011000_0;
      patterns[12395] = 25'b00110000_01101001_10011001_0;
      patterns[12396] = 25'b00110000_01101010_10011010_0;
      patterns[12397] = 25'b00110000_01101011_10011011_0;
      patterns[12398] = 25'b00110000_01101100_10011100_0;
      patterns[12399] = 25'b00110000_01101101_10011101_0;
      patterns[12400] = 25'b00110000_01101110_10011110_0;
      patterns[12401] = 25'b00110000_01101111_10011111_0;
      patterns[12402] = 25'b00110000_01110000_10100000_0;
      patterns[12403] = 25'b00110000_01110001_10100001_0;
      patterns[12404] = 25'b00110000_01110010_10100010_0;
      patterns[12405] = 25'b00110000_01110011_10100011_0;
      patterns[12406] = 25'b00110000_01110100_10100100_0;
      patterns[12407] = 25'b00110000_01110101_10100101_0;
      patterns[12408] = 25'b00110000_01110110_10100110_0;
      patterns[12409] = 25'b00110000_01110111_10100111_0;
      patterns[12410] = 25'b00110000_01111000_10101000_0;
      patterns[12411] = 25'b00110000_01111001_10101001_0;
      patterns[12412] = 25'b00110000_01111010_10101010_0;
      patterns[12413] = 25'b00110000_01111011_10101011_0;
      patterns[12414] = 25'b00110000_01111100_10101100_0;
      patterns[12415] = 25'b00110000_01111101_10101101_0;
      patterns[12416] = 25'b00110000_01111110_10101110_0;
      patterns[12417] = 25'b00110000_01111111_10101111_0;
      patterns[12418] = 25'b00110000_10000000_10110000_0;
      patterns[12419] = 25'b00110000_10000001_10110001_0;
      patterns[12420] = 25'b00110000_10000010_10110010_0;
      patterns[12421] = 25'b00110000_10000011_10110011_0;
      patterns[12422] = 25'b00110000_10000100_10110100_0;
      patterns[12423] = 25'b00110000_10000101_10110101_0;
      patterns[12424] = 25'b00110000_10000110_10110110_0;
      patterns[12425] = 25'b00110000_10000111_10110111_0;
      patterns[12426] = 25'b00110000_10001000_10111000_0;
      patterns[12427] = 25'b00110000_10001001_10111001_0;
      patterns[12428] = 25'b00110000_10001010_10111010_0;
      patterns[12429] = 25'b00110000_10001011_10111011_0;
      patterns[12430] = 25'b00110000_10001100_10111100_0;
      patterns[12431] = 25'b00110000_10001101_10111101_0;
      patterns[12432] = 25'b00110000_10001110_10111110_0;
      patterns[12433] = 25'b00110000_10001111_10111111_0;
      patterns[12434] = 25'b00110000_10010000_11000000_0;
      patterns[12435] = 25'b00110000_10010001_11000001_0;
      patterns[12436] = 25'b00110000_10010010_11000010_0;
      patterns[12437] = 25'b00110000_10010011_11000011_0;
      patterns[12438] = 25'b00110000_10010100_11000100_0;
      patterns[12439] = 25'b00110000_10010101_11000101_0;
      patterns[12440] = 25'b00110000_10010110_11000110_0;
      patterns[12441] = 25'b00110000_10010111_11000111_0;
      patterns[12442] = 25'b00110000_10011000_11001000_0;
      patterns[12443] = 25'b00110000_10011001_11001001_0;
      patterns[12444] = 25'b00110000_10011010_11001010_0;
      patterns[12445] = 25'b00110000_10011011_11001011_0;
      patterns[12446] = 25'b00110000_10011100_11001100_0;
      patterns[12447] = 25'b00110000_10011101_11001101_0;
      patterns[12448] = 25'b00110000_10011110_11001110_0;
      patterns[12449] = 25'b00110000_10011111_11001111_0;
      patterns[12450] = 25'b00110000_10100000_11010000_0;
      patterns[12451] = 25'b00110000_10100001_11010001_0;
      patterns[12452] = 25'b00110000_10100010_11010010_0;
      patterns[12453] = 25'b00110000_10100011_11010011_0;
      patterns[12454] = 25'b00110000_10100100_11010100_0;
      patterns[12455] = 25'b00110000_10100101_11010101_0;
      patterns[12456] = 25'b00110000_10100110_11010110_0;
      patterns[12457] = 25'b00110000_10100111_11010111_0;
      patterns[12458] = 25'b00110000_10101000_11011000_0;
      patterns[12459] = 25'b00110000_10101001_11011001_0;
      patterns[12460] = 25'b00110000_10101010_11011010_0;
      patterns[12461] = 25'b00110000_10101011_11011011_0;
      patterns[12462] = 25'b00110000_10101100_11011100_0;
      patterns[12463] = 25'b00110000_10101101_11011101_0;
      patterns[12464] = 25'b00110000_10101110_11011110_0;
      patterns[12465] = 25'b00110000_10101111_11011111_0;
      patterns[12466] = 25'b00110000_10110000_11100000_0;
      patterns[12467] = 25'b00110000_10110001_11100001_0;
      patterns[12468] = 25'b00110000_10110010_11100010_0;
      patterns[12469] = 25'b00110000_10110011_11100011_0;
      patterns[12470] = 25'b00110000_10110100_11100100_0;
      patterns[12471] = 25'b00110000_10110101_11100101_0;
      patterns[12472] = 25'b00110000_10110110_11100110_0;
      patterns[12473] = 25'b00110000_10110111_11100111_0;
      patterns[12474] = 25'b00110000_10111000_11101000_0;
      patterns[12475] = 25'b00110000_10111001_11101001_0;
      patterns[12476] = 25'b00110000_10111010_11101010_0;
      patterns[12477] = 25'b00110000_10111011_11101011_0;
      patterns[12478] = 25'b00110000_10111100_11101100_0;
      patterns[12479] = 25'b00110000_10111101_11101101_0;
      patterns[12480] = 25'b00110000_10111110_11101110_0;
      patterns[12481] = 25'b00110000_10111111_11101111_0;
      patterns[12482] = 25'b00110000_11000000_11110000_0;
      patterns[12483] = 25'b00110000_11000001_11110001_0;
      patterns[12484] = 25'b00110000_11000010_11110010_0;
      patterns[12485] = 25'b00110000_11000011_11110011_0;
      patterns[12486] = 25'b00110000_11000100_11110100_0;
      patterns[12487] = 25'b00110000_11000101_11110101_0;
      patterns[12488] = 25'b00110000_11000110_11110110_0;
      patterns[12489] = 25'b00110000_11000111_11110111_0;
      patterns[12490] = 25'b00110000_11001000_11111000_0;
      patterns[12491] = 25'b00110000_11001001_11111001_0;
      patterns[12492] = 25'b00110000_11001010_11111010_0;
      patterns[12493] = 25'b00110000_11001011_11111011_0;
      patterns[12494] = 25'b00110000_11001100_11111100_0;
      patterns[12495] = 25'b00110000_11001101_11111101_0;
      patterns[12496] = 25'b00110000_11001110_11111110_0;
      patterns[12497] = 25'b00110000_11001111_11111111_0;
      patterns[12498] = 25'b00110000_11010000_00000000_1;
      patterns[12499] = 25'b00110000_11010001_00000001_1;
      patterns[12500] = 25'b00110000_11010010_00000010_1;
      patterns[12501] = 25'b00110000_11010011_00000011_1;
      patterns[12502] = 25'b00110000_11010100_00000100_1;
      patterns[12503] = 25'b00110000_11010101_00000101_1;
      patterns[12504] = 25'b00110000_11010110_00000110_1;
      patterns[12505] = 25'b00110000_11010111_00000111_1;
      patterns[12506] = 25'b00110000_11011000_00001000_1;
      patterns[12507] = 25'b00110000_11011001_00001001_1;
      patterns[12508] = 25'b00110000_11011010_00001010_1;
      patterns[12509] = 25'b00110000_11011011_00001011_1;
      patterns[12510] = 25'b00110000_11011100_00001100_1;
      patterns[12511] = 25'b00110000_11011101_00001101_1;
      patterns[12512] = 25'b00110000_11011110_00001110_1;
      patterns[12513] = 25'b00110000_11011111_00001111_1;
      patterns[12514] = 25'b00110000_11100000_00010000_1;
      patterns[12515] = 25'b00110000_11100001_00010001_1;
      patterns[12516] = 25'b00110000_11100010_00010010_1;
      patterns[12517] = 25'b00110000_11100011_00010011_1;
      patterns[12518] = 25'b00110000_11100100_00010100_1;
      patterns[12519] = 25'b00110000_11100101_00010101_1;
      patterns[12520] = 25'b00110000_11100110_00010110_1;
      patterns[12521] = 25'b00110000_11100111_00010111_1;
      patterns[12522] = 25'b00110000_11101000_00011000_1;
      patterns[12523] = 25'b00110000_11101001_00011001_1;
      patterns[12524] = 25'b00110000_11101010_00011010_1;
      patterns[12525] = 25'b00110000_11101011_00011011_1;
      patterns[12526] = 25'b00110000_11101100_00011100_1;
      patterns[12527] = 25'b00110000_11101101_00011101_1;
      patterns[12528] = 25'b00110000_11101110_00011110_1;
      patterns[12529] = 25'b00110000_11101111_00011111_1;
      patterns[12530] = 25'b00110000_11110000_00100000_1;
      patterns[12531] = 25'b00110000_11110001_00100001_1;
      patterns[12532] = 25'b00110000_11110010_00100010_1;
      patterns[12533] = 25'b00110000_11110011_00100011_1;
      patterns[12534] = 25'b00110000_11110100_00100100_1;
      patterns[12535] = 25'b00110000_11110101_00100101_1;
      patterns[12536] = 25'b00110000_11110110_00100110_1;
      patterns[12537] = 25'b00110000_11110111_00100111_1;
      patterns[12538] = 25'b00110000_11111000_00101000_1;
      patterns[12539] = 25'b00110000_11111001_00101001_1;
      patterns[12540] = 25'b00110000_11111010_00101010_1;
      patterns[12541] = 25'b00110000_11111011_00101011_1;
      patterns[12542] = 25'b00110000_11111100_00101100_1;
      patterns[12543] = 25'b00110000_11111101_00101101_1;
      patterns[12544] = 25'b00110000_11111110_00101110_1;
      patterns[12545] = 25'b00110000_11111111_00101111_1;
      patterns[12546] = 25'b00110001_00000000_00110001_0;
      patterns[12547] = 25'b00110001_00000001_00110010_0;
      patterns[12548] = 25'b00110001_00000010_00110011_0;
      patterns[12549] = 25'b00110001_00000011_00110100_0;
      patterns[12550] = 25'b00110001_00000100_00110101_0;
      patterns[12551] = 25'b00110001_00000101_00110110_0;
      patterns[12552] = 25'b00110001_00000110_00110111_0;
      patterns[12553] = 25'b00110001_00000111_00111000_0;
      patterns[12554] = 25'b00110001_00001000_00111001_0;
      patterns[12555] = 25'b00110001_00001001_00111010_0;
      patterns[12556] = 25'b00110001_00001010_00111011_0;
      patterns[12557] = 25'b00110001_00001011_00111100_0;
      patterns[12558] = 25'b00110001_00001100_00111101_0;
      patterns[12559] = 25'b00110001_00001101_00111110_0;
      patterns[12560] = 25'b00110001_00001110_00111111_0;
      patterns[12561] = 25'b00110001_00001111_01000000_0;
      patterns[12562] = 25'b00110001_00010000_01000001_0;
      patterns[12563] = 25'b00110001_00010001_01000010_0;
      patterns[12564] = 25'b00110001_00010010_01000011_0;
      patterns[12565] = 25'b00110001_00010011_01000100_0;
      patterns[12566] = 25'b00110001_00010100_01000101_0;
      patterns[12567] = 25'b00110001_00010101_01000110_0;
      patterns[12568] = 25'b00110001_00010110_01000111_0;
      patterns[12569] = 25'b00110001_00010111_01001000_0;
      patterns[12570] = 25'b00110001_00011000_01001001_0;
      patterns[12571] = 25'b00110001_00011001_01001010_0;
      patterns[12572] = 25'b00110001_00011010_01001011_0;
      patterns[12573] = 25'b00110001_00011011_01001100_0;
      patterns[12574] = 25'b00110001_00011100_01001101_0;
      patterns[12575] = 25'b00110001_00011101_01001110_0;
      patterns[12576] = 25'b00110001_00011110_01001111_0;
      patterns[12577] = 25'b00110001_00011111_01010000_0;
      patterns[12578] = 25'b00110001_00100000_01010001_0;
      patterns[12579] = 25'b00110001_00100001_01010010_0;
      patterns[12580] = 25'b00110001_00100010_01010011_0;
      patterns[12581] = 25'b00110001_00100011_01010100_0;
      patterns[12582] = 25'b00110001_00100100_01010101_0;
      patterns[12583] = 25'b00110001_00100101_01010110_0;
      patterns[12584] = 25'b00110001_00100110_01010111_0;
      patterns[12585] = 25'b00110001_00100111_01011000_0;
      patterns[12586] = 25'b00110001_00101000_01011001_0;
      patterns[12587] = 25'b00110001_00101001_01011010_0;
      patterns[12588] = 25'b00110001_00101010_01011011_0;
      patterns[12589] = 25'b00110001_00101011_01011100_0;
      patterns[12590] = 25'b00110001_00101100_01011101_0;
      patterns[12591] = 25'b00110001_00101101_01011110_0;
      patterns[12592] = 25'b00110001_00101110_01011111_0;
      patterns[12593] = 25'b00110001_00101111_01100000_0;
      patterns[12594] = 25'b00110001_00110000_01100001_0;
      patterns[12595] = 25'b00110001_00110001_01100010_0;
      patterns[12596] = 25'b00110001_00110010_01100011_0;
      patterns[12597] = 25'b00110001_00110011_01100100_0;
      patterns[12598] = 25'b00110001_00110100_01100101_0;
      patterns[12599] = 25'b00110001_00110101_01100110_0;
      patterns[12600] = 25'b00110001_00110110_01100111_0;
      patterns[12601] = 25'b00110001_00110111_01101000_0;
      patterns[12602] = 25'b00110001_00111000_01101001_0;
      patterns[12603] = 25'b00110001_00111001_01101010_0;
      patterns[12604] = 25'b00110001_00111010_01101011_0;
      patterns[12605] = 25'b00110001_00111011_01101100_0;
      patterns[12606] = 25'b00110001_00111100_01101101_0;
      patterns[12607] = 25'b00110001_00111101_01101110_0;
      patterns[12608] = 25'b00110001_00111110_01101111_0;
      patterns[12609] = 25'b00110001_00111111_01110000_0;
      patterns[12610] = 25'b00110001_01000000_01110001_0;
      patterns[12611] = 25'b00110001_01000001_01110010_0;
      patterns[12612] = 25'b00110001_01000010_01110011_0;
      patterns[12613] = 25'b00110001_01000011_01110100_0;
      patterns[12614] = 25'b00110001_01000100_01110101_0;
      patterns[12615] = 25'b00110001_01000101_01110110_0;
      patterns[12616] = 25'b00110001_01000110_01110111_0;
      patterns[12617] = 25'b00110001_01000111_01111000_0;
      patterns[12618] = 25'b00110001_01001000_01111001_0;
      patterns[12619] = 25'b00110001_01001001_01111010_0;
      patterns[12620] = 25'b00110001_01001010_01111011_0;
      patterns[12621] = 25'b00110001_01001011_01111100_0;
      patterns[12622] = 25'b00110001_01001100_01111101_0;
      patterns[12623] = 25'b00110001_01001101_01111110_0;
      patterns[12624] = 25'b00110001_01001110_01111111_0;
      patterns[12625] = 25'b00110001_01001111_10000000_0;
      patterns[12626] = 25'b00110001_01010000_10000001_0;
      patterns[12627] = 25'b00110001_01010001_10000010_0;
      patterns[12628] = 25'b00110001_01010010_10000011_0;
      patterns[12629] = 25'b00110001_01010011_10000100_0;
      patterns[12630] = 25'b00110001_01010100_10000101_0;
      patterns[12631] = 25'b00110001_01010101_10000110_0;
      patterns[12632] = 25'b00110001_01010110_10000111_0;
      patterns[12633] = 25'b00110001_01010111_10001000_0;
      patterns[12634] = 25'b00110001_01011000_10001001_0;
      patterns[12635] = 25'b00110001_01011001_10001010_0;
      patterns[12636] = 25'b00110001_01011010_10001011_0;
      patterns[12637] = 25'b00110001_01011011_10001100_0;
      patterns[12638] = 25'b00110001_01011100_10001101_0;
      patterns[12639] = 25'b00110001_01011101_10001110_0;
      patterns[12640] = 25'b00110001_01011110_10001111_0;
      patterns[12641] = 25'b00110001_01011111_10010000_0;
      patterns[12642] = 25'b00110001_01100000_10010001_0;
      patterns[12643] = 25'b00110001_01100001_10010010_0;
      patterns[12644] = 25'b00110001_01100010_10010011_0;
      patterns[12645] = 25'b00110001_01100011_10010100_0;
      patterns[12646] = 25'b00110001_01100100_10010101_0;
      patterns[12647] = 25'b00110001_01100101_10010110_0;
      patterns[12648] = 25'b00110001_01100110_10010111_0;
      patterns[12649] = 25'b00110001_01100111_10011000_0;
      patterns[12650] = 25'b00110001_01101000_10011001_0;
      patterns[12651] = 25'b00110001_01101001_10011010_0;
      patterns[12652] = 25'b00110001_01101010_10011011_0;
      patterns[12653] = 25'b00110001_01101011_10011100_0;
      patterns[12654] = 25'b00110001_01101100_10011101_0;
      patterns[12655] = 25'b00110001_01101101_10011110_0;
      patterns[12656] = 25'b00110001_01101110_10011111_0;
      patterns[12657] = 25'b00110001_01101111_10100000_0;
      patterns[12658] = 25'b00110001_01110000_10100001_0;
      patterns[12659] = 25'b00110001_01110001_10100010_0;
      patterns[12660] = 25'b00110001_01110010_10100011_0;
      patterns[12661] = 25'b00110001_01110011_10100100_0;
      patterns[12662] = 25'b00110001_01110100_10100101_0;
      patterns[12663] = 25'b00110001_01110101_10100110_0;
      patterns[12664] = 25'b00110001_01110110_10100111_0;
      patterns[12665] = 25'b00110001_01110111_10101000_0;
      patterns[12666] = 25'b00110001_01111000_10101001_0;
      patterns[12667] = 25'b00110001_01111001_10101010_0;
      patterns[12668] = 25'b00110001_01111010_10101011_0;
      patterns[12669] = 25'b00110001_01111011_10101100_0;
      patterns[12670] = 25'b00110001_01111100_10101101_0;
      patterns[12671] = 25'b00110001_01111101_10101110_0;
      patterns[12672] = 25'b00110001_01111110_10101111_0;
      patterns[12673] = 25'b00110001_01111111_10110000_0;
      patterns[12674] = 25'b00110001_10000000_10110001_0;
      patterns[12675] = 25'b00110001_10000001_10110010_0;
      patterns[12676] = 25'b00110001_10000010_10110011_0;
      patterns[12677] = 25'b00110001_10000011_10110100_0;
      patterns[12678] = 25'b00110001_10000100_10110101_0;
      patterns[12679] = 25'b00110001_10000101_10110110_0;
      patterns[12680] = 25'b00110001_10000110_10110111_0;
      patterns[12681] = 25'b00110001_10000111_10111000_0;
      patterns[12682] = 25'b00110001_10001000_10111001_0;
      patterns[12683] = 25'b00110001_10001001_10111010_0;
      patterns[12684] = 25'b00110001_10001010_10111011_0;
      patterns[12685] = 25'b00110001_10001011_10111100_0;
      patterns[12686] = 25'b00110001_10001100_10111101_0;
      patterns[12687] = 25'b00110001_10001101_10111110_0;
      patterns[12688] = 25'b00110001_10001110_10111111_0;
      patterns[12689] = 25'b00110001_10001111_11000000_0;
      patterns[12690] = 25'b00110001_10010000_11000001_0;
      patterns[12691] = 25'b00110001_10010001_11000010_0;
      patterns[12692] = 25'b00110001_10010010_11000011_0;
      patterns[12693] = 25'b00110001_10010011_11000100_0;
      patterns[12694] = 25'b00110001_10010100_11000101_0;
      patterns[12695] = 25'b00110001_10010101_11000110_0;
      patterns[12696] = 25'b00110001_10010110_11000111_0;
      patterns[12697] = 25'b00110001_10010111_11001000_0;
      patterns[12698] = 25'b00110001_10011000_11001001_0;
      patterns[12699] = 25'b00110001_10011001_11001010_0;
      patterns[12700] = 25'b00110001_10011010_11001011_0;
      patterns[12701] = 25'b00110001_10011011_11001100_0;
      patterns[12702] = 25'b00110001_10011100_11001101_0;
      patterns[12703] = 25'b00110001_10011101_11001110_0;
      patterns[12704] = 25'b00110001_10011110_11001111_0;
      patterns[12705] = 25'b00110001_10011111_11010000_0;
      patterns[12706] = 25'b00110001_10100000_11010001_0;
      patterns[12707] = 25'b00110001_10100001_11010010_0;
      patterns[12708] = 25'b00110001_10100010_11010011_0;
      patterns[12709] = 25'b00110001_10100011_11010100_0;
      patterns[12710] = 25'b00110001_10100100_11010101_0;
      patterns[12711] = 25'b00110001_10100101_11010110_0;
      patterns[12712] = 25'b00110001_10100110_11010111_0;
      patterns[12713] = 25'b00110001_10100111_11011000_0;
      patterns[12714] = 25'b00110001_10101000_11011001_0;
      patterns[12715] = 25'b00110001_10101001_11011010_0;
      patterns[12716] = 25'b00110001_10101010_11011011_0;
      patterns[12717] = 25'b00110001_10101011_11011100_0;
      patterns[12718] = 25'b00110001_10101100_11011101_0;
      patterns[12719] = 25'b00110001_10101101_11011110_0;
      patterns[12720] = 25'b00110001_10101110_11011111_0;
      patterns[12721] = 25'b00110001_10101111_11100000_0;
      patterns[12722] = 25'b00110001_10110000_11100001_0;
      patterns[12723] = 25'b00110001_10110001_11100010_0;
      patterns[12724] = 25'b00110001_10110010_11100011_0;
      patterns[12725] = 25'b00110001_10110011_11100100_0;
      patterns[12726] = 25'b00110001_10110100_11100101_0;
      patterns[12727] = 25'b00110001_10110101_11100110_0;
      patterns[12728] = 25'b00110001_10110110_11100111_0;
      patterns[12729] = 25'b00110001_10110111_11101000_0;
      patterns[12730] = 25'b00110001_10111000_11101001_0;
      patterns[12731] = 25'b00110001_10111001_11101010_0;
      patterns[12732] = 25'b00110001_10111010_11101011_0;
      patterns[12733] = 25'b00110001_10111011_11101100_0;
      patterns[12734] = 25'b00110001_10111100_11101101_0;
      patterns[12735] = 25'b00110001_10111101_11101110_0;
      patterns[12736] = 25'b00110001_10111110_11101111_0;
      patterns[12737] = 25'b00110001_10111111_11110000_0;
      patterns[12738] = 25'b00110001_11000000_11110001_0;
      patterns[12739] = 25'b00110001_11000001_11110010_0;
      patterns[12740] = 25'b00110001_11000010_11110011_0;
      patterns[12741] = 25'b00110001_11000011_11110100_0;
      patterns[12742] = 25'b00110001_11000100_11110101_0;
      patterns[12743] = 25'b00110001_11000101_11110110_0;
      patterns[12744] = 25'b00110001_11000110_11110111_0;
      patterns[12745] = 25'b00110001_11000111_11111000_0;
      patterns[12746] = 25'b00110001_11001000_11111001_0;
      patterns[12747] = 25'b00110001_11001001_11111010_0;
      patterns[12748] = 25'b00110001_11001010_11111011_0;
      patterns[12749] = 25'b00110001_11001011_11111100_0;
      patterns[12750] = 25'b00110001_11001100_11111101_0;
      patterns[12751] = 25'b00110001_11001101_11111110_0;
      patterns[12752] = 25'b00110001_11001110_11111111_0;
      patterns[12753] = 25'b00110001_11001111_00000000_1;
      patterns[12754] = 25'b00110001_11010000_00000001_1;
      patterns[12755] = 25'b00110001_11010001_00000010_1;
      patterns[12756] = 25'b00110001_11010010_00000011_1;
      patterns[12757] = 25'b00110001_11010011_00000100_1;
      patterns[12758] = 25'b00110001_11010100_00000101_1;
      patterns[12759] = 25'b00110001_11010101_00000110_1;
      patterns[12760] = 25'b00110001_11010110_00000111_1;
      patterns[12761] = 25'b00110001_11010111_00001000_1;
      patterns[12762] = 25'b00110001_11011000_00001001_1;
      patterns[12763] = 25'b00110001_11011001_00001010_1;
      patterns[12764] = 25'b00110001_11011010_00001011_1;
      patterns[12765] = 25'b00110001_11011011_00001100_1;
      patterns[12766] = 25'b00110001_11011100_00001101_1;
      patterns[12767] = 25'b00110001_11011101_00001110_1;
      patterns[12768] = 25'b00110001_11011110_00001111_1;
      patterns[12769] = 25'b00110001_11011111_00010000_1;
      patterns[12770] = 25'b00110001_11100000_00010001_1;
      patterns[12771] = 25'b00110001_11100001_00010010_1;
      patterns[12772] = 25'b00110001_11100010_00010011_1;
      patterns[12773] = 25'b00110001_11100011_00010100_1;
      patterns[12774] = 25'b00110001_11100100_00010101_1;
      patterns[12775] = 25'b00110001_11100101_00010110_1;
      patterns[12776] = 25'b00110001_11100110_00010111_1;
      patterns[12777] = 25'b00110001_11100111_00011000_1;
      patterns[12778] = 25'b00110001_11101000_00011001_1;
      patterns[12779] = 25'b00110001_11101001_00011010_1;
      patterns[12780] = 25'b00110001_11101010_00011011_1;
      patterns[12781] = 25'b00110001_11101011_00011100_1;
      patterns[12782] = 25'b00110001_11101100_00011101_1;
      patterns[12783] = 25'b00110001_11101101_00011110_1;
      patterns[12784] = 25'b00110001_11101110_00011111_1;
      patterns[12785] = 25'b00110001_11101111_00100000_1;
      patterns[12786] = 25'b00110001_11110000_00100001_1;
      patterns[12787] = 25'b00110001_11110001_00100010_1;
      patterns[12788] = 25'b00110001_11110010_00100011_1;
      patterns[12789] = 25'b00110001_11110011_00100100_1;
      patterns[12790] = 25'b00110001_11110100_00100101_1;
      patterns[12791] = 25'b00110001_11110101_00100110_1;
      patterns[12792] = 25'b00110001_11110110_00100111_1;
      patterns[12793] = 25'b00110001_11110111_00101000_1;
      patterns[12794] = 25'b00110001_11111000_00101001_1;
      patterns[12795] = 25'b00110001_11111001_00101010_1;
      patterns[12796] = 25'b00110001_11111010_00101011_1;
      patterns[12797] = 25'b00110001_11111011_00101100_1;
      patterns[12798] = 25'b00110001_11111100_00101101_1;
      patterns[12799] = 25'b00110001_11111101_00101110_1;
      patterns[12800] = 25'b00110001_11111110_00101111_1;
      patterns[12801] = 25'b00110001_11111111_00110000_1;
      patterns[12802] = 25'b00110010_00000000_00110010_0;
      patterns[12803] = 25'b00110010_00000001_00110011_0;
      patterns[12804] = 25'b00110010_00000010_00110100_0;
      patterns[12805] = 25'b00110010_00000011_00110101_0;
      patterns[12806] = 25'b00110010_00000100_00110110_0;
      patterns[12807] = 25'b00110010_00000101_00110111_0;
      patterns[12808] = 25'b00110010_00000110_00111000_0;
      patterns[12809] = 25'b00110010_00000111_00111001_0;
      patterns[12810] = 25'b00110010_00001000_00111010_0;
      patterns[12811] = 25'b00110010_00001001_00111011_0;
      patterns[12812] = 25'b00110010_00001010_00111100_0;
      patterns[12813] = 25'b00110010_00001011_00111101_0;
      patterns[12814] = 25'b00110010_00001100_00111110_0;
      patterns[12815] = 25'b00110010_00001101_00111111_0;
      patterns[12816] = 25'b00110010_00001110_01000000_0;
      patterns[12817] = 25'b00110010_00001111_01000001_0;
      patterns[12818] = 25'b00110010_00010000_01000010_0;
      patterns[12819] = 25'b00110010_00010001_01000011_0;
      patterns[12820] = 25'b00110010_00010010_01000100_0;
      patterns[12821] = 25'b00110010_00010011_01000101_0;
      patterns[12822] = 25'b00110010_00010100_01000110_0;
      patterns[12823] = 25'b00110010_00010101_01000111_0;
      patterns[12824] = 25'b00110010_00010110_01001000_0;
      patterns[12825] = 25'b00110010_00010111_01001001_0;
      patterns[12826] = 25'b00110010_00011000_01001010_0;
      patterns[12827] = 25'b00110010_00011001_01001011_0;
      patterns[12828] = 25'b00110010_00011010_01001100_0;
      patterns[12829] = 25'b00110010_00011011_01001101_0;
      patterns[12830] = 25'b00110010_00011100_01001110_0;
      patterns[12831] = 25'b00110010_00011101_01001111_0;
      patterns[12832] = 25'b00110010_00011110_01010000_0;
      patterns[12833] = 25'b00110010_00011111_01010001_0;
      patterns[12834] = 25'b00110010_00100000_01010010_0;
      patterns[12835] = 25'b00110010_00100001_01010011_0;
      patterns[12836] = 25'b00110010_00100010_01010100_0;
      patterns[12837] = 25'b00110010_00100011_01010101_0;
      patterns[12838] = 25'b00110010_00100100_01010110_0;
      patterns[12839] = 25'b00110010_00100101_01010111_0;
      patterns[12840] = 25'b00110010_00100110_01011000_0;
      patterns[12841] = 25'b00110010_00100111_01011001_0;
      patterns[12842] = 25'b00110010_00101000_01011010_0;
      patterns[12843] = 25'b00110010_00101001_01011011_0;
      patterns[12844] = 25'b00110010_00101010_01011100_0;
      patterns[12845] = 25'b00110010_00101011_01011101_0;
      patterns[12846] = 25'b00110010_00101100_01011110_0;
      patterns[12847] = 25'b00110010_00101101_01011111_0;
      patterns[12848] = 25'b00110010_00101110_01100000_0;
      patterns[12849] = 25'b00110010_00101111_01100001_0;
      patterns[12850] = 25'b00110010_00110000_01100010_0;
      patterns[12851] = 25'b00110010_00110001_01100011_0;
      patterns[12852] = 25'b00110010_00110010_01100100_0;
      patterns[12853] = 25'b00110010_00110011_01100101_0;
      patterns[12854] = 25'b00110010_00110100_01100110_0;
      patterns[12855] = 25'b00110010_00110101_01100111_0;
      patterns[12856] = 25'b00110010_00110110_01101000_0;
      patterns[12857] = 25'b00110010_00110111_01101001_0;
      patterns[12858] = 25'b00110010_00111000_01101010_0;
      patterns[12859] = 25'b00110010_00111001_01101011_0;
      patterns[12860] = 25'b00110010_00111010_01101100_0;
      patterns[12861] = 25'b00110010_00111011_01101101_0;
      patterns[12862] = 25'b00110010_00111100_01101110_0;
      patterns[12863] = 25'b00110010_00111101_01101111_0;
      patterns[12864] = 25'b00110010_00111110_01110000_0;
      patterns[12865] = 25'b00110010_00111111_01110001_0;
      patterns[12866] = 25'b00110010_01000000_01110010_0;
      patterns[12867] = 25'b00110010_01000001_01110011_0;
      patterns[12868] = 25'b00110010_01000010_01110100_0;
      patterns[12869] = 25'b00110010_01000011_01110101_0;
      patterns[12870] = 25'b00110010_01000100_01110110_0;
      patterns[12871] = 25'b00110010_01000101_01110111_0;
      patterns[12872] = 25'b00110010_01000110_01111000_0;
      patterns[12873] = 25'b00110010_01000111_01111001_0;
      patterns[12874] = 25'b00110010_01001000_01111010_0;
      patterns[12875] = 25'b00110010_01001001_01111011_0;
      patterns[12876] = 25'b00110010_01001010_01111100_0;
      patterns[12877] = 25'b00110010_01001011_01111101_0;
      patterns[12878] = 25'b00110010_01001100_01111110_0;
      patterns[12879] = 25'b00110010_01001101_01111111_0;
      patterns[12880] = 25'b00110010_01001110_10000000_0;
      patterns[12881] = 25'b00110010_01001111_10000001_0;
      patterns[12882] = 25'b00110010_01010000_10000010_0;
      patterns[12883] = 25'b00110010_01010001_10000011_0;
      patterns[12884] = 25'b00110010_01010010_10000100_0;
      patterns[12885] = 25'b00110010_01010011_10000101_0;
      patterns[12886] = 25'b00110010_01010100_10000110_0;
      patterns[12887] = 25'b00110010_01010101_10000111_0;
      patterns[12888] = 25'b00110010_01010110_10001000_0;
      patterns[12889] = 25'b00110010_01010111_10001001_0;
      patterns[12890] = 25'b00110010_01011000_10001010_0;
      patterns[12891] = 25'b00110010_01011001_10001011_0;
      patterns[12892] = 25'b00110010_01011010_10001100_0;
      patterns[12893] = 25'b00110010_01011011_10001101_0;
      patterns[12894] = 25'b00110010_01011100_10001110_0;
      patterns[12895] = 25'b00110010_01011101_10001111_0;
      patterns[12896] = 25'b00110010_01011110_10010000_0;
      patterns[12897] = 25'b00110010_01011111_10010001_0;
      patterns[12898] = 25'b00110010_01100000_10010010_0;
      patterns[12899] = 25'b00110010_01100001_10010011_0;
      patterns[12900] = 25'b00110010_01100010_10010100_0;
      patterns[12901] = 25'b00110010_01100011_10010101_0;
      patterns[12902] = 25'b00110010_01100100_10010110_0;
      patterns[12903] = 25'b00110010_01100101_10010111_0;
      patterns[12904] = 25'b00110010_01100110_10011000_0;
      patterns[12905] = 25'b00110010_01100111_10011001_0;
      patterns[12906] = 25'b00110010_01101000_10011010_0;
      patterns[12907] = 25'b00110010_01101001_10011011_0;
      patterns[12908] = 25'b00110010_01101010_10011100_0;
      patterns[12909] = 25'b00110010_01101011_10011101_0;
      patterns[12910] = 25'b00110010_01101100_10011110_0;
      patterns[12911] = 25'b00110010_01101101_10011111_0;
      patterns[12912] = 25'b00110010_01101110_10100000_0;
      patterns[12913] = 25'b00110010_01101111_10100001_0;
      patterns[12914] = 25'b00110010_01110000_10100010_0;
      patterns[12915] = 25'b00110010_01110001_10100011_0;
      patterns[12916] = 25'b00110010_01110010_10100100_0;
      patterns[12917] = 25'b00110010_01110011_10100101_0;
      patterns[12918] = 25'b00110010_01110100_10100110_0;
      patterns[12919] = 25'b00110010_01110101_10100111_0;
      patterns[12920] = 25'b00110010_01110110_10101000_0;
      patterns[12921] = 25'b00110010_01110111_10101001_0;
      patterns[12922] = 25'b00110010_01111000_10101010_0;
      patterns[12923] = 25'b00110010_01111001_10101011_0;
      patterns[12924] = 25'b00110010_01111010_10101100_0;
      patterns[12925] = 25'b00110010_01111011_10101101_0;
      patterns[12926] = 25'b00110010_01111100_10101110_0;
      patterns[12927] = 25'b00110010_01111101_10101111_0;
      patterns[12928] = 25'b00110010_01111110_10110000_0;
      patterns[12929] = 25'b00110010_01111111_10110001_0;
      patterns[12930] = 25'b00110010_10000000_10110010_0;
      patterns[12931] = 25'b00110010_10000001_10110011_0;
      patterns[12932] = 25'b00110010_10000010_10110100_0;
      patterns[12933] = 25'b00110010_10000011_10110101_0;
      patterns[12934] = 25'b00110010_10000100_10110110_0;
      patterns[12935] = 25'b00110010_10000101_10110111_0;
      patterns[12936] = 25'b00110010_10000110_10111000_0;
      patterns[12937] = 25'b00110010_10000111_10111001_0;
      patterns[12938] = 25'b00110010_10001000_10111010_0;
      patterns[12939] = 25'b00110010_10001001_10111011_0;
      patterns[12940] = 25'b00110010_10001010_10111100_0;
      patterns[12941] = 25'b00110010_10001011_10111101_0;
      patterns[12942] = 25'b00110010_10001100_10111110_0;
      patterns[12943] = 25'b00110010_10001101_10111111_0;
      patterns[12944] = 25'b00110010_10001110_11000000_0;
      patterns[12945] = 25'b00110010_10001111_11000001_0;
      patterns[12946] = 25'b00110010_10010000_11000010_0;
      patterns[12947] = 25'b00110010_10010001_11000011_0;
      patterns[12948] = 25'b00110010_10010010_11000100_0;
      patterns[12949] = 25'b00110010_10010011_11000101_0;
      patterns[12950] = 25'b00110010_10010100_11000110_0;
      patterns[12951] = 25'b00110010_10010101_11000111_0;
      patterns[12952] = 25'b00110010_10010110_11001000_0;
      patterns[12953] = 25'b00110010_10010111_11001001_0;
      patterns[12954] = 25'b00110010_10011000_11001010_0;
      patterns[12955] = 25'b00110010_10011001_11001011_0;
      patterns[12956] = 25'b00110010_10011010_11001100_0;
      patterns[12957] = 25'b00110010_10011011_11001101_0;
      patterns[12958] = 25'b00110010_10011100_11001110_0;
      patterns[12959] = 25'b00110010_10011101_11001111_0;
      patterns[12960] = 25'b00110010_10011110_11010000_0;
      patterns[12961] = 25'b00110010_10011111_11010001_0;
      patterns[12962] = 25'b00110010_10100000_11010010_0;
      patterns[12963] = 25'b00110010_10100001_11010011_0;
      patterns[12964] = 25'b00110010_10100010_11010100_0;
      patterns[12965] = 25'b00110010_10100011_11010101_0;
      patterns[12966] = 25'b00110010_10100100_11010110_0;
      patterns[12967] = 25'b00110010_10100101_11010111_0;
      patterns[12968] = 25'b00110010_10100110_11011000_0;
      patterns[12969] = 25'b00110010_10100111_11011001_0;
      patterns[12970] = 25'b00110010_10101000_11011010_0;
      patterns[12971] = 25'b00110010_10101001_11011011_0;
      patterns[12972] = 25'b00110010_10101010_11011100_0;
      patterns[12973] = 25'b00110010_10101011_11011101_0;
      patterns[12974] = 25'b00110010_10101100_11011110_0;
      patterns[12975] = 25'b00110010_10101101_11011111_0;
      patterns[12976] = 25'b00110010_10101110_11100000_0;
      patterns[12977] = 25'b00110010_10101111_11100001_0;
      patterns[12978] = 25'b00110010_10110000_11100010_0;
      patterns[12979] = 25'b00110010_10110001_11100011_0;
      patterns[12980] = 25'b00110010_10110010_11100100_0;
      patterns[12981] = 25'b00110010_10110011_11100101_0;
      patterns[12982] = 25'b00110010_10110100_11100110_0;
      patterns[12983] = 25'b00110010_10110101_11100111_0;
      patterns[12984] = 25'b00110010_10110110_11101000_0;
      patterns[12985] = 25'b00110010_10110111_11101001_0;
      patterns[12986] = 25'b00110010_10111000_11101010_0;
      patterns[12987] = 25'b00110010_10111001_11101011_0;
      patterns[12988] = 25'b00110010_10111010_11101100_0;
      patterns[12989] = 25'b00110010_10111011_11101101_0;
      patterns[12990] = 25'b00110010_10111100_11101110_0;
      patterns[12991] = 25'b00110010_10111101_11101111_0;
      patterns[12992] = 25'b00110010_10111110_11110000_0;
      patterns[12993] = 25'b00110010_10111111_11110001_0;
      patterns[12994] = 25'b00110010_11000000_11110010_0;
      patterns[12995] = 25'b00110010_11000001_11110011_0;
      patterns[12996] = 25'b00110010_11000010_11110100_0;
      patterns[12997] = 25'b00110010_11000011_11110101_0;
      patterns[12998] = 25'b00110010_11000100_11110110_0;
      patterns[12999] = 25'b00110010_11000101_11110111_0;
      patterns[13000] = 25'b00110010_11000110_11111000_0;
      patterns[13001] = 25'b00110010_11000111_11111001_0;
      patterns[13002] = 25'b00110010_11001000_11111010_0;
      patterns[13003] = 25'b00110010_11001001_11111011_0;
      patterns[13004] = 25'b00110010_11001010_11111100_0;
      patterns[13005] = 25'b00110010_11001011_11111101_0;
      patterns[13006] = 25'b00110010_11001100_11111110_0;
      patterns[13007] = 25'b00110010_11001101_11111111_0;
      patterns[13008] = 25'b00110010_11001110_00000000_1;
      patterns[13009] = 25'b00110010_11001111_00000001_1;
      patterns[13010] = 25'b00110010_11010000_00000010_1;
      patterns[13011] = 25'b00110010_11010001_00000011_1;
      patterns[13012] = 25'b00110010_11010010_00000100_1;
      patterns[13013] = 25'b00110010_11010011_00000101_1;
      patterns[13014] = 25'b00110010_11010100_00000110_1;
      patterns[13015] = 25'b00110010_11010101_00000111_1;
      patterns[13016] = 25'b00110010_11010110_00001000_1;
      patterns[13017] = 25'b00110010_11010111_00001001_1;
      patterns[13018] = 25'b00110010_11011000_00001010_1;
      patterns[13019] = 25'b00110010_11011001_00001011_1;
      patterns[13020] = 25'b00110010_11011010_00001100_1;
      patterns[13021] = 25'b00110010_11011011_00001101_1;
      patterns[13022] = 25'b00110010_11011100_00001110_1;
      patterns[13023] = 25'b00110010_11011101_00001111_1;
      patterns[13024] = 25'b00110010_11011110_00010000_1;
      patterns[13025] = 25'b00110010_11011111_00010001_1;
      patterns[13026] = 25'b00110010_11100000_00010010_1;
      patterns[13027] = 25'b00110010_11100001_00010011_1;
      patterns[13028] = 25'b00110010_11100010_00010100_1;
      patterns[13029] = 25'b00110010_11100011_00010101_1;
      patterns[13030] = 25'b00110010_11100100_00010110_1;
      patterns[13031] = 25'b00110010_11100101_00010111_1;
      patterns[13032] = 25'b00110010_11100110_00011000_1;
      patterns[13033] = 25'b00110010_11100111_00011001_1;
      patterns[13034] = 25'b00110010_11101000_00011010_1;
      patterns[13035] = 25'b00110010_11101001_00011011_1;
      patterns[13036] = 25'b00110010_11101010_00011100_1;
      patterns[13037] = 25'b00110010_11101011_00011101_1;
      patterns[13038] = 25'b00110010_11101100_00011110_1;
      patterns[13039] = 25'b00110010_11101101_00011111_1;
      patterns[13040] = 25'b00110010_11101110_00100000_1;
      patterns[13041] = 25'b00110010_11101111_00100001_1;
      patterns[13042] = 25'b00110010_11110000_00100010_1;
      patterns[13043] = 25'b00110010_11110001_00100011_1;
      patterns[13044] = 25'b00110010_11110010_00100100_1;
      patterns[13045] = 25'b00110010_11110011_00100101_1;
      patterns[13046] = 25'b00110010_11110100_00100110_1;
      patterns[13047] = 25'b00110010_11110101_00100111_1;
      patterns[13048] = 25'b00110010_11110110_00101000_1;
      patterns[13049] = 25'b00110010_11110111_00101001_1;
      patterns[13050] = 25'b00110010_11111000_00101010_1;
      patterns[13051] = 25'b00110010_11111001_00101011_1;
      patterns[13052] = 25'b00110010_11111010_00101100_1;
      patterns[13053] = 25'b00110010_11111011_00101101_1;
      patterns[13054] = 25'b00110010_11111100_00101110_1;
      patterns[13055] = 25'b00110010_11111101_00101111_1;
      patterns[13056] = 25'b00110010_11111110_00110000_1;
      patterns[13057] = 25'b00110010_11111111_00110001_1;
      patterns[13058] = 25'b00110011_00000000_00110011_0;
      patterns[13059] = 25'b00110011_00000001_00110100_0;
      patterns[13060] = 25'b00110011_00000010_00110101_0;
      patterns[13061] = 25'b00110011_00000011_00110110_0;
      patterns[13062] = 25'b00110011_00000100_00110111_0;
      patterns[13063] = 25'b00110011_00000101_00111000_0;
      patterns[13064] = 25'b00110011_00000110_00111001_0;
      patterns[13065] = 25'b00110011_00000111_00111010_0;
      patterns[13066] = 25'b00110011_00001000_00111011_0;
      patterns[13067] = 25'b00110011_00001001_00111100_0;
      patterns[13068] = 25'b00110011_00001010_00111101_0;
      patterns[13069] = 25'b00110011_00001011_00111110_0;
      patterns[13070] = 25'b00110011_00001100_00111111_0;
      patterns[13071] = 25'b00110011_00001101_01000000_0;
      patterns[13072] = 25'b00110011_00001110_01000001_0;
      patterns[13073] = 25'b00110011_00001111_01000010_0;
      patterns[13074] = 25'b00110011_00010000_01000011_0;
      patterns[13075] = 25'b00110011_00010001_01000100_0;
      patterns[13076] = 25'b00110011_00010010_01000101_0;
      patterns[13077] = 25'b00110011_00010011_01000110_0;
      patterns[13078] = 25'b00110011_00010100_01000111_0;
      patterns[13079] = 25'b00110011_00010101_01001000_0;
      patterns[13080] = 25'b00110011_00010110_01001001_0;
      patterns[13081] = 25'b00110011_00010111_01001010_0;
      patterns[13082] = 25'b00110011_00011000_01001011_0;
      patterns[13083] = 25'b00110011_00011001_01001100_0;
      patterns[13084] = 25'b00110011_00011010_01001101_0;
      patterns[13085] = 25'b00110011_00011011_01001110_0;
      patterns[13086] = 25'b00110011_00011100_01001111_0;
      patterns[13087] = 25'b00110011_00011101_01010000_0;
      patterns[13088] = 25'b00110011_00011110_01010001_0;
      patterns[13089] = 25'b00110011_00011111_01010010_0;
      patterns[13090] = 25'b00110011_00100000_01010011_0;
      patterns[13091] = 25'b00110011_00100001_01010100_0;
      patterns[13092] = 25'b00110011_00100010_01010101_0;
      patterns[13093] = 25'b00110011_00100011_01010110_0;
      patterns[13094] = 25'b00110011_00100100_01010111_0;
      patterns[13095] = 25'b00110011_00100101_01011000_0;
      patterns[13096] = 25'b00110011_00100110_01011001_0;
      patterns[13097] = 25'b00110011_00100111_01011010_0;
      patterns[13098] = 25'b00110011_00101000_01011011_0;
      patterns[13099] = 25'b00110011_00101001_01011100_0;
      patterns[13100] = 25'b00110011_00101010_01011101_0;
      patterns[13101] = 25'b00110011_00101011_01011110_0;
      patterns[13102] = 25'b00110011_00101100_01011111_0;
      patterns[13103] = 25'b00110011_00101101_01100000_0;
      patterns[13104] = 25'b00110011_00101110_01100001_0;
      patterns[13105] = 25'b00110011_00101111_01100010_0;
      patterns[13106] = 25'b00110011_00110000_01100011_0;
      patterns[13107] = 25'b00110011_00110001_01100100_0;
      patterns[13108] = 25'b00110011_00110010_01100101_0;
      patterns[13109] = 25'b00110011_00110011_01100110_0;
      patterns[13110] = 25'b00110011_00110100_01100111_0;
      patterns[13111] = 25'b00110011_00110101_01101000_0;
      patterns[13112] = 25'b00110011_00110110_01101001_0;
      patterns[13113] = 25'b00110011_00110111_01101010_0;
      patterns[13114] = 25'b00110011_00111000_01101011_0;
      patterns[13115] = 25'b00110011_00111001_01101100_0;
      patterns[13116] = 25'b00110011_00111010_01101101_0;
      patterns[13117] = 25'b00110011_00111011_01101110_0;
      patterns[13118] = 25'b00110011_00111100_01101111_0;
      patterns[13119] = 25'b00110011_00111101_01110000_0;
      patterns[13120] = 25'b00110011_00111110_01110001_0;
      patterns[13121] = 25'b00110011_00111111_01110010_0;
      patterns[13122] = 25'b00110011_01000000_01110011_0;
      patterns[13123] = 25'b00110011_01000001_01110100_0;
      patterns[13124] = 25'b00110011_01000010_01110101_0;
      patterns[13125] = 25'b00110011_01000011_01110110_0;
      patterns[13126] = 25'b00110011_01000100_01110111_0;
      patterns[13127] = 25'b00110011_01000101_01111000_0;
      patterns[13128] = 25'b00110011_01000110_01111001_0;
      patterns[13129] = 25'b00110011_01000111_01111010_0;
      patterns[13130] = 25'b00110011_01001000_01111011_0;
      patterns[13131] = 25'b00110011_01001001_01111100_0;
      patterns[13132] = 25'b00110011_01001010_01111101_0;
      patterns[13133] = 25'b00110011_01001011_01111110_0;
      patterns[13134] = 25'b00110011_01001100_01111111_0;
      patterns[13135] = 25'b00110011_01001101_10000000_0;
      patterns[13136] = 25'b00110011_01001110_10000001_0;
      patterns[13137] = 25'b00110011_01001111_10000010_0;
      patterns[13138] = 25'b00110011_01010000_10000011_0;
      patterns[13139] = 25'b00110011_01010001_10000100_0;
      patterns[13140] = 25'b00110011_01010010_10000101_0;
      patterns[13141] = 25'b00110011_01010011_10000110_0;
      patterns[13142] = 25'b00110011_01010100_10000111_0;
      patterns[13143] = 25'b00110011_01010101_10001000_0;
      patterns[13144] = 25'b00110011_01010110_10001001_0;
      patterns[13145] = 25'b00110011_01010111_10001010_0;
      patterns[13146] = 25'b00110011_01011000_10001011_0;
      patterns[13147] = 25'b00110011_01011001_10001100_0;
      patterns[13148] = 25'b00110011_01011010_10001101_0;
      patterns[13149] = 25'b00110011_01011011_10001110_0;
      patterns[13150] = 25'b00110011_01011100_10001111_0;
      patterns[13151] = 25'b00110011_01011101_10010000_0;
      patterns[13152] = 25'b00110011_01011110_10010001_0;
      patterns[13153] = 25'b00110011_01011111_10010010_0;
      patterns[13154] = 25'b00110011_01100000_10010011_0;
      patterns[13155] = 25'b00110011_01100001_10010100_0;
      patterns[13156] = 25'b00110011_01100010_10010101_0;
      patterns[13157] = 25'b00110011_01100011_10010110_0;
      patterns[13158] = 25'b00110011_01100100_10010111_0;
      patterns[13159] = 25'b00110011_01100101_10011000_0;
      patterns[13160] = 25'b00110011_01100110_10011001_0;
      patterns[13161] = 25'b00110011_01100111_10011010_0;
      patterns[13162] = 25'b00110011_01101000_10011011_0;
      patterns[13163] = 25'b00110011_01101001_10011100_0;
      patterns[13164] = 25'b00110011_01101010_10011101_0;
      patterns[13165] = 25'b00110011_01101011_10011110_0;
      patterns[13166] = 25'b00110011_01101100_10011111_0;
      patterns[13167] = 25'b00110011_01101101_10100000_0;
      patterns[13168] = 25'b00110011_01101110_10100001_0;
      patterns[13169] = 25'b00110011_01101111_10100010_0;
      patterns[13170] = 25'b00110011_01110000_10100011_0;
      patterns[13171] = 25'b00110011_01110001_10100100_0;
      patterns[13172] = 25'b00110011_01110010_10100101_0;
      patterns[13173] = 25'b00110011_01110011_10100110_0;
      patterns[13174] = 25'b00110011_01110100_10100111_0;
      patterns[13175] = 25'b00110011_01110101_10101000_0;
      patterns[13176] = 25'b00110011_01110110_10101001_0;
      patterns[13177] = 25'b00110011_01110111_10101010_0;
      patterns[13178] = 25'b00110011_01111000_10101011_0;
      patterns[13179] = 25'b00110011_01111001_10101100_0;
      patterns[13180] = 25'b00110011_01111010_10101101_0;
      patterns[13181] = 25'b00110011_01111011_10101110_0;
      patterns[13182] = 25'b00110011_01111100_10101111_0;
      patterns[13183] = 25'b00110011_01111101_10110000_0;
      patterns[13184] = 25'b00110011_01111110_10110001_0;
      patterns[13185] = 25'b00110011_01111111_10110010_0;
      patterns[13186] = 25'b00110011_10000000_10110011_0;
      patterns[13187] = 25'b00110011_10000001_10110100_0;
      patterns[13188] = 25'b00110011_10000010_10110101_0;
      patterns[13189] = 25'b00110011_10000011_10110110_0;
      patterns[13190] = 25'b00110011_10000100_10110111_0;
      patterns[13191] = 25'b00110011_10000101_10111000_0;
      patterns[13192] = 25'b00110011_10000110_10111001_0;
      patterns[13193] = 25'b00110011_10000111_10111010_0;
      patterns[13194] = 25'b00110011_10001000_10111011_0;
      patterns[13195] = 25'b00110011_10001001_10111100_0;
      patterns[13196] = 25'b00110011_10001010_10111101_0;
      patterns[13197] = 25'b00110011_10001011_10111110_0;
      patterns[13198] = 25'b00110011_10001100_10111111_0;
      patterns[13199] = 25'b00110011_10001101_11000000_0;
      patterns[13200] = 25'b00110011_10001110_11000001_0;
      patterns[13201] = 25'b00110011_10001111_11000010_0;
      patterns[13202] = 25'b00110011_10010000_11000011_0;
      patterns[13203] = 25'b00110011_10010001_11000100_0;
      patterns[13204] = 25'b00110011_10010010_11000101_0;
      patterns[13205] = 25'b00110011_10010011_11000110_0;
      patterns[13206] = 25'b00110011_10010100_11000111_0;
      patterns[13207] = 25'b00110011_10010101_11001000_0;
      patterns[13208] = 25'b00110011_10010110_11001001_0;
      patterns[13209] = 25'b00110011_10010111_11001010_0;
      patterns[13210] = 25'b00110011_10011000_11001011_0;
      patterns[13211] = 25'b00110011_10011001_11001100_0;
      patterns[13212] = 25'b00110011_10011010_11001101_0;
      patterns[13213] = 25'b00110011_10011011_11001110_0;
      patterns[13214] = 25'b00110011_10011100_11001111_0;
      patterns[13215] = 25'b00110011_10011101_11010000_0;
      patterns[13216] = 25'b00110011_10011110_11010001_0;
      patterns[13217] = 25'b00110011_10011111_11010010_0;
      patterns[13218] = 25'b00110011_10100000_11010011_0;
      patterns[13219] = 25'b00110011_10100001_11010100_0;
      patterns[13220] = 25'b00110011_10100010_11010101_0;
      patterns[13221] = 25'b00110011_10100011_11010110_0;
      patterns[13222] = 25'b00110011_10100100_11010111_0;
      patterns[13223] = 25'b00110011_10100101_11011000_0;
      patterns[13224] = 25'b00110011_10100110_11011001_0;
      patterns[13225] = 25'b00110011_10100111_11011010_0;
      patterns[13226] = 25'b00110011_10101000_11011011_0;
      patterns[13227] = 25'b00110011_10101001_11011100_0;
      patterns[13228] = 25'b00110011_10101010_11011101_0;
      patterns[13229] = 25'b00110011_10101011_11011110_0;
      patterns[13230] = 25'b00110011_10101100_11011111_0;
      patterns[13231] = 25'b00110011_10101101_11100000_0;
      patterns[13232] = 25'b00110011_10101110_11100001_0;
      patterns[13233] = 25'b00110011_10101111_11100010_0;
      patterns[13234] = 25'b00110011_10110000_11100011_0;
      patterns[13235] = 25'b00110011_10110001_11100100_0;
      patterns[13236] = 25'b00110011_10110010_11100101_0;
      patterns[13237] = 25'b00110011_10110011_11100110_0;
      patterns[13238] = 25'b00110011_10110100_11100111_0;
      patterns[13239] = 25'b00110011_10110101_11101000_0;
      patterns[13240] = 25'b00110011_10110110_11101001_0;
      patterns[13241] = 25'b00110011_10110111_11101010_0;
      patterns[13242] = 25'b00110011_10111000_11101011_0;
      patterns[13243] = 25'b00110011_10111001_11101100_0;
      patterns[13244] = 25'b00110011_10111010_11101101_0;
      patterns[13245] = 25'b00110011_10111011_11101110_0;
      patterns[13246] = 25'b00110011_10111100_11101111_0;
      patterns[13247] = 25'b00110011_10111101_11110000_0;
      patterns[13248] = 25'b00110011_10111110_11110001_0;
      patterns[13249] = 25'b00110011_10111111_11110010_0;
      patterns[13250] = 25'b00110011_11000000_11110011_0;
      patterns[13251] = 25'b00110011_11000001_11110100_0;
      patterns[13252] = 25'b00110011_11000010_11110101_0;
      patterns[13253] = 25'b00110011_11000011_11110110_0;
      patterns[13254] = 25'b00110011_11000100_11110111_0;
      patterns[13255] = 25'b00110011_11000101_11111000_0;
      patterns[13256] = 25'b00110011_11000110_11111001_0;
      patterns[13257] = 25'b00110011_11000111_11111010_0;
      patterns[13258] = 25'b00110011_11001000_11111011_0;
      patterns[13259] = 25'b00110011_11001001_11111100_0;
      patterns[13260] = 25'b00110011_11001010_11111101_0;
      patterns[13261] = 25'b00110011_11001011_11111110_0;
      patterns[13262] = 25'b00110011_11001100_11111111_0;
      patterns[13263] = 25'b00110011_11001101_00000000_1;
      patterns[13264] = 25'b00110011_11001110_00000001_1;
      patterns[13265] = 25'b00110011_11001111_00000010_1;
      patterns[13266] = 25'b00110011_11010000_00000011_1;
      patterns[13267] = 25'b00110011_11010001_00000100_1;
      patterns[13268] = 25'b00110011_11010010_00000101_1;
      patterns[13269] = 25'b00110011_11010011_00000110_1;
      patterns[13270] = 25'b00110011_11010100_00000111_1;
      patterns[13271] = 25'b00110011_11010101_00001000_1;
      patterns[13272] = 25'b00110011_11010110_00001001_1;
      patterns[13273] = 25'b00110011_11010111_00001010_1;
      patterns[13274] = 25'b00110011_11011000_00001011_1;
      patterns[13275] = 25'b00110011_11011001_00001100_1;
      patterns[13276] = 25'b00110011_11011010_00001101_1;
      patterns[13277] = 25'b00110011_11011011_00001110_1;
      patterns[13278] = 25'b00110011_11011100_00001111_1;
      patterns[13279] = 25'b00110011_11011101_00010000_1;
      patterns[13280] = 25'b00110011_11011110_00010001_1;
      patterns[13281] = 25'b00110011_11011111_00010010_1;
      patterns[13282] = 25'b00110011_11100000_00010011_1;
      patterns[13283] = 25'b00110011_11100001_00010100_1;
      patterns[13284] = 25'b00110011_11100010_00010101_1;
      patterns[13285] = 25'b00110011_11100011_00010110_1;
      patterns[13286] = 25'b00110011_11100100_00010111_1;
      patterns[13287] = 25'b00110011_11100101_00011000_1;
      patterns[13288] = 25'b00110011_11100110_00011001_1;
      patterns[13289] = 25'b00110011_11100111_00011010_1;
      patterns[13290] = 25'b00110011_11101000_00011011_1;
      patterns[13291] = 25'b00110011_11101001_00011100_1;
      patterns[13292] = 25'b00110011_11101010_00011101_1;
      patterns[13293] = 25'b00110011_11101011_00011110_1;
      patterns[13294] = 25'b00110011_11101100_00011111_1;
      patterns[13295] = 25'b00110011_11101101_00100000_1;
      patterns[13296] = 25'b00110011_11101110_00100001_1;
      patterns[13297] = 25'b00110011_11101111_00100010_1;
      patterns[13298] = 25'b00110011_11110000_00100011_1;
      patterns[13299] = 25'b00110011_11110001_00100100_1;
      patterns[13300] = 25'b00110011_11110010_00100101_1;
      patterns[13301] = 25'b00110011_11110011_00100110_1;
      patterns[13302] = 25'b00110011_11110100_00100111_1;
      patterns[13303] = 25'b00110011_11110101_00101000_1;
      patterns[13304] = 25'b00110011_11110110_00101001_1;
      patterns[13305] = 25'b00110011_11110111_00101010_1;
      patterns[13306] = 25'b00110011_11111000_00101011_1;
      patterns[13307] = 25'b00110011_11111001_00101100_1;
      patterns[13308] = 25'b00110011_11111010_00101101_1;
      patterns[13309] = 25'b00110011_11111011_00101110_1;
      patterns[13310] = 25'b00110011_11111100_00101111_1;
      patterns[13311] = 25'b00110011_11111101_00110000_1;
      patterns[13312] = 25'b00110011_11111110_00110001_1;
      patterns[13313] = 25'b00110011_11111111_00110010_1;
      patterns[13314] = 25'b00110100_00000000_00110100_0;
      patterns[13315] = 25'b00110100_00000001_00110101_0;
      patterns[13316] = 25'b00110100_00000010_00110110_0;
      patterns[13317] = 25'b00110100_00000011_00110111_0;
      patterns[13318] = 25'b00110100_00000100_00111000_0;
      patterns[13319] = 25'b00110100_00000101_00111001_0;
      patterns[13320] = 25'b00110100_00000110_00111010_0;
      patterns[13321] = 25'b00110100_00000111_00111011_0;
      patterns[13322] = 25'b00110100_00001000_00111100_0;
      patterns[13323] = 25'b00110100_00001001_00111101_0;
      patterns[13324] = 25'b00110100_00001010_00111110_0;
      patterns[13325] = 25'b00110100_00001011_00111111_0;
      patterns[13326] = 25'b00110100_00001100_01000000_0;
      patterns[13327] = 25'b00110100_00001101_01000001_0;
      patterns[13328] = 25'b00110100_00001110_01000010_0;
      patterns[13329] = 25'b00110100_00001111_01000011_0;
      patterns[13330] = 25'b00110100_00010000_01000100_0;
      patterns[13331] = 25'b00110100_00010001_01000101_0;
      patterns[13332] = 25'b00110100_00010010_01000110_0;
      patterns[13333] = 25'b00110100_00010011_01000111_0;
      patterns[13334] = 25'b00110100_00010100_01001000_0;
      patterns[13335] = 25'b00110100_00010101_01001001_0;
      patterns[13336] = 25'b00110100_00010110_01001010_0;
      patterns[13337] = 25'b00110100_00010111_01001011_0;
      patterns[13338] = 25'b00110100_00011000_01001100_0;
      patterns[13339] = 25'b00110100_00011001_01001101_0;
      patterns[13340] = 25'b00110100_00011010_01001110_0;
      patterns[13341] = 25'b00110100_00011011_01001111_0;
      patterns[13342] = 25'b00110100_00011100_01010000_0;
      patterns[13343] = 25'b00110100_00011101_01010001_0;
      patterns[13344] = 25'b00110100_00011110_01010010_0;
      patterns[13345] = 25'b00110100_00011111_01010011_0;
      patterns[13346] = 25'b00110100_00100000_01010100_0;
      patterns[13347] = 25'b00110100_00100001_01010101_0;
      patterns[13348] = 25'b00110100_00100010_01010110_0;
      patterns[13349] = 25'b00110100_00100011_01010111_0;
      patterns[13350] = 25'b00110100_00100100_01011000_0;
      patterns[13351] = 25'b00110100_00100101_01011001_0;
      patterns[13352] = 25'b00110100_00100110_01011010_0;
      patterns[13353] = 25'b00110100_00100111_01011011_0;
      patterns[13354] = 25'b00110100_00101000_01011100_0;
      patterns[13355] = 25'b00110100_00101001_01011101_0;
      patterns[13356] = 25'b00110100_00101010_01011110_0;
      patterns[13357] = 25'b00110100_00101011_01011111_0;
      patterns[13358] = 25'b00110100_00101100_01100000_0;
      patterns[13359] = 25'b00110100_00101101_01100001_0;
      patterns[13360] = 25'b00110100_00101110_01100010_0;
      patterns[13361] = 25'b00110100_00101111_01100011_0;
      patterns[13362] = 25'b00110100_00110000_01100100_0;
      patterns[13363] = 25'b00110100_00110001_01100101_0;
      patterns[13364] = 25'b00110100_00110010_01100110_0;
      patterns[13365] = 25'b00110100_00110011_01100111_0;
      patterns[13366] = 25'b00110100_00110100_01101000_0;
      patterns[13367] = 25'b00110100_00110101_01101001_0;
      patterns[13368] = 25'b00110100_00110110_01101010_0;
      patterns[13369] = 25'b00110100_00110111_01101011_0;
      patterns[13370] = 25'b00110100_00111000_01101100_0;
      patterns[13371] = 25'b00110100_00111001_01101101_0;
      patterns[13372] = 25'b00110100_00111010_01101110_0;
      patterns[13373] = 25'b00110100_00111011_01101111_0;
      patterns[13374] = 25'b00110100_00111100_01110000_0;
      patterns[13375] = 25'b00110100_00111101_01110001_0;
      patterns[13376] = 25'b00110100_00111110_01110010_0;
      patterns[13377] = 25'b00110100_00111111_01110011_0;
      patterns[13378] = 25'b00110100_01000000_01110100_0;
      patterns[13379] = 25'b00110100_01000001_01110101_0;
      patterns[13380] = 25'b00110100_01000010_01110110_0;
      patterns[13381] = 25'b00110100_01000011_01110111_0;
      patterns[13382] = 25'b00110100_01000100_01111000_0;
      patterns[13383] = 25'b00110100_01000101_01111001_0;
      patterns[13384] = 25'b00110100_01000110_01111010_0;
      patterns[13385] = 25'b00110100_01000111_01111011_0;
      patterns[13386] = 25'b00110100_01001000_01111100_0;
      patterns[13387] = 25'b00110100_01001001_01111101_0;
      patterns[13388] = 25'b00110100_01001010_01111110_0;
      patterns[13389] = 25'b00110100_01001011_01111111_0;
      patterns[13390] = 25'b00110100_01001100_10000000_0;
      patterns[13391] = 25'b00110100_01001101_10000001_0;
      patterns[13392] = 25'b00110100_01001110_10000010_0;
      patterns[13393] = 25'b00110100_01001111_10000011_0;
      patterns[13394] = 25'b00110100_01010000_10000100_0;
      patterns[13395] = 25'b00110100_01010001_10000101_0;
      patterns[13396] = 25'b00110100_01010010_10000110_0;
      patterns[13397] = 25'b00110100_01010011_10000111_0;
      patterns[13398] = 25'b00110100_01010100_10001000_0;
      patterns[13399] = 25'b00110100_01010101_10001001_0;
      patterns[13400] = 25'b00110100_01010110_10001010_0;
      patterns[13401] = 25'b00110100_01010111_10001011_0;
      patterns[13402] = 25'b00110100_01011000_10001100_0;
      patterns[13403] = 25'b00110100_01011001_10001101_0;
      patterns[13404] = 25'b00110100_01011010_10001110_0;
      patterns[13405] = 25'b00110100_01011011_10001111_0;
      patterns[13406] = 25'b00110100_01011100_10010000_0;
      patterns[13407] = 25'b00110100_01011101_10010001_0;
      patterns[13408] = 25'b00110100_01011110_10010010_0;
      patterns[13409] = 25'b00110100_01011111_10010011_0;
      patterns[13410] = 25'b00110100_01100000_10010100_0;
      patterns[13411] = 25'b00110100_01100001_10010101_0;
      patterns[13412] = 25'b00110100_01100010_10010110_0;
      patterns[13413] = 25'b00110100_01100011_10010111_0;
      patterns[13414] = 25'b00110100_01100100_10011000_0;
      patterns[13415] = 25'b00110100_01100101_10011001_0;
      patterns[13416] = 25'b00110100_01100110_10011010_0;
      patterns[13417] = 25'b00110100_01100111_10011011_0;
      patterns[13418] = 25'b00110100_01101000_10011100_0;
      patterns[13419] = 25'b00110100_01101001_10011101_0;
      patterns[13420] = 25'b00110100_01101010_10011110_0;
      patterns[13421] = 25'b00110100_01101011_10011111_0;
      patterns[13422] = 25'b00110100_01101100_10100000_0;
      patterns[13423] = 25'b00110100_01101101_10100001_0;
      patterns[13424] = 25'b00110100_01101110_10100010_0;
      patterns[13425] = 25'b00110100_01101111_10100011_0;
      patterns[13426] = 25'b00110100_01110000_10100100_0;
      patterns[13427] = 25'b00110100_01110001_10100101_0;
      patterns[13428] = 25'b00110100_01110010_10100110_0;
      patterns[13429] = 25'b00110100_01110011_10100111_0;
      patterns[13430] = 25'b00110100_01110100_10101000_0;
      patterns[13431] = 25'b00110100_01110101_10101001_0;
      patterns[13432] = 25'b00110100_01110110_10101010_0;
      patterns[13433] = 25'b00110100_01110111_10101011_0;
      patterns[13434] = 25'b00110100_01111000_10101100_0;
      patterns[13435] = 25'b00110100_01111001_10101101_0;
      patterns[13436] = 25'b00110100_01111010_10101110_0;
      patterns[13437] = 25'b00110100_01111011_10101111_0;
      patterns[13438] = 25'b00110100_01111100_10110000_0;
      patterns[13439] = 25'b00110100_01111101_10110001_0;
      patterns[13440] = 25'b00110100_01111110_10110010_0;
      patterns[13441] = 25'b00110100_01111111_10110011_0;
      patterns[13442] = 25'b00110100_10000000_10110100_0;
      patterns[13443] = 25'b00110100_10000001_10110101_0;
      patterns[13444] = 25'b00110100_10000010_10110110_0;
      patterns[13445] = 25'b00110100_10000011_10110111_0;
      patterns[13446] = 25'b00110100_10000100_10111000_0;
      patterns[13447] = 25'b00110100_10000101_10111001_0;
      patterns[13448] = 25'b00110100_10000110_10111010_0;
      patterns[13449] = 25'b00110100_10000111_10111011_0;
      patterns[13450] = 25'b00110100_10001000_10111100_0;
      patterns[13451] = 25'b00110100_10001001_10111101_0;
      patterns[13452] = 25'b00110100_10001010_10111110_0;
      patterns[13453] = 25'b00110100_10001011_10111111_0;
      patterns[13454] = 25'b00110100_10001100_11000000_0;
      patterns[13455] = 25'b00110100_10001101_11000001_0;
      patterns[13456] = 25'b00110100_10001110_11000010_0;
      patterns[13457] = 25'b00110100_10001111_11000011_0;
      patterns[13458] = 25'b00110100_10010000_11000100_0;
      patterns[13459] = 25'b00110100_10010001_11000101_0;
      patterns[13460] = 25'b00110100_10010010_11000110_0;
      patterns[13461] = 25'b00110100_10010011_11000111_0;
      patterns[13462] = 25'b00110100_10010100_11001000_0;
      patterns[13463] = 25'b00110100_10010101_11001001_0;
      patterns[13464] = 25'b00110100_10010110_11001010_0;
      patterns[13465] = 25'b00110100_10010111_11001011_0;
      patterns[13466] = 25'b00110100_10011000_11001100_0;
      patterns[13467] = 25'b00110100_10011001_11001101_0;
      patterns[13468] = 25'b00110100_10011010_11001110_0;
      patterns[13469] = 25'b00110100_10011011_11001111_0;
      patterns[13470] = 25'b00110100_10011100_11010000_0;
      patterns[13471] = 25'b00110100_10011101_11010001_0;
      patterns[13472] = 25'b00110100_10011110_11010010_0;
      patterns[13473] = 25'b00110100_10011111_11010011_0;
      patterns[13474] = 25'b00110100_10100000_11010100_0;
      patterns[13475] = 25'b00110100_10100001_11010101_0;
      patterns[13476] = 25'b00110100_10100010_11010110_0;
      patterns[13477] = 25'b00110100_10100011_11010111_0;
      patterns[13478] = 25'b00110100_10100100_11011000_0;
      patterns[13479] = 25'b00110100_10100101_11011001_0;
      patterns[13480] = 25'b00110100_10100110_11011010_0;
      patterns[13481] = 25'b00110100_10100111_11011011_0;
      patterns[13482] = 25'b00110100_10101000_11011100_0;
      patterns[13483] = 25'b00110100_10101001_11011101_0;
      patterns[13484] = 25'b00110100_10101010_11011110_0;
      patterns[13485] = 25'b00110100_10101011_11011111_0;
      patterns[13486] = 25'b00110100_10101100_11100000_0;
      patterns[13487] = 25'b00110100_10101101_11100001_0;
      patterns[13488] = 25'b00110100_10101110_11100010_0;
      patterns[13489] = 25'b00110100_10101111_11100011_0;
      patterns[13490] = 25'b00110100_10110000_11100100_0;
      patterns[13491] = 25'b00110100_10110001_11100101_0;
      patterns[13492] = 25'b00110100_10110010_11100110_0;
      patterns[13493] = 25'b00110100_10110011_11100111_0;
      patterns[13494] = 25'b00110100_10110100_11101000_0;
      patterns[13495] = 25'b00110100_10110101_11101001_0;
      patterns[13496] = 25'b00110100_10110110_11101010_0;
      patterns[13497] = 25'b00110100_10110111_11101011_0;
      patterns[13498] = 25'b00110100_10111000_11101100_0;
      patterns[13499] = 25'b00110100_10111001_11101101_0;
      patterns[13500] = 25'b00110100_10111010_11101110_0;
      patterns[13501] = 25'b00110100_10111011_11101111_0;
      patterns[13502] = 25'b00110100_10111100_11110000_0;
      patterns[13503] = 25'b00110100_10111101_11110001_0;
      patterns[13504] = 25'b00110100_10111110_11110010_0;
      patterns[13505] = 25'b00110100_10111111_11110011_0;
      patterns[13506] = 25'b00110100_11000000_11110100_0;
      patterns[13507] = 25'b00110100_11000001_11110101_0;
      patterns[13508] = 25'b00110100_11000010_11110110_0;
      patterns[13509] = 25'b00110100_11000011_11110111_0;
      patterns[13510] = 25'b00110100_11000100_11111000_0;
      patterns[13511] = 25'b00110100_11000101_11111001_0;
      patterns[13512] = 25'b00110100_11000110_11111010_0;
      patterns[13513] = 25'b00110100_11000111_11111011_0;
      patterns[13514] = 25'b00110100_11001000_11111100_0;
      patterns[13515] = 25'b00110100_11001001_11111101_0;
      patterns[13516] = 25'b00110100_11001010_11111110_0;
      patterns[13517] = 25'b00110100_11001011_11111111_0;
      patterns[13518] = 25'b00110100_11001100_00000000_1;
      patterns[13519] = 25'b00110100_11001101_00000001_1;
      patterns[13520] = 25'b00110100_11001110_00000010_1;
      patterns[13521] = 25'b00110100_11001111_00000011_1;
      patterns[13522] = 25'b00110100_11010000_00000100_1;
      patterns[13523] = 25'b00110100_11010001_00000101_1;
      patterns[13524] = 25'b00110100_11010010_00000110_1;
      patterns[13525] = 25'b00110100_11010011_00000111_1;
      patterns[13526] = 25'b00110100_11010100_00001000_1;
      patterns[13527] = 25'b00110100_11010101_00001001_1;
      patterns[13528] = 25'b00110100_11010110_00001010_1;
      patterns[13529] = 25'b00110100_11010111_00001011_1;
      patterns[13530] = 25'b00110100_11011000_00001100_1;
      patterns[13531] = 25'b00110100_11011001_00001101_1;
      patterns[13532] = 25'b00110100_11011010_00001110_1;
      patterns[13533] = 25'b00110100_11011011_00001111_1;
      patterns[13534] = 25'b00110100_11011100_00010000_1;
      patterns[13535] = 25'b00110100_11011101_00010001_1;
      patterns[13536] = 25'b00110100_11011110_00010010_1;
      patterns[13537] = 25'b00110100_11011111_00010011_1;
      patterns[13538] = 25'b00110100_11100000_00010100_1;
      patterns[13539] = 25'b00110100_11100001_00010101_1;
      patterns[13540] = 25'b00110100_11100010_00010110_1;
      patterns[13541] = 25'b00110100_11100011_00010111_1;
      patterns[13542] = 25'b00110100_11100100_00011000_1;
      patterns[13543] = 25'b00110100_11100101_00011001_1;
      patterns[13544] = 25'b00110100_11100110_00011010_1;
      patterns[13545] = 25'b00110100_11100111_00011011_1;
      patterns[13546] = 25'b00110100_11101000_00011100_1;
      patterns[13547] = 25'b00110100_11101001_00011101_1;
      patterns[13548] = 25'b00110100_11101010_00011110_1;
      patterns[13549] = 25'b00110100_11101011_00011111_1;
      patterns[13550] = 25'b00110100_11101100_00100000_1;
      patterns[13551] = 25'b00110100_11101101_00100001_1;
      patterns[13552] = 25'b00110100_11101110_00100010_1;
      patterns[13553] = 25'b00110100_11101111_00100011_1;
      patterns[13554] = 25'b00110100_11110000_00100100_1;
      patterns[13555] = 25'b00110100_11110001_00100101_1;
      patterns[13556] = 25'b00110100_11110010_00100110_1;
      patterns[13557] = 25'b00110100_11110011_00100111_1;
      patterns[13558] = 25'b00110100_11110100_00101000_1;
      patterns[13559] = 25'b00110100_11110101_00101001_1;
      patterns[13560] = 25'b00110100_11110110_00101010_1;
      patterns[13561] = 25'b00110100_11110111_00101011_1;
      patterns[13562] = 25'b00110100_11111000_00101100_1;
      patterns[13563] = 25'b00110100_11111001_00101101_1;
      patterns[13564] = 25'b00110100_11111010_00101110_1;
      patterns[13565] = 25'b00110100_11111011_00101111_1;
      patterns[13566] = 25'b00110100_11111100_00110000_1;
      patterns[13567] = 25'b00110100_11111101_00110001_1;
      patterns[13568] = 25'b00110100_11111110_00110010_1;
      patterns[13569] = 25'b00110100_11111111_00110011_1;
      patterns[13570] = 25'b00110101_00000000_00110101_0;
      patterns[13571] = 25'b00110101_00000001_00110110_0;
      patterns[13572] = 25'b00110101_00000010_00110111_0;
      patterns[13573] = 25'b00110101_00000011_00111000_0;
      patterns[13574] = 25'b00110101_00000100_00111001_0;
      patterns[13575] = 25'b00110101_00000101_00111010_0;
      patterns[13576] = 25'b00110101_00000110_00111011_0;
      patterns[13577] = 25'b00110101_00000111_00111100_0;
      patterns[13578] = 25'b00110101_00001000_00111101_0;
      patterns[13579] = 25'b00110101_00001001_00111110_0;
      patterns[13580] = 25'b00110101_00001010_00111111_0;
      patterns[13581] = 25'b00110101_00001011_01000000_0;
      patterns[13582] = 25'b00110101_00001100_01000001_0;
      patterns[13583] = 25'b00110101_00001101_01000010_0;
      patterns[13584] = 25'b00110101_00001110_01000011_0;
      patterns[13585] = 25'b00110101_00001111_01000100_0;
      patterns[13586] = 25'b00110101_00010000_01000101_0;
      patterns[13587] = 25'b00110101_00010001_01000110_0;
      patterns[13588] = 25'b00110101_00010010_01000111_0;
      patterns[13589] = 25'b00110101_00010011_01001000_0;
      patterns[13590] = 25'b00110101_00010100_01001001_0;
      patterns[13591] = 25'b00110101_00010101_01001010_0;
      patterns[13592] = 25'b00110101_00010110_01001011_0;
      patterns[13593] = 25'b00110101_00010111_01001100_0;
      patterns[13594] = 25'b00110101_00011000_01001101_0;
      patterns[13595] = 25'b00110101_00011001_01001110_0;
      patterns[13596] = 25'b00110101_00011010_01001111_0;
      patterns[13597] = 25'b00110101_00011011_01010000_0;
      patterns[13598] = 25'b00110101_00011100_01010001_0;
      patterns[13599] = 25'b00110101_00011101_01010010_0;
      patterns[13600] = 25'b00110101_00011110_01010011_0;
      patterns[13601] = 25'b00110101_00011111_01010100_0;
      patterns[13602] = 25'b00110101_00100000_01010101_0;
      patterns[13603] = 25'b00110101_00100001_01010110_0;
      patterns[13604] = 25'b00110101_00100010_01010111_0;
      patterns[13605] = 25'b00110101_00100011_01011000_0;
      patterns[13606] = 25'b00110101_00100100_01011001_0;
      patterns[13607] = 25'b00110101_00100101_01011010_0;
      patterns[13608] = 25'b00110101_00100110_01011011_0;
      patterns[13609] = 25'b00110101_00100111_01011100_0;
      patterns[13610] = 25'b00110101_00101000_01011101_0;
      patterns[13611] = 25'b00110101_00101001_01011110_0;
      patterns[13612] = 25'b00110101_00101010_01011111_0;
      patterns[13613] = 25'b00110101_00101011_01100000_0;
      patterns[13614] = 25'b00110101_00101100_01100001_0;
      patterns[13615] = 25'b00110101_00101101_01100010_0;
      patterns[13616] = 25'b00110101_00101110_01100011_0;
      patterns[13617] = 25'b00110101_00101111_01100100_0;
      patterns[13618] = 25'b00110101_00110000_01100101_0;
      patterns[13619] = 25'b00110101_00110001_01100110_0;
      patterns[13620] = 25'b00110101_00110010_01100111_0;
      patterns[13621] = 25'b00110101_00110011_01101000_0;
      patterns[13622] = 25'b00110101_00110100_01101001_0;
      patterns[13623] = 25'b00110101_00110101_01101010_0;
      patterns[13624] = 25'b00110101_00110110_01101011_0;
      patterns[13625] = 25'b00110101_00110111_01101100_0;
      patterns[13626] = 25'b00110101_00111000_01101101_0;
      patterns[13627] = 25'b00110101_00111001_01101110_0;
      patterns[13628] = 25'b00110101_00111010_01101111_0;
      patterns[13629] = 25'b00110101_00111011_01110000_0;
      patterns[13630] = 25'b00110101_00111100_01110001_0;
      patterns[13631] = 25'b00110101_00111101_01110010_0;
      patterns[13632] = 25'b00110101_00111110_01110011_0;
      patterns[13633] = 25'b00110101_00111111_01110100_0;
      patterns[13634] = 25'b00110101_01000000_01110101_0;
      patterns[13635] = 25'b00110101_01000001_01110110_0;
      patterns[13636] = 25'b00110101_01000010_01110111_0;
      patterns[13637] = 25'b00110101_01000011_01111000_0;
      patterns[13638] = 25'b00110101_01000100_01111001_0;
      patterns[13639] = 25'b00110101_01000101_01111010_0;
      patterns[13640] = 25'b00110101_01000110_01111011_0;
      patterns[13641] = 25'b00110101_01000111_01111100_0;
      patterns[13642] = 25'b00110101_01001000_01111101_0;
      patterns[13643] = 25'b00110101_01001001_01111110_0;
      patterns[13644] = 25'b00110101_01001010_01111111_0;
      patterns[13645] = 25'b00110101_01001011_10000000_0;
      patterns[13646] = 25'b00110101_01001100_10000001_0;
      patterns[13647] = 25'b00110101_01001101_10000010_0;
      patterns[13648] = 25'b00110101_01001110_10000011_0;
      patterns[13649] = 25'b00110101_01001111_10000100_0;
      patterns[13650] = 25'b00110101_01010000_10000101_0;
      patterns[13651] = 25'b00110101_01010001_10000110_0;
      patterns[13652] = 25'b00110101_01010010_10000111_0;
      patterns[13653] = 25'b00110101_01010011_10001000_0;
      patterns[13654] = 25'b00110101_01010100_10001001_0;
      patterns[13655] = 25'b00110101_01010101_10001010_0;
      patterns[13656] = 25'b00110101_01010110_10001011_0;
      patterns[13657] = 25'b00110101_01010111_10001100_0;
      patterns[13658] = 25'b00110101_01011000_10001101_0;
      patterns[13659] = 25'b00110101_01011001_10001110_0;
      patterns[13660] = 25'b00110101_01011010_10001111_0;
      patterns[13661] = 25'b00110101_01011011_10010000_0;
      patterns[13662] = 25'b00110101_01011100_10010001_0;
      patterns[13663] = 25'b00110101_01011101_10010010_0;
      patterns[13664] = 25'b00110101_01011110_10010011_0;
      patterns[13665] = 25'b00110101_01011111_10010100_0;
      patterns[13666] = 25'b00110101_01100000_10010101_0;
      patterns[13667] = 25'b00110101_01100001_10010110_0;
      patterns[13668] = 25'b00110101_01100010_10010111_0;
      patterns[13669] = 25'b00110101_01100011_10011000_0;
      patterns[13670] = 25'b00110101_01100100_10011001_0;
      patterns[13671] = 25'b00110101_01100101_10011010_0;
      patterns[13672] = 25'b00110101_01100110_10011011_0;
      patterns[13673] = 25'b00110101_01100111_10011100_0;
      patterns[13674] = 25'b00110101_01101000_10011101_0;
      patterns[13675] = 25'b00110101_01101001_10011110_0;
      patterns[13676] = 25'b00110101_01101010_10011111_0;
      patterns[13677] = 25'b00110101_01101011_10100000_0;
      patterns[13678] = 25'b00110101_01101100_10100001_0;
      patterns[13679] = 25'b00110101_01101101_10100010_0;
      patterns[13680] = 25'b00110101_01101110_10100011_0;
      patterns[13681] = 25'b00110101_01101111_10100100_0;
      patterns[13682] = 25'b00110101_01110000_10100101_0;
      patterns[13683] = 25'b00110101_01110001_10100110_0;
      patterns[13684] = 25'b00110101_01110010_10100111_0;
      patterns[13685] = 25'b00110101_01110011_10101000_0;
      patterns[13686] = 25'b00110101_01110100_10101001_0;
      patterns[13687] = 25'b00110101_01110101_10101010_0;
      patterns[13688] = 25'b00110101_01110110_10101011_0;
      patterns[13689] = 25'b00110101_01110111_10101100_0;
      patterns[13690] = 25'b00110101_01111000_10101101_0;
      patterns[13691] = 25'b00110101_01111001_10101110_0;
      patterns[13692] = 25'b00110101_01111010_10101111_0;
      patterns[13693] = 25'b00110101_01111011_10110000_0;
      patterns[13694] = 25'b00110101_01111100_10110001_0;
      patterns[13695] = 25'b00110101_01111101_10110010_0;
      patterns[13696] = 25'b00110101_01111110_10110011_0;
      patterns[13697] = 25'b00110101_01111111_10110100_0;
      patterns[13698] = 25'b00110101_10000000_10110101_0;
      patterns[13699] = 25'b00110101_10000001_10110110_0;
      patterns[13700] = 25'b00110101_10000010_10110111_0;
      patterns[13701] = 25'b00110101_10000011_10111000_0;
      patterns[13702] = 25'b00110101_10000100_10111001_0;
      patterns[13703] = 25'b00110101_10000101_10111010_0;
      patterns[13704] = 25'b00110101_10000110_10111011_0;
      patterns[13705] = 25'b00110101_10000111_10111100_0;
      patterns[13706] = 25'b00110101_10001000_10111101_0;
      patterns[13707] = 25'b00110101_10001001_10111110_0;
      patterns[13708] = 25'b00110101_10001010_10111111_0;
      patterns[13709] = 25'b00110101_10001011_11000000_0;
      patterns[13710] = 25'b00110101_10001100_11000001_0;
      patterns[13711] = 25'b00110101_10001101_11000010_0;
      patterns[13712] = 25'b00110101_10001110_11000011_0;
      patterns[13713] = 25'b00110101_10001111_11000100_0;
      patterns[13714] = 25'b00110101_10010000_11000101_0;
      patterns[13715] = 25'b00110101_10010001_11000110_0;
      patterns[13716] = 25'b00110101_10010010_11000111_0;
      patterns[13717] = 25'b00110101_10010011_11001000_0;
      patterns[13718] = 25'b00110101_10010100_11001001_0;
      patterns[13719] = 25'b00110101_10010101_11001010_0;
      patterns[13720] = 25'b00110101_10010110_11001011_0;
      patterns[13721] = 25'b00110101_10010111_11001100_0;
      patterns[13722] = 25'b00110101_10011000_11001101_0;
      patterns[13723] = 25'b00110101_10011001_11001110_0;
      patterns[13724] = 25'b00110101_10011010_11001111_0;
      patterns[13725] = 25'b00110101_10011011_11010000_0;
      patterns[13726] = 25'b00110101_10011100_11010001_0;
      patterns[13727] = 25'b00110101_10011101_11010010_0;
      patterns[13728] = 25'b00110101_10011110_11010011_0;
      patterns[13729] = 25'b00110101_10011111_11010100_0;
      patterns[13730] = 25'b00110101_10100000_11010101_0;
      patterns[13731] = 25'b00110101_10100001_11010110_0;
      patterns[13732] = 25'b00110101_10100010_11010111_0;
      patterns[13733] = 25'b00110101_10100011_11011000_0;
      patterns[13734] = 25'b00110101_10100100_11011001_0;
      patterns[13735] = 25'b00110101_10100101_11011010_0;
      patterns[13736] = 25'b00110101_10100110_11011011_0;
      patterns[13737] = 25'b00110101_10100111_11011100_0;
      patterns[13738] = 25'b00110101_10101000_11011101_0;
      patterns[13739] = 25'b00110101_10101001_11011110_0;
      patterns[13740] = 25'b00110101_10101010_11011111_0;
      patterns[13741] = 25'b00110101_10101011_11100000_0;
      patterns[13742] = 25'b00110101_10101100_11100001_0;
      patterns[13743] = 25'b00110101_10101101_11100010_0;
      patterns[13744] = 25'b00110101_10101110_11100011_0;
      patterns[13745] = 25'b00110101_10101111_11100100_0;
      patterns[13746] = 25'b00110101_10110000_11100101_0;
      patterns[13747] = 25'b00110101_10110001_11100110_0;
      patterns[13748] = 25'b00110101_10110010_11100111_0;
      patterns[13749] = 25'b00110101_10110011_11101000_0;
      patterns[13750] = 25'b00110101_10110100_11101001_0;
      patterns[13751] = 25'b00110101_10110101_11101010_0;
      patterns[13752] = 25'b00110101_10110110_11101011_0;
      patterns[13753] = 25'b00110101_10110111_11101100_0;
      patterns[13754] = 25'b00110101_10111000_11101101_0;
      patterns[13755] = 25'b00110101_10111001_11101110_0;
      patterns[13756] = 25'b00110101_10111010_11101111_0;
      patterns[13757] = 25'b00110101_10111011_11110000_0;
      patterns[13758] = 25'b00110101_10111100_11110001_0;
      patterns[13759] = 25'b00110101_10111101_11110010_0;
      patterns[13760] = 25'b00110101_10111110_11110011_0;
      patterns[13761] = 25'b00110101_10111111_11110100_0;
      patterns[13762] = 25'b00110101_11000000_11110101_0;
      patterns[13763] = 25'b00110101_11000001_11110110_0;
      patterns[13764] = 25'b00110101_11000010_11110111_0;
      patterns[13765] = 25'b00110101_11000011_11111000_0;
      patterns[13766] = 25'b00110101_11000100_11111001_0;
      patterns[13767] = 25'b00110101_11000101_11111010_0;
      patterns[13768] = 25'b00110101_11000110_11111011_0;
      patterns[13769] = 25'b00110101_11000111_11111100_0;
      patterns[13770] = 25'b00110101_11001000_11111101_0;
      patterns[13771] = 25'b00110101_11001001_11111110_0;
      patterns[13772] = 25'b00110101_11001010_11111111_0;
      patterns[13773] = 25'b00110101_11001011_00000000_1;
      patterns[13774] = 25'b00110101_11001100_00000001_1;
      patterns[13775] = 25'b00110101_11001101_00000010_1;
      patterns[13776] = 25'b00110101_11001110_00000011_1;
      patterns[13777] = 25'b00110101_11001111_00000100_1;
      patterns[13778] = 25'b00110101_11010000_00000101_1;
      patterns[13779] = 25'b00110101_11010001_00000110_1;
      patterns[13780] = 25'b00110101_11010010_00000111_1;
      patterns[13781] = 25'b00110101_11010011_00001000_1;
      patterns[13782] = 25'b00110101_11010100_00001001_1;
      patterns[13783] = 25'b00110101_11010101_00001010_1;
      patterns[13784] = 25'b00110101_11010110_00001011_1;
      patterns[13785] = 25'b00110101_11010111_00001100_1;
      patterns[13786] = 25'b00110101_11011000_00001101_1;
      patterns[13787] = 25'b00110101_11011001_00001110_1;
      patterns[13788] = 25'b00110101_11011010_00001111_1;
      patterns[13789] = 25'b00110101_11011011_00010000_1;
      patterns[13790] = 25'b00110101_11011100_00010001_1;
      patterns[13791] = 25'b00110101_11011101_00010010_1;
      patterns[13792] = 25'b00110101_11011110_00010011_1;
      patterns[13793] = 25'b00110101_11011111_00010100_1;
      patterns[13794] = 25'b00110101_11100000_00010101_1;
      patterns[13795] = 25'b00110101_11100001_00010110_1;
      patterns[13796] = 25'b00110101_11100010_00010111_1;
      patterns[13797] = 25'b00110101_11100011_00011000_1;
      patterns[13798] = 25'b00110101_11100100_00011001_1;
      patterns[13799] = 25'b00110101_11100101_00011010_1;
      patterns[13800] = 25'b00110101_11100110_00011011_1;
      patterns[13801] = 25'b00110101_11100111_00011100_1;
      patterns[13802] = 25'b00110101_11101000_00011101_1;
      patterns[13803] = 25'b00110101_11101001_00011110_1;
      patterns[13804] = 25'b00110101_11101010_00011111_1;
      patterns[13805] = 25'b00110101_11101011_00100000_1;
      patterns[13806] = 25'b00110101_11101100_00100001_1;
      patterns[13807] = 25'b00110101_11101101_00100010_1;
      patterns[13808] = 25'b00110101_11101110_00100011_1;
      patterns[13809] = 25'b00110101_11101111_00100100_1;
      patterns[13810] = 25'b00110101_11110000_00100101_1;
      patterns[13811] = 25'b00110101_11110001_00100110_1;
      patterns[13812] = 25'b00110101_11110010_00100111_1;
      patterns[13813] = 25'b00110101_11110011_00101000_1;
      patterns[13814] = 25'b00110101_11110100_00101001_1;
      patterns[13815] = 25'b00110101_11110101_00101010_1;
      patterns[13816] = 25'b00110101_11110110_00101011_1;
      patterns[13817] = 25'b00110101_11110111_00101100_1;
      patterns[13818] = 25'b00110101_11111000_00101101_1;
      patterns[13819] = 25'b00110101_11111001_00101110_1;
      patterns[13820] = 25'b00110101_11111010_00101111_1;
      patterns[13821] = 25'b00110101_11111011_00110000_1;
      patterns[13822] = 25'b00110101_11111100_00110001_1;
      patterns[13823] = 25'b00110101_11111101_00110010_1;
      patterns[13824] = 25'b00110101_11111110_00110011_1;
      patterns[13825] = 25'b00110101_11111111_00110100_1;
      patterns[13826] = 25'b00110110_00000000_00110110_0;
      patterns[13827] = 25'b00110110_00000001_00110111_0;
      patterns[13828] = 25'b00110110_00000010_00111000_0;
      patterns[13829] = 25'b00110110_00000011_00111001_0;
      patterns[13830] = 25'b00110110_00000100_00111010_0;
      patterns[13831] = 25'b00110110_00000101_00111011_0;
      patterns[13832] = 25'b00110110_00000110_00111100_0;
      patterns[13833] = 25'b00110110_00000111_00111101_0;
      patterns[13834] = 25'b00110110_00001000_00111110_0;
      patterns[13835] = 25'b00110110_00001001_00111111_0;
      patterns[13836] = 25'b00110110_00001010_01000000_0;
      patterns[13837] = 25'b00110110_00001011_01000001_0;
      patterns[13838] = 25'b00110110_00001100_01000010_0;
      patterns[13839] = 25'b00110110_00001101_01000011_0;
      patterns[13840] = 25'b00110110_00001110_01000100_0;
      patterns[13841] = 25'b00110110_00001111_01000101_0;
      patterns[13842] = 25'b00110110_00010000_01000110_0;
      patterns[13843] = 25'b00110110_00010001_01000111_0;
      patterns[13844] = 25'b00110110_00010010_01001000_0;
      patterns[13845] = 25'b00110110_00010011_01001001_0;
      patterns[13846] = 25'b00110110_00010100_01001010_0;
      patterns[13847] = 25'b00110110_00010101_01001011_0;
      patterns[13848] = 25'b00110110_00010110_01001100_0;
      patterns[13849] = 25'b00110110_00010111_01001101_0;
      patterns[13850] = 25'b00110110_00011000_01001110_0;
      patterns[13851] = 25'b00110110_00011001_01001111_0;
      patterns[13852] = 25'b00110110_00011010_01010000_0;
      patterns[13853] = 25'b00110110_00011011_01010001_0;
      patterns[13854] = 25'b00110110_00011100_01010010_0;
      patterns[13855] = 25'b00110110_00011101_01010011_0;
      patterns[13856] = 25'b00110110_00011110_01010100_0;
      patterns[13857] = 25'b00110110_00011111_01010101_0;
      patterns[13858] = 25'b00110110_00100000_01010110_0;
      patterns[13859] = 25'b00110110_00100001_01010111_0;
      patterns[13860] = 25'b00110110_00100010_01011000_0;
      patterns[13861] = 25'b00110110_00100011_01011001_0;
      patterns[13862] = 25'b00110110_00100100_01011010_0;
      patterns[13863] = 25'b00110110_00100101_01011011_0;
      patterns[13864] = 25'b00110110_00100110_01011100_0;
      patterns[13865] = 25'b00110110_00100111_01011101_0;
      patterns[13866] = 25'b00110110_00101000_01011110_0;
      patterns[13867] = 25'b00110110_00101001_01011111_0;
      patterns[13868] = 25'b00110110_00101010_01100000_0;
      patterns[13869] = 25'b00110110_00101011_01100001_0;
      patterns[13870] = 25'b00110110_00101100_01100010_0;
      patterns[13871] = 25'b00110110_00101101_01100011_0;
      patterns[13872] = 25'b00110110_00101110_01100100_0;
      patterns[13873] = 25'b00110110_00101111_01100101_0;
      patterns[13874] = 25'b00110110_00110000_01100110_0;
      patterns[13875] = 25'b00110110_00110001_01100111_0;
      patterns[13876] = 25'b00110110_00110010_01101000_0;
      patterns[13877] = 25'b00110110_00110011_01101001_0;
      patterns[13878] = 25'b00110110_00110100_01101010_0;
      patterns[13879] = 25'b00110110_00110101_01101011_0;
      patterns[13880] = 25'b00110110_00110110_01101100_0;
      patterns[13881] = 25'b00110110_00110111_01101101_0;
      patterns[13882] = 25'b00110110_00111000_01101110_0;
      patterns[13883] = 25'b00110110_00111001_01101111_0;
      patterns[13884] = 25'b00110110_00111010_01110000_0;
      patterns[13885] = 25'b00110110_00111011_01110001_0;
      patterns[13886] = 25'b00110110_00111100_01110010_0;
      patterns[13887] = 25'b00110110_00111101_01110011_0;
      patterns[13888] = 25'b00110110_00111110_01110100_0;
      patterns[13889] = 25'b00110110_00111111_01110101_0;
      patterns[13890] = 25'b00110110_01000000_01110110_0;
      patterns[13891] = 25'b00110110_01000001_01110111_0;
      patterns[13892] = 25'b00110110_01000010_01111000_0;
      patterns[13893] = 25'b00110110_01000011_01111001_0;
      patterns[13894] = 25'b00110110_01000100_01111010_0;
      patterns[13895] = 25'b00110110_01000101_01111011_0;
      patterns[13896] = 25'b00110110_01000110_01111100_0;
      patterns[13897] = 25'b00110110_01000111_01111101_0;
      patterns[13898] = 25'b00110110_01001000_01111110_0;
      patterns[13899] = 25'b00110110_01001001_01111111_0;
      patterns[13900] = 25'b00110110_01001010_10000000_0;
      patterns[13901] = 25'b00110110_01001011_10000001_0;
      patterns[13902] = 25'b00110110_01001100_10000010_0;
      patterns[13903] = 25'b00110110_01001101_10000011_0;
      patterns[13904] = 25'b00110110_01001110_10000100_0;
      patterns[13905] = 25'b00110110_01001111_10000101_0;
      patterns[13906] = 25'b00110110_01010000_10000110_0;
      patterns[13907] = 25'b00110110_01010001_10000111_0;
      patterns[13908] = 25'b00110110_01010010_10001000_0;
      patterns[13909] = 25'b00110110_01010011_10001001_0;
      patterns[13910] = 25'b00110110_01010100_10001010_0;
      patterns[13911] = 25'b00110110_01010101_10001011_0;
      patterns[13912] = 25'b00110110_01010110_10001100_0;
      patterns[13913] = 25'b00110110_01010111_10001101_0;
      patterns[13914] = 25'b00110110_01011000_10001110_0;
      patterns[13915] = 25'b00110110_01011001_10001111_0;
      patterns[13916] = 25'b00110110_01011010_10010000_0;
      patterns[13917] = 25'b00110110_01011011_10010001_0;
      patterns[13918] = 25'b00110110_01011100_10010010_0;
      patterns[13919] = 25'b00110110_01011101_10010011_0;
      patterns[13920] = 25'b00110110_01011110_10010100_0;
      patterns[13921] = 25'b00110110_01011111_10010101_0;
      patterns[13922] = 25'b00110110_01100000_10010110_0;
      patterns[13923] = 25'b00110110_01100001_10010111_0;
      patterns[13924] = 25'b00110110_01100010_10011000_0;
      patterns[13925] = 25'b00110110_01100011_10011001_0;
      patterns[13926] = 25'b00110110_01100100_10011010_0;
      patterns[13927] = 25'b00110110_01100101_10011011_0;
      patterns[13928] = 25'b00110110_01100110_10011100_0;
      patterns[13929] = 25'b00110110_01100111_10011101_0;
      patterns[13930] = 25'b00110110_01101000_10011110_0;
      patterns[13931] = 25'b00110110_01101001_10011111_0;
      patterns[13932] = 25'b00110110_01101010_10100000_0;
      patterns[13933] = 25'b00110110_01101011_10100001_0;
      patterns[13934] = 25'b00110110_01101100_10100010_0;
      patterns[13935] = 25'b00110110_01101101_10100011_0;
      patterns[13936] = 25'b00110110_01101110_10100100_0;
      patterns[13937] = 25'b00110110_01101111_10100101_0;
      patterns[13938] = 25'b00110110_01110000_10100110_0;
      patterns[13939] = 25'b00110110_01110001_10100111_0;
      patterns[13940] = 25'b00110110_01110010_10101000_0;
      patterns[13941] = 25'b00110110_01110011_10101001_0;
      patterns[13942] = 25'b00110110_01110100_10101010_0;
      patterns[13943] = 25'b00110110_01110101_10101011_0;
      patterns[13944] = 25'b00110110_01110110_10101100_0;
      patterns[13945] = 25'b00110110_01110111_10101101_0;
      patterns[13946] = 25'b00110110_01111000_10101110_0;
      patterns[13947] = 25'b00110110_01111001_10101111_0;
      patterns[13948] = 25'b00110110_01111010_10110000_0;
      patterns[13949] = 25'b00110110_01111011_10110001_0;
      patterns[13950] = 25'b00110110_01111100_10110010_0;
      patterns[13951] = 25'b00110110_01111101_10110011_0;
      patterns[13952] = 25'b00110110_01111110_10110100_0;
      patterns[13953] = 25'b00110110_01111111_10110101_0;
      patterns[13954] = 25'b00110110_10000000_10110110_0;
      patterns[13955] = 25'b00110110_10000001_10110111_0;
      patterns[13956] = 25'b00110110_10000010_10111000_0;
      patterns[13957] = 25'b00110110_10000011_10111001_0;
      patterns[13958] = 25'b00110110_10000100_10111010_0;
      patterns[13959] = 25'b00110110_10000101_10111011_0;
      patterns[13960] = 25'b00110110_10000110_10111100_0;
      patterns[13961] = 25'b00110110_10000111_10111101_0;
      patterns[13962] = 25'b00110110_10001000_10111110_0;
      patterns[13963] = 25'b00110110_10001001_10111111_0;
      patterns[13964] = 25'b00110110_10001010_11000000_0;
      patterns[13965] = 25'b00110110_10001011_11000001_0;
      patterns[13966] = 25'b00110110_10001100_11000010_0;
      patterns[13967] = 25'b00110110_10001101_11000011_0;
      patterns[13968] = 25'b00110110_10001110_11000100_0;
      patterns[13969] = 25'b00110110_10001111_11000101_0;
      patterns[13970] = 25'b00110110_10010000_11000110_0;
      patterns[13971] = 25'b00110110_10010001_11000111_0;
      patterns[13972] = 25'b00110110_10010010_11001000_0;
      patterns[13973] = 25'b00110110_10010011_11001001_0;
      patterns[13974] = 25'b00110110_10010100_11001010_0;
      patterns[13975] = 25'b00110110_10010101_11001011_0;
      patterns[13976] = 25'b00110110_10010110_11001100_0;
      patterns[13977] = 25'b00110110_10010111_11001101_0;
      patterns[13978] = 25'b00110110_10011000_11001110_0;
      patterns[13979] = 25'b00110110_10011001_11001111_0;
      patterns[13980] = 25'b00110110_10011010_11010000_0;
      patterns[13981] = 25'b00110110_10011011_11010001_0;
      patterns[13982] = 25'b00110110_10011100_11010010_0;
      patterns[13983] = 25'b00110110_10011101_11010011_0;
      patterns[13984] = 25'b00110110_10011110_11010100_0;
      patterns[13985] = 25'b00110110_10011111_11010101_0;
      patterns[13986] = 25'b00110110_10100000_11010110_0;
      patterns[13987] = 25'b00110110_10100001_11010111_0;
      patterns[13988] = 25'b00110110_10100010_11011000_0;
      patterns[13989] = 25'b00110110_10100011_11011001_0;
      patterns[13990] = 25'b00110110_10100100_11011010_0;
      patterns[13991] = 25'b00110110_10100101_11011011_0;
      patterns[13992] = 25'b00110110_10100110_11011100_0;
      patterns[13993] = 25'b00110110_10100111_11011101_0;
      patterns[13994] = 25'b00110110_10101000_11011110_0;
      patterns[13995] = 25'b00110110_10101001_11011111_0;
      patterns[13996] = 25'b00110110_10101010_11100000_0;
      patterns[13997] = 25'b00110110_10101011_11100001_0;
      patterns[13998] = 25'b00110110_10101100_11100010_0;
      patterns[13999] = 25'b00110110_10101101_11100011_0;
      patterns[14000] = 25'b00110110_10101110_11100100_0;
      patterns[14001] = 25'b00110110_10101111_11100101_0;
      patterns[14002] = 25'b00110110_10110000_11100110_0;
      patterns[14003] = 25'b00110110_10110001_11100111_0;
      patterns[14004] = 25'b00110110_10110010_11101000_0;
      patterns[14005] = 25'b00110110_10110011_11101001_0;
      patterns[14006] = 25'b00110110_10110100_11101010_0;
      patterns[14007] = 25'b00110110_10110101_11101011_0;
      patterns[14008] = 25'b00110110_10110110_11101100_0;
      patterns[14009] = 25'b00110110_10110111_11101101_0;
      patterns[14010] = 25'b00110110_10111000_11101110_0;
      patterns[14011] = 25'b00110110_10111001_11101111_0;
      patterns[14012] = 25'b00110110_10111010_11110000_0;
      patterns[14013] = 25'b00110110_10111011_11110001_0;
      patterns[14014] = 25'b00110110_10111100_11110010_0;
      patterns[14015] = 25'b00110110_10111101_11110011_0;
      patterns[14016] = 25'b00110110_10111110_11110100_0;
      patterns[14017] = 25'b00110110_10111111_11110101_0;
      patterns[14018] = 25'b00110110_11000000_11110110_0;
      patterns[14019] = 25'b00110110_11000001_11110111_0;
      patterns[14020] = 25'b00110110_11000010_11111000_0;
      patterns[14021] = 25'b00110110_11000011_11111001_0;
      patterns[14022] = 25'b00110110_11000100_11111010_0;
      patterns[14023] = 25'b00110110_11000101_11111011_0;
      patterns[14024] = 25'b00110110_11000110_11111100_0;
      patterns[14025] = 25'b00110110_11000111_11111101_0;
      patterns[14026] = 25'b00110110_11001000_11111110_0;
      patterns[14027] = 25'b00110110_11001001_11111111_0;
      patterns[14028] = 25'b00110110_11001010_00000000_1;
      patterns[14029] = 25'b00110110_11001011_00000001_1;
      patterns[14030] = 25'b00110110_11001100_00000010_1;
      patterns[14031] = 25'b00110110_11001101_00000011_1;
      patterns[14032] = 25'b00110110_11001110_00000100_1;
      patterns[14033] = 25'b00110110_11001111_00000101_1;
      patterns[14034] = 25'b00110110_11010000_00000110_1;
      patterns[14035] = 25'b00110110_11010001_00000111_1;
      patterns[14036] = 25'b00110110_11010010_00001000_1;
      patterns[14037] = 25'b00110110_11010011_00001001_1;
      patterns[14038] = 25'b00110110_11010100_00001010_1;
      patterns[14039] = 25'b00110110_11010101_00001011_1;
      patterns[14040] = 25'b00110110_11010110_00001100_1;
      patterns[14041] = 25'b00110110_11010111_00001101_1;
      patterns[14042] = 25'b00110110_11011000_00001110_1;
      patterns[14043] = 25'b00110110_11011001_00001111_1;
      patterns[14044] = 25'b00110110_11011010_00010000_1;
      patterns[14045] = 25'b00110110_11011011_00010001_1;
      patterns[14046] = 25'b00110110_11011100_00010010_1;
      patterns[14047] = 25'b00110110_11011101_00010011_1;
      patterns[14048] = 25'b00110110_11011110_00010100_1;
      patterns[14049] = 25'b00110110_11011111_00010101_1;
      patterns[14050] = 25'b00110110_11100000_00010110_1;
      patterns[14051] = 25'b00110110_11100001_00010111_1;
      patterns[14052] = 25'b00110110_11100010_00011000_1;
      patterns[14053] = 25'b00110110_11100011_00011001_1;
      patterns[14054] = 25'b00110110_11100100_00011010_1;
      patterns[14055] = 25'b00110110_11100101_00011011_1;
      patterns[14056] = 25'b00110110_11100110_00011100_1;
      patterns[14057] = 25'b00110110_11100111_00011101_1;
      patterns[14058] = 25'b00110110_11101000_00011110_1;
      patterns[14059] = 25'b00110110_11101001_00011111_1;
      patterns[14060] = 25'b00110110_11101010_00100000_1;
      patterns[14061] = 25'b00110110_11101011_00100001_1;
      patterns[14062] = 25'b00110110_11101100_00100010_1;
      patterns[14063] = 25'b00110110_11101101_00100011_1;
      patterns[14064] = 25'b00110110_11101110_00100100_1;
      patterns[14065] = 25'b00110110_11101111_00100101_1;
      patterns[14066] = 25'b00110110_11110000_00100110_1;
      patterns[14067] = 25'b00110110_11110001_00100111_1;
      patterns[14068] = 25'b00110110_11110010_00101000_1;
      patterns[14069] = 25'b00110110_11110011_00101001_1;
      patterns[14070] = 25'b00110110_11110100_00101010_1;
      patterns[14071] = 25'b00110110_11110101_00101011_1;
      patterns[14072] = 25'b00110110_11110110_00101100_1;
      patterns[14073] = 25'b00110110_11110111_00101101_1;
      patterns[14074] = 25'b00110110_11111000_00101110_1;
      patterns[14075] = 25'b00110110_11111001_00101111_1;
      patterns[14076] = 25'b00110110_11111010_00110000_1;
      patterns[14077] = 25'b00110110_11111011_00110001_1;
      patterns[14078] = 25'b00110110_11111100_00110010_1;
      patterns[14079] = 25'b00110110_11111101_00110011_1;
      patterns[14080] = 25'b00110110_11111110_00110100_1;
      patterns[14081] = 25'b00110110_11111111_00110101_1;
      patterns[14082] = 25'b00110111_00000000_00110111_0;
      patterns[14083] = 25'b00110111_00000001_00111000_0;
      patterns[14084] = 25'b00110111_00000010_00111001_0;
      patterns[14085] = 25'b00110111_00000011_00111010_0;
      patterns[14086] = 25'b00110111_00000100_00111011_0;
      patterns[14087] = 25'b00110111_00000101_00111100_0;
      patterns[14088] = 25'b00110111_00000110_00111101_0;
      patterns[14089] = 25'b00110111_00000111_00111110_0;
      patterns[14090] = 25'b00110111_00001000_00111111_0;
      patterns[14091] = 25'b00110111_00001001_01000000_0;
      patterns[14092] = 25'b00110111_00001010_01000001_0;
      patterns[14093] = 25'b00110111_00001011_01000010_0;
      patterns[14094] = 25'b00110111_00001100_01000011_0;
      patterns[14095] = 25'b00110111_00001101_01000100_0;
      patterns[14096] = 25'b00110111_00001110_01000101_0;
      patterns[14097] = 25'b00110111_00001111_01000110_0;
      patterns[14098] = 25'b00110111_00010000_01000111_0;
      patterns[14099] = 25'b00110111_00010001_01001000_0;
      patterns[14100] = 25'b00110111_00010010_01001001_0;
      patterns[14101] = 25'b00110111_00010011_01001010_0;
      patterns[14102] = 25'b00110111_00010100_01001011_0;
      patterns[14103] = 25'b00110111_00010101_01001100_0;
      patterns[14104] = 25'b00110111_00010110_01001101_0;
      patterns[14105] = 25'b00110111_00010111_01001110_0;
      patterns[14106] = 25'b00110111_00011000_01001111_0;
      patterns[14107] = 25'b00110111_00011001_01010000_0;
      patterns[14108] = 25'b00110111_00011010_01010001_0;
      patterns[14109] = 25'b00110111_00011011_01010010_0;
      patterns[14110] = 25'b00110111_00011100_01010011_0;
      patterns[14111] = 25'b00110111_00011101_01010100_0;
      patterns[14112] = 25'b00110111_00011110_01010101_0;
      patterns[14113] = 25'b00110111_00011111_01010110_0;
      patterns[14114] = 25'b00110111_00100000_01010111_0;
      patterns[14115] = 25'b00110111_00100001_01011000_0;
      patterns[14116] = 25'b00110111_00100010_01011001_0;
      patterns[14117] = 25'b00110111_00100011_01011010_0;
      patterns[14118] = 25'b00110111_00100100_01011011_0;
      patterns[14119] = 25'b00110111_00100101_01011100_0;
      patterns[14120] = 25'b00110111_00100110_01011101_0;
      patterns[14121] = 25'b00110111_00100111_01011110_0;
      patterns[14122] = 25'b00110111_00101000_01011111_0;
      patterns[14123] = 25'b00110111_00101001_01100000_0;
      patterns[14124] = 25'b00110111_00101010_01100001_0;
      patterns[14125] = 25'b00110111_00101011_01100010_0;
      patterns[14126] = 25'b00110111_00101100_01100011_0;
      patterns[14127] = 25'b00110111_00101101_01100100_0;
      patterns[14128] = 25'b00110111_00101110_01100101_0;
      patterns[14129] = 25'b00110111_00101111_01100110_0;
      patterns[14130] = 25'b00110111_00110000_01100111_0;
      patterns[14131] = 25'b00110111_00110001_01101000_0;
      patterns[14132] = 25'b00110111_00110010_01101001_0;
      patterns[14133] = 25'b00110111_00110011_01101010_0;
      patterns[14134] = 25'b00110111_00110100_01101011_0;
      patterns[14135] = 25'b00110111_00110101_01101100_0;
      patterns[14136] = 25'b00110111_00110110_01101101_0;
      patterns[14137] = 25'b00110111_00110111_01101110_0;
      patterns[14138] = 25'b00110111_00111000_01101111_0;
      patterns[14139] = 25'b00110111_00111001_01110000_0;
      patterns[14140] = 25'b00110111_00111010_01110001_0;
      patterns[14141] = 25'b00110111_00111011_01110010_0;
      patterns[14142] = 25'b00110111_00111100_01110011_0;
      patterns[14143] = 25'b00110111_00111101_01110100_0;
      patterns[14144] = 25'b00110111_00111110_01110101_0;
      patterns[14145] = 25'b00110111_00111111_01110110_0;
      patterns[14146] = 25'b00110111_01000000_01110111_0;
      patterns[14147] = 25'b00110111_01000001_01111000_0;
      patterns[14148] = 25'b00110111_01000010_01111001_0;
      patterns[14149] = 25'b00110111_01000011_01111010_0;
      patterns[14150] = 25'b00110111_01000100_01111011_0;
      patterns[14151] = 25'b00110111_01000101_01111100_0;
      patterns[14152] = 25'b00110111_01000110_01111101_0;
      patterns[14153] = 25'b00110111_01000111_01111110_0;
      patterns[14154] = 25'b00110111_01001000_01111111_0;
      patterns[14155] = 25'b00110111_01001001_10000000_0;
      patterns[14156] = 25'b00110111_01001010_10000001_0;
      patterns[14157] = 25'b00110111_01001011_10000010_0;
      patterns[14158] = 25'b00110111_01001100_10000011_0;
      patterns[14159] = 25'b00110111_01001101_10000100_0;
      patterns[14160] = 25'b00110111_01001110_10000101_0;
      patterns[14161] = 25'b00110111_01001111_10000110_0;
      patterns[14162] = 25'b00110111_01010000_10000111_0;
      patterns[14163] = 25'b00110111_01010001_10001000_0;
      patterns[14164] = 25'b00110111_01010010_10001001_0;
      patterns[14165] = 25'b00110111_01010011_10001010_0;
      patterns[14166] = 25'b00110111_01010100_10001011_0;
      patterns[14167] = 25'b00110111_01010101_10001100_0;
      patterns[14168] = 25'b00110111_01010110_10001101_0;
      patterns[14169] = 25'b00110111_01010111_10001110_0;
      patterns[14170] = 25'b00110111_01011000_10001111_0;
      patterns[14171] = 25'b00110111_01011001_10010000_0;
      patterns[14172] = 25'b00110111_01011010_10010001_0;
      patterns[14173] = 25'b00110111_01011011_10010010_0;
      patterns[14174] = 25'b00110111_01011100_10010011_0;
      patterns[14175] = 25'b00110111_01011101_10010100_0;
      patterns[14176] = 25'b00110111_01011110_10010101_0;
      patterns[14177] = 25'b00110111_01011111_10010110_0;
      patterns[14178] = 25'b00110111_01100000_10010111_0;
      patterns[14179] = 25'b00110111_01100001_10011000_0;
      patterns[14180] = 25'b00110111_01100010_10011001_0;
      patterns[14181] = 25'b00110111_01100011_10011010_0;
      patterns[14182] = 25'b00110111_01100100_10011011_0;
      patterns[14183] = 25'b00110111_01100101_10011100_0;
      patterns[14184] = 25'b00110111_01100110_10011101_0;
      patterns[14185] = 25'b00110111_01100111_10011110_0;
      patterns[14186] = 25'b00110111_01101000_10011111_0;
      patterns[14187] = 25'b00110111_01101001_10100000_0;
      patterns[14188] = 25'b00110111_01101010_10100001_0;
      patterns[14189] = 25'b00110111_01101011_10100010_0;
      patterns[14190] = 25'b00110111_01101100_10100011_0;
      patterns[14191] = 25'b00110111_01101101_10100100_0;
      patterns[14192] = 25'b00110111_01101110_10100101_0;
      patterns[14193] = 25'b00110111_01101111_10100110_0;
      patterns[14194] = 25'b00110111_01110000_10100111_0;
      patterns[14195] = 25'b00110111_01110001_10101000_0;
      patterns[14196] = 25'b00110111_01110010_10101001_0;
      patterns[14197] = 25'b00110111_01110011_10101010_0;
      patterns[14198] = 25'b00110111_01110100_10101011_0;
      patterns[14199] = 25'b00110111_01110101_10101100_0;
      patterns[14200] = 25'b00110111_01110110_10101101_0;
      patterns[14201] = 25'b00110111_01110111_10101110_0;
      patterns[14202] = 25'b00110111_01111000_10101111_0;
      patterns[14203] = 25'b00110111_01111001_10110000_0;
      patterns[14204] = 25'b00110111_01111010_10110001_0;
      patterns[14205] = 25'b00110111_01111011_10110010_0;
      patterns[14206] = 25'b00110111_01111100_10110011_0;
      patterns[14207] = 25'b00110111_01111101_10110100_0;
      patterns[14208] = 25'b00110111_01111110_10110101_0;
      patterns[14209] = 25'b00110111_01111111_10110110_0;
      patterns[14210] = 25'b00110111_10000000_10110111_0;
      patterns[14211] = 25'b00110111_10000001_10111000_0;
      patterns[14212] = 25'b00110111_10000010_10111001_0;
      patterns[14213] = 25'b00110111_10000011_10111010_0;
      patterns[14214] = 25'b00110111_10000100_10111011_0;
      patterns[14215] = 25'b00110111_10000101_10111100_0;
      patterns[14216] = 25'b00110111_10000110_10111101_0;
      patterns[14217] = 25'b00110111_10000111_10111110_0;
      patterns[14218] = 25'b00110111_10001000_10111111_0;
      patterns[14219] = 25'b00110111_10001001_11000000_0;
      patterns[14220] = 25'b00110111_10001010_11000001_0;
      patterns[14221] = 25'b00110111_10001011_11000010_0;
      patterns[14222] = 25'b00110111_10001100_11000011_0;
      patterns[14223] = 25'b00110111_10001101_11000100_0;
      patterns[14224] = 25'b00110111_10001110_11000101_0;
      patterns[14225] = 25'b00110111_10001111_11000110_0;
      patterns[14226] = 25'b00110111_10010000_11000111_0;
      patterns[14227] = 25'b00110111_10010001_11001000_0;
      patterns[14228] = 25'b00110111_10010010_11001001_0;
      patterns[14229] = 25'b00110111_10010011_11001010_0;
      patterns[14230] = 25'b00110111_10010100_11001011_0;
      patterns[14231] = 25'b00110111_10010101_11001100_0;
      patterns[14232] = 25'b00110111_10010110_11001101_0;
      patterns[14233] = 25'b00110111_10010111_11001110_0;
      patterns[14234] = 25'b00110111_10011000_11001111_0;
      patterns[14235] = 25'b00110111_10011001_11010000_0;
      patterns[14236] = 25'b00110111_10011010_11010001_0;
      patterns[14237] = 25'b00110111_10011011_11010010_0;
      patterns[14238] = 25'b00110111_10011100_11010011_0;
      patterns[14239] = 25'b00110111_10011101_11010100_0;
      patterns[14240] = 25'b00110111_10011110_11010101_0;
      patterns[14241] = 25'b00110111_10011111_11010110_0;
      patterns[14242] = 25'b00110111_10100000_11010111_0;
      patterns[14243] = 25'b00110111_10100001_11011000_0;
      patterns[14244] = 25'b00110111_10100010_11011001_0;
      patterns[14245] = 25'b00110111_10100011_11011010_0;
      patterns[14246] = 25'b00110111_10100100_11011011_0;
      patterns[14247] = 25'b00110111_10100101_11011100_0;
      patterns[14248] = 25'b00110111_10100110_11011101_0;
      patterns[14249] = 25'b00110111_10100111_11011110_0;
      patterns[14250] = 25'b00110111_10101000_11011111_0;
      patterns[14251] = 25'b00110111_10101001_11100000_0;
      patterns[14252] = 25'b00110111_10101010_11100001_0;
      patterns[14253] = 25'b00110111_10101011_11100010_0;
      patterns[14254] = 25'b00110111_10101100_11100011_0;
      patterns[14255] = 25'b00110111_10101101_11100100_0;
      patterns[14256] = 25'b00110111_10101110_11100101_0;
      patterns[14257] = 25'b00110111_10101111_11100110_0;
      patterns[14258] = 25'b00110111_10110000_11100111_0;
      patterns[14259] = 25'b00110111_10110001_11101000_0;
      patterns[14260] = 25'b00110111_10110010_11101001_0;
      patterns[14261] = 25'b00110111_10110011_11101010_0;
      patterns[14262] = 25'b00110111_10110100_11101011_0;
      patterns[14263] = 25'b00110111_10110101_11101100_0;
      patterns[14264] = 25'b00110111_10110110_11101101_0;
      patterns[14265] = 25'b00110111_10110111_11101110_0;
      patterns[14266] = 25'b00110111_10111000_11101111_0;
      patterns[14267] = 25'b00110111_10111001_11110000_0;
      patterns[14268] = 25'b00110111_10111010_11110001_0;
      patterns[14269] = 25'b00110111_10111011_11110010_0;
      patterns[14270] = 25'b00110111_10111100_11110011_0;
      patterns[14271] = 25'b00110111_10111101_11110100_0;
      patterns[14272] = 25'b00110111_10111110_11110101_0;
      patterns[14273] = 25'b00110111_10111111_11110110_0;
      patterns[14274] = 25'b00110111_11000000_11110111_0;
      patterns[14275] = 25'b00110111_11000001_11111000_0;
      patterns[14276] = 25'b00110111_11000010_11111001_0;
      patterns[14277] = 25'b00110111_11000011_11111010_0;
      patterns[14278] = 25'b00110111_11000100_11111011_0;
      patterns[14279] = 25'b00110111_11000101_11111100_0;
      patterns[14280] = 25'b00110111_11000110_11111101_0;
      patterns[14281] = 25'b00110111_11000111_11111110_0;
      patterns[14282] = 25'b00110111_11001000_11111111_0;
      patterns[14283] = 25'b00110111_11001001_00000000_1;
      patterns[14284] = 25'b00110111_11001010_00000001_1;
      patterns[14285] = 25'b00110111_11001011_00000010_1;
      patterns[14286] = 25'b00110111_11001100_00000011_1;
      patterns[14287] = 25'b00110111_11001101_00000100_1;
      patterns[14288] = 25'b00110111_11001110_00000101_1;
      patterns[14289] = 25'b00110111_11001111_00000110_1;
      patterns[14290] = 25'b00110111_11010000_00000111_1;
      patterns[14291] = 25'b00110111_11010001_00001000_1;
      patterns[14292] = 25'b00110111_11010010_00001001_1;
      patterns[14293] = 25'b00110111_11010011_00001010_1;
      patterns[14294] = 25'b00110111_11010100_00001011_1;
      patterns[14295] = 25'b00110111_11010101_00001100_1;
      patterns[14296] = 25'b00110111_11010110_00001101_1;
      patterns[14297] = 25'b00110111_11010111_00001110_1;
      patterns[14298] = 25'b00110111_11011000_00001111_1;
      patterns[14299] = 25'b00110111_11011001_00010000_1;
      patterns[14300] = 25'b00110111_11011010_00010001_1;
      patterns[14301] = 25'b00110111_11011011_00010010_1;
      patterns[14302] = 25'b00110111_11011100_00010011_1;
      patterns[14303] = 25'b00110111_11011101_00010100_1;
      patterns[14304] = 25'b00110111_11011110_00010101_1;
      patterns[14305] = 25'b00110111_11011111_00010110_1;
      patterns[14306] = 25'b00110111_11100000_00010111_1;
      patterns[14307] = 25'b00110111_11100001_00011000_1;
      patterns[14308] = 25'b00110111_11100010_00011001_1;
      patterns[14309] = 25'b00110111_11100011_00011010_1;
      patterns[14310] = 25'b00110111_11100100_00011011_1;
      patterns[14311] = 25'b00110111_11100101_00011100_1;
      patterns[14312] = 25'b00110111_11100110_00011101_1;
      patterns[14313] = 25'b00110111_11100111_00011110_1;
      patterns[14314] = 25'b00110111_11101000_00011111_1;
      patterns[14315] = 25'b00110111_11101001_00100000_1;
      patterns[14316] = 25'b00110111_11101010_00100001_1;
      patterns[14317] = 25'b00110111_11101011_00100010_1;
      patterns[14318] = 25'b00110111_11101100_00100011_1;
      patterns[14319] = 25'b00110111_11101101_00100100_1;
      patterns[14320] = 25'b00110111_11101110_00100101_1;
      patterns[14321] = 25'b00110111_11101111_00100110_1;
      patterns[14322] = 25'b00110111_11110000_00100111_1;
      patterns[14323] = 25'b00110111_11110001_00101000_1;
      patterns[14324] = 25'b00110111_11110010_00101001_1;
      patterns[14325] = 25'b00110111_11110011_00101010_1;
      patterns[14326] = 25'b00110111_11110100_00101011_1;
      patterns[14327] = 25'b00110111_11110101_00101100_1;
      patterns[14328] = 25'b00110111_11110110_00101101_1;
      patterns[14329] = 25'b00110111_11110111_00101110_1;
      patterns[14330] = 25'b00110111_11111000_00101111_1;
      patterns[14331] = 25'b00110111_11111001_00110000_1;
      patterns[14332] = 25'b00110111_11111010_00110001_1;
      patterns[14333] = 25'b00110111_11111011_00110010_1;
      patterns[14334] = 25'b00110111_11111100_00110011_1;
      patterns[14335] = 25'b00110111_11111101_00110100_1;
      patterns[14336] = 25'b00110111_11111110_00110101_1;
      patterns[14337] = 25'b00110111_11111111_00110110_1;
      patterns[14338] = 25'b00111000_00000000_00111000_0;
      patterns[14339] = 25'b00111000_00000001_00111001_0;
      patterns[14340] = 25'b00111000_00000010_00111010_0;
      patterns[14341] = 25'b00111000_00000011_00111011_0;
      patterns[14342] = 25'b00111000_00000100_00111100_0;
      patterns[14343] = 25'b00111000_00000101_00111101_0;
      patterns[14344] = 25'b00111000_00000110_00111110_0;
      patterns[14345] = 25'b00111000_00000111_00111111_0;
      patterns[14346] = 25'b00111000_00001000_01000000_0;
      patterns[14347] = 25'b00111000_00001001_01000001_0;
      patterns[14348] = 25'b00111000_00001010_01000010_0;
      patterns[14349] = 25'b00111000_00001011_01000011_0;
      patterns[14350] = 25'b00111000_00001100_01000100_0;
      patterns[14351] = 25'b00111000_00001101_01000101_0;
      patterns[14352] = 25'b00111000_00001110_01000110_0;
      patterns[14353] = 25'b00111000_00001111_01000111_0;
      patterns[14354] = 25'b00111000_00010000_01001000_0;
      patterns[14355] = 25'b00111000_00010001_01001001_0;
      patterns[14356] = 25'b00111000_00010010_01001010_0;
      patterns[14357] = 25'b00111000_00010011_01001011_0;
      patterns[14358] = 25'b00111000_00010100_01001100_0;
      patterns[14359] = 25'b00111000_00010101_01001101_0;
      patterns[14360] = 25'b00111000_00010110_01001110_0;
      patterns[14361] = 25'b00111000_00010111_01001111_0;
      patterns[14362] = 25'b00111000_00011000_01010000_0;
      patterns[14363] = 25'b00111000_00011001_01010001_0;
      patterns[14364] = 25'b00111000_00011010_01010010_0;
      patterns[14365] = 25'b00111000_00011011_01010011_0;
      patterns[14366] = 25'b00111000_00011100_01010100_0;
      patterns[14367] = 25'b00111000_00011101_01010101_0;
      patterns[14368] = 25'b00111000_00011110_01010110_0;
      patterns[14369] = 25'b00111000_00011111_01010111_0;
      patterns[14370] = 25'b00111000_00100000_01011000_0;
      patterns[14371] = 25'b00111000_00100001_01011001_0;
      patterns[14372] = 25'b00111000_00100010_01011010_0;
      patterns[14373] = 25'b00111000_00100011_01011011_0;
      patterns[14374] = 25'b00111000_00100100_01011100_0;
      patterns[14375] = 25'b00111000_00100101_01011101_0;
      patterns[14376] = 25'b00111000_00100110_01011110_0;
      patterns[14377] = 25'b00111000_00100111_01011111_0;
      patterns[14378] = 25'b00111000_00101000_01100000_0;
      patterns[14379] = 25'b00111000_00101001_01100001_0;
      patterns[14380] = 25'b00111000_00101010_01100010_0;
      patterns[14381] = 25'b00111000_00101011_01100011_0;
      patterns[14382] = 25'b00111000_00101100_01100100_0;
      patterns[14383] = 25'b00111000_00101101_01100101_0;
      patterns[14384] = 25'b00111000_00101110_01100110_0;
      patterns[14385] = 25'b00111000_00101111_01100111_0;
      patterns[14386] = 25'b00111000_00110000_01101000_0;
      patterns[14387] = 25'b00111000_00110001_01101001_0;
      patterns[14388] = 25'b00111000_00110010_01101010_0;
      patterns[14389] = 25'b00111000_00110011_01101011_0;
      patterns[14390] = 25'b00111000_00110100_01101100_0;
      patterns[14391] = 25'b00111000_00110101_01101101_0;
      patterns[14392] = 25'b00111000_00110110_01101110_0;
      patterns[14393] = 25'b00111000_00110111_01101111_0;
      patterns[14394] = 25'b00111000_00111000_01110000_0;
      patterns[14395] = 25'b00111000_00111001_01110001_0;
      patterns[14396] = 25'b00111000_00111010_01110010_0;
      patterns[14397] = 25'b00111000_00111011_01110011_0;
      patterns[14398] = 25'b00111000_00111100_01110100_0;
      patterns[14399] = 25'b00111000_00111101_01110101_0;
      patterns[14400] = 25'b00111000_00111110_01110110_0;
      patterns[14401] = 25'b00111000_00111111_01110111_0;
      patterns[14402] = 25'b00111000_01000000_01111000_0;
      patterns[14403] = 25'b00111000_01000001_01111001_0;
      patterns[14404] = 25'b00111000_01000010_01111010_0;
      patterns[14405] = 25'b00111000_01000011_01111011_0;
      patterns[14406] = 25'b00111000_01000100_01111100_0;
      patterns[14407] = 25'b00111000_01000101_01111101_0;
      patterns[14408] = 25'b00111000_01000110_01111110_0;
      patterns[14409] = 25'b00111000_01000111_01111111_0;
      patterns[14410] = 25'b00111000_01001000_10000000_0;
      patterns[14411] = 25'b00111000_01001001_10000001_0;
      patterns[14412] = 25'b00111000_01001010_10000010_0;
      patterns[14413] = 25'b00111000_01001011_10000011_0;
      patterns[14414] = 25'b00111000_01001100_10000100_0;
      patterns[14415] = 25'b00111000_01001101_10000101_0;
      patterns[14416] = 25'b00111000_01001110_10000110_0;
      patterns[14417] = 25'b00111000_01001111_10000111_0;
      patterns[14418] = 25'b00111000_01010000_10001000_0;
      patterns[14419] = 25'b00111000_01010001_10001001_0;
      patterns[14420] = 25'b00111000_01010010_10001010_0;
      patterns[14421] = 25'b00111000_01010011_10001011_0;
      patterns[14422] = 25'b00111000_01010100_10001100_0;
      patterns[14423] = 25'b00111000_01010101_10001101_0;
      patterns[14424] = 25'b00111000_01010110_10001110_0;
      patterns[14425] = 25'b00111000_01010111_10001111_0;
      patterns[14426] = 25'b00111000_01011000_10010000_0;
      patterns[14427] = 25'b00111000_01011001_10010001_0;
      patterns[14428] = 25'b00111000_01011010_10010010_0;
      patterns[14429] = 25'b00111000_01011011_10010011_0;
      patterns[14430] = 25'b00111000_01011100_10010100_0;
      patterns[14431] = 25'b00111000_01011101_10010101_0;
      patterns[14432] = 25'b00111000_01011110_10010110_0;
      patterns[14433] = 25'b00111000_01011111_10010111_0;
      patterns[14434] = 25'b00111000_01100000_10011000_0;
      patterns[14435] = 25'b00111000_01100001_10011001_0;
      patterns[14436] = 25'b00111000_01100010_10011010_0;
      patterns[14437] = 25'b00111000_01100011_10011011_0;
      patterns[14438] = 25'b00111000_01100100_10011100_0;
      patterns[14439] = 25'b00111000_01100101_10011101_0;
      patterns[14440] = 25'b00111000_01100110_10011110_0;
      patterns[14441] = 25'b00111000_01100111_10011111_0;
      patterns[14442] = 25'b00111000_01101000_10100000_0;
      patterns[14443] = 25'b00111000_01101001_10100001_0;
      patterns[14444] = 25'b00111000_01101010_10100010_0;
      patterns[14445] = 25'b00111000_01101011_10100011_0;
      patterns[14446] = 25'b00111000_01101100_10100100_0;
      patterns[14447] = 25'b00111000_01101101_10100101_0;
      patterns[14448] = 25'b00111000_01101110_10100110_0;
      patterns[14449] = 25'b00111000_01101111_10100111_0;
      patterns[14450] = 25'b00111000_01110000_10101000_0;
      patterns[14451] = 25'b00111000_01110001_10101001_0;
      patterns[14452] = 25'b00111000_01110010_10101010_0;
      patterns[14453] = 25'b00111000_01110011_10101011_0;
      patterns[14454] = 25'b00111000_01110100_10101100_0;
      patterns[14455] = 25'b00111000_01110101_10101101_0;
      patterns[14456] = 25'b00111000_01110110_10101110_0;
      patterns[14457] = 25'b00111000_01110111_10101111_0;
      patterns[14458] = 25'b00111000_01111000_10110000_0;
      patterns[14459] = 25'b00111000_01111001_10110001_0;
      patterns[14460] = 25'b00111000_01111010_10110010_0;
      patterns[14461] = 25'b00111000_01111011_10110011_0;
      patterns[14462] = 25'b00111000_01111100_10110100_0;
      patterns[14463] = 25'b00111000_01111101_10110101_0;
      patterns[14464] = 25'b00111000_01111110_10110110_0;
      patterns[14465] = 25'b00111000_01111111_10110111_0;
      patterns[14466] = 25'b00111000_10000000_10111000_0;
      patterns[14467] = 25'b00111000_10000001_10111001_0;
      patterns[14468] = 25'b00111000_10000010_10111010_0;
      patterns[14469] = 25'b00111000_10000011_10111011_0;
      patterns[14470] = 25'b00111000_10000100_10111100_0;
      patterns[14471] = 25'b00111000_10000101_10111101_0;
      patterns[14472] = 25'b00111000_10000110_10111110_0;
      patterns[14473] = 25'b00111000_10000111_10111111_0;
      patterns[14474] = 25'b00111000_10001000_11000000_0;
      patterns[14475] = 25'b00111000_10001001_11000001_0;
      patterns[14476] = 25'b00111000_10001010_11000010_0;
      patterns[14477] = 25'b00111000_10001011_11000011_0;
      patterns[14478] = 25'b00111000_10001100_11000100_0;
      patterns[14479] = 25'b00111000_10001101_11000101_0;
      patterns[14480] = 25'b00111000_10001110_11000110_0;
      patterns[14481] = 25'b00111000_10001111_11000111_0;
      patterns[14482] = 25'b00111000_10010000_11001000_0;
      patterns[14483] = 25'b00111000_10010001_11001001_0;
      patterns[14484] = 25'b00111000_10010010_11001010_0;
      patterns[14485] = 25'b00111000_10010011_11001011_0;
      patterns[14486] = 25'b00111000_10010100_11001100_0;
      patterns[14487] = 25'b00111000_10010101_11001101_0;
      patterns[14488] = 25'b00111000_10010110_11001110_0;
      patterns[14489] = 25'b00111000_10010111_11001111_0;
      patterns[14490] = 25'b00111000_10011000_11010000_0;
      patterns[14491] = 25'b00111000_10011001_11010001_0;
      patterns[14492] = 25'b00111000_10011010_11010010_0;
      patterns[14493] = 25'b00111000_10011011_11010011_0;
      patterns[14494] = 25'b00111000_10011100_11010100_0;
      patterns[14495] = 25'b00111000_10011101_11010101_0;
      patterns[14496] = 25'b00111000_10011110_11010110_0;
      patterns[14497] = 25'b00111000_10011111_11010111_0;
      patterns[14498] = 25'b00111000_10100000_11011000_0;
      patterns[14499] = 25'b00111000_10100001_11011001_0;
      patterns[14500] = 25'b00111000_10100010_11011010_0;
      patterns[14501] = 25'b00111000_10100011_11011011_0;
      patterns[14502] = 25'b00111000_10100100_11011100_0;
      patterns[14503] = 25'b00111000_10100101_11011101_0;
      patterns[14504] = 25'b00111000_10100110_11011110_0;
      patterns[14505] = 25'b00111000_10100111_11011111_0;
      patterns[14506] = 25'b00111000_10101000_11100000_0;
      patterns[14507] = 25'b00111000_10101001_11100001_0;
      patterns[14508] = 25'b00111000_10101010_11100010_0;
      patterns[14509] = 25'b00111000_10101011_11100011_0;
      patterns[14510] = 25'b00111000_10101100_11100100_0;
      patterns[14511] = 25'b00111000_10101101_11100101_0;
      patterns[14512] = 25'b00111000_10101110_11100110_0;
      patterns[14513] = 25'b00111000_10101111_11100111_0;
      patterns[14514] = 25'b00111000_10110000_11101000_0;
      patterns[14515] = 25'b00111000_10110001_11101001_0;
      patterns[14516] = 25'b00111000_10110010_11101010_0;
      patterns[14517] = 25'b00111000_10110011_11101011_0;
      patterns[14518] = 25'b00111000_10110100_11101100_0;
      patterns[14519] = 25'b00111000_10110101_11101101_0;
      patterns[14520] = 25'b00111000_10110110_11101110_0;
      patterns[14521] = 25'b00111000_10110111_11101111_0;
      patterns[14522] = 25'b00111000_10111000_11110000_0;
      patterns[14523] = 25'b00111000_10111001_11110001_0;
      patterns[14524] = 25'b00111000_10111010_11110010_0;
      patterns[14525] = 25'b00111000_10111011_11110011_0;
      patterns[14526] = 25'b00111000_10111100_11110100_0;
      patterns[14527] = 25'b00111000_10111101_11110101_0;
      patterns[14528] = 25'b00111000_10111110_11110110_0;
      patterns[14529] = 25'b00111000_10111111_11110111_0;
      patterns[14530] = 25'b00111000_11000000_11111000_0;
      patterns[14531] = 25'b00111000_11000001_11111001_0;
      patterns[14532] = 25'b00111000_11000010_11111010_0;
      patterns[14533] = 25'b00111000_11000011_11111011_0;
      patterns[14534] = 25'b00111000_11000100_11111100_0;
      patterns[14535] = 25'b00111000_11000101_11111101_0;
      patterns[14536] = 25'b00111000_11000110_11111110_0;
      patterns[14537] = 25'b00111000_11000111_11111111_0;
      patterns[14538] = 25'b00111000_11001000_00000000_1;
      patterns[14539] = 25'b00111000_11001001_00000001_1;
      patterns[14540] = 25'b00111000_11001010_00000010_1;
      patterns[14541] = 25'b00111000_11001011_00000011_1;
      patterns[14542] = 25'b00111000_11001100_00000100_1;
      patterns[14543] = 25'b00111000_11001101_00000101_1;
      patterns[14544] = 25'b00111000_11001110_00000110_1;
      patterns[14545] = 25'b00111000_11001111_00000111_1;
      patterns[14546] = 25'b00111000_11010000_00001000_1;
      patterns[14547] = 25'b00111000_11010001_00001001_1;
      patterns[14548] = 25'b00111000_11010010_00001010_1;
      patterns[14549] = 25'b00111000_11010011_00001011_1;
      patterns[14550] = 25'b00111000_11010100_00001100_1;
      patterns[14551] = 25'b00111000_11010101_00001101_1;
      patterns[14552] = 25'b00111000_11010110_00001110_1;
      patterns[14553] = 25'b00111000_11010111_00001111_1;
      patterns[14554] = 25'b00111000_11011000_00010000_1;
      patterns[14555] = 25'b00111000_11011001_00010001_1;
      patterns[14556] = 25'b00111000_11011010_00010010_1;
      patterns[14557] = 25'b00111000_11011011_00010011_1;
      patterns[14558] = 25'b00111000_11011100_00010100_1;
      patterns[14559] = 25'b00111000_11011101_00010101_1;
      patterns[14560] = 25'b00111000_11011110_00010110_1;
      patterns[14561] = 25'b00111000_11011111_00010111_1;
      patterns[14562] = 25'b00111000_11100000_00011000_1;
      patterns[14563] = 25'b00111000_11100001_00011001_1;
      patterns[14564] = 25'b00111000_11100010_00011010_1;
      patterns[14565] = 25'b00111000_11100011_00011011_1;
      patterns[14566] = 25'b00111000_11100100_00011100_1;
      patterns[14567] = 25'b00111000_11100101_00011101_1;
      patterns[14568] = 25'b00111000_11100110_00011110_1;
      patterns[14569] = 25'b00111000_11100111_00011111_1;
      patterns[14570] = 25'b00111000_11101000_00100000_1;
      patterns[14571] = 25'b00111000_11101001_00100001_1;
      patterns[14572] = 25'b00111000_11101010_00100010_1;
      patterns[14573] = 25'b00111000_11101011_00100011_1;
      patterns[14574] = 25'b00111000_11101100_00100100_1;
      patterns[14575] = 25'b00111000_11101101_00100101_1;
      patterns[14576] = 25'b00111000_11101110_00100110_1;
      patterns[14577] = 25'b00111000_11101111_00100111_1;
      patterns[14578] = 25'b00111000_11110000_00101000_1;
      patterns[14579] = 25'b00111000_11110001_00101001_1;
      patterns[14580] = 25'b00111000_11110010_00101010_1;
      patterns[14581] = 25'b00111000_11110011_00101011_1;
      patterns[14582] = 25'b00111000_11110100_00101100_1;
      patterns[14583] = 25'b00111000_11110101_00101101_1;
      patterns[14584] = 25'b00111000_11110110_00101110_1;
      patterns[14585] = 25'b00111000_11110111_00101111_1;
      patterns[14586] = 25'b00111000_11111000_00110000_1;
      patterns[14587] = 25'b00111000_11111001_00110001_1;
      patterns[14588] = 25'b00111000_11111010_00110010_1;
      patterns[14589] = 25'b00111000_11111011_00110011_1;
      patterns[14590] = 25'b00111000_11111100_00110100_1;
      patterns[14591] = 25'b00111000_11111101_00110101_1;
      patterns[14592] = 25'b00111000_11111110_00110110_1;
      patterns[14593] = 25'b00111000_11111111_00110111_1;
      patterns[14594] = 25'b00111001_00000000_00111001_0;
      patterns[14595] = 25'b00111001_00000001_00111010_0;
      patterns[14596] = 25'b00111001_00000010_00111011_0;
      patterns[14597] = 25'b00111001_00000011_00111100_0;
      patterns[14598] = 25'b00111001_00000100_00111101_0;
      patterns[14599] = 25'b00111001_00000101_00111110_0;
      patterns[14600] = 25'b00111001_00000110_00111111_0;
      patterns[14601] = 25'b00111001_00000111_01000000_0;
      patterns[14602] = 25'b00111001_00001000_01000001_0;
      patterns[14603] = 25'b00111001_00001001_01000010_0;
      patterns[14604] = 25'b00111001_00001010_01000011_0;
      patterns[14605] = 25'b00111001_00001011_01000100_0;
      patterns[14606] = 25'b00111001_00001100_01000101_0;
      patterns[14607] = 25'b00111001_00001101_01000110_0;
      patterns[14608] = 25'b00111001_00001110_01000111_0;
      patterns[14609] = 25'b00111001_00001111_01001000_0;
      patterns[14610] = 25'b00111001_00010000_01001001_0;
      patterns[14611] = 25'b00111001_00010001_01001010_0;
      patterns[14612] = 25'b00111001_00010010_01001011_0;
      patterns[14613] = 25'b00111001_00010011_01001100_0;
      patterns[14614] = 25'b00111001_00010100_01001101_0;
      patterns[14615] = 25'b00111001_00010101_01001110_0;
      patterns[14616] = 25'b00111001_00010110_01001111_0;
      patterns[14617] = 25'b00111001_00010111_01010000_0;
      patterns[14618] = 25'b00111001_00011000_01010001_0;
      patterns[14619] = 25'b00111001_00011001_01010010_0;
      patterns[14620] = 25'b00111001_00011010_01010011_0;
      patterns[14621] = 25'b00111001_00011011_01010100_0;
      patterns[14622] = 25'b00111001_00011100_01010101_0;
      patterns[14623] = 25'b00111001_00011101_01010110_0;
      patterns[14624] = 25'b00111001_00011110_01010111_0;
      patterns[14625] = 25'b00111001_00011111_01011000_0;
      patterns[14626] = 25'b00111001_00100000_01011001_0;
      patterns[14627] = 25'b00111001_00100001_01011010_0;
      patterns[14628] = 25'b00111001_00100010_01011011_0;
      patterns[14629] = 25'b00111001_00100011_01011100_0;
      patterns[14630] = 25'b00111001_00100100_01011101_0;
      patterns[14631] = 25'b00111001_00100101_01011110_0;
      patterns[14632] = 25'b00111001_00100110_01011111_0;
      patterns[14633] = 25'b00111001_00100111_01100000_0;
      patterns[14634] = 25'b00111001_00101000_01100001_0;
      patterns[14635] = 25'b00111001_00101001_01100010_0;
      patterns[14636] = 25'b00111001_00101010_01100011_0;
      patterns[14637] = 25'b00111001_00101011_01100100_0;
      patterns[14638] = 25'b00111001_00101100_01100101_0;
      patterns[14639] = 25'b00111001_00101101_01100110_0;
      patterns[14640] = 25'b00111001_00101110_01100111_0;
      patterns[14641] = 25'b00111001_00101111_01101000_0;
      patterns[14642] = 25'b00111001_00110000_01101001_0;
      patterns[14643] = 25'b00111001_00110001_01101010_0;
      patterns[14644] = 25'b00111001_00110010_01101011_0;
      patterns[14645] = 25'b00111001_00110011_01101100_0;
      patterns[14646] = 25'b00111001_00110100_01101101_0;
      patterns[14647] = 25'b00111001_00110101_01101110_0;
      patterns[14648] = 25'b00111001_00110110_01101111_0;
      patterns[14649] = 25'b00111001_00110111_01110000_0;
      patterns[14650] = 25'b00111001_00111000_01110001_0;
      patterns[14651] = 25'b00111001_00111001_01110010_0;
      patterns[14652] = 25'b00111001_00111010_01110011_0;
      patterns[14653] = 25'b00111001_00111011_01110100_0;
      patterns[14654] = 25'b00111001_00111100_01110101_0;
      patterns[14655] = 25'b00111001_00111101_01110110_0;
      patterns[14656] = 25'b00111001_00111110_01110111_0;
      patterns[14657] = 25'b00111001_00111111_01111000_0;
      patterns[14658] = 25'b00111001_01000000_01111001_0;
      patterns[14659] = 25'b00111001_01000001_01111010_0;
      patterns[14660] = 25'b00111001_01000010_01111011_0;
      patterns[14661] = 25'b00111001_01000011_01111100_0;
      patterns[14662] = 25'b00111001_01000100_01111101_0;
      patterns[14663] = 25'b00111001_01000101_01111110_0;
      patterns[14664] = 25'b00111001_01000110_01111111_0;
      patterns[14665] = 25'b00111001_01000111_10000000_0;
      patterns[14666] = 25'b00111001_01001000_10000001_0;
      patterns[14667] = 25'b00111001_01001001_10000010_0;
      patterns[14668] = 25'b00111001_01001010_10000011_0;
      patterns[14669] = 25'b00111001_01001011_10000100_0;
      patterns[14670] = 25'b00111001_01001100_10000101_0;
      patterns[14671] = 25'b00111001_01001101_10000110_0;
      patterns[14672] = 25'b00111001_01001110_10000111_0;
      patterns[14673] = 25'b00111001_01001111_10001000_0;
      patterns[14674] = 25'b00111001_01010000_10001001_0;
      patterns[14675] = 25'b00111001_01010001_10001010_0;
      patterns[14676] = 25'b00111001_01010010_10001011_0;
      patterns[14677] = 25'b00111001_01010011_10001100_0;
      patterns[14678] = 25'b00111001_01010100_10001101_0;
      patterns[14679] = 25'b00111001_01010101_10001110_0;
      patterns[14680] = 25'b00111001_01010110_10001111_0;
      patterns[14681] = 25'b00111001_01010111_10010000_0;
      patterns[14682] = 25'b00111001_01011000_10010001_0;
      patterns[14683] = 25'b00111001_01011001_10010010_0;
      patterns[14684] = 25'b00111001_01011010_10010011_0;
      patterns[14685] = 25'b00111001_01011011_10010100_0;
      patterns[14686] = 25'b00111001_01011100_10010101_0;
      patterns[14687] = 25'b00111001_01011101_10010110_0;
      patterns[14688] = 25'b00111001_01011110_10010111_0;
      patterns[14689] = 25'b00111001_01011111_10011000_0;
      patterns[14690] = 25'b00111001_01100000_10011001_0;
      patterns[14691] = 25'b00111001_01100001_10011010_0;
      patterns[14692] = 25'b00111001_01100010_10011011_0;
      patterns[14693] = 25'b00111001_01100011_10011100_0;
      patterns[14694] = 25'b00111001_01100100_10011101_0;
      patterns[14695] = 25'b00111001_01100101_10011110_0;
      patterns[14696] = 25'b00111001_01100110_10011111_0;
      patterns[14697] = 25'b00111001_01100111_10100000_0;
      patterns[14698] = 25'b00111001_01101000_10100001_0;
      patterns[14699] = 25'b00111001_01101001_10100010_0;
      patterns[14700] = 25'b00111001_01101010_10100011_0;
      patterns[14701] = 25'b00111001_01101011_10100100_0;
      patterns[14702] = 25'b00111001_01101100_10100101_0;
      patterns[14703] = 25'b00111001_01101101_10100110_0;
      patterns[14704] = 25'b00111001_01101110_10100111_0;
      patterns[14705] = 25'b00111001_01101111_10101000_0;
      patterns[14706] = 25'b00111001_01110000_10101001_0;
      patterns[14707] = 25'b00111001_01110001_10101010_0;
      patterns[14708] = 25'b00111001_01110010_10101011_0;
      patterns[14709] = 25'b00111001_01110011_10101100_0;
      patterns[14710] = 25'b00111001_01110100_10101101_0;
      patterns[14711] = 25'b00111001_01110101_10101110_0;
      patterns[14712] = 25'b00111001_01110110_10101111_0;
      patterns[14713] = 25'b00111001_01110111_10110000_0;
      patterns[14714] = 25'b00111001_01111000_10110001_0;
      patterns[14715] = 25'b00111001_01111001_10110010_0;
      patterns[14716] = 25'b00111001_01111010_10110011_0;
      patterns[14717] = 25'b00111001_01111011_10110100_0;
      patterns[14718] = 25'b00111001_01111100_10110101_0;
      patterns[14719] = 25'b00111001_01111101_10110110_0;
      patterns[14720] = 25'b00111001_01111110_10110111_0;
      patterns[14721] = 25'b00111001_01111111_10111000_0;
      patterns[14722] = 25'b00111001_10000000_10111001_0;
      patterns[14723] = 25'b00111001_10000001_10111010_0;
      patterns[14724] = 25'b00111001_10000010_10111011_0;
      patterns[14725] = 25'b00111001_10000011_10111100_0;
      patterns[14726] = 25'b00111001_10000100_10111101_0;
      patterns[14727] = 25'b00111001_10000101_10111110_0;
      patterns[14728] = 25'b00111001_10000110_10111111_0;
      patterns[14729] = 25'b00111001_10000111_11000000_0;
      patterns[14730] = 25'b00111001_10001000_11000001_0;
      patterns[14731] = 25'b00111001_10001001_11000010_0;
      patterns[14732] = 25'b00111001_10001010_11000011_0;
      patterns[14733] = 25'b00111001_10001011_11000100_0;
      patterns[14734] = 25'b00111001_10001100_11000101_0;
      patterns[14735] = 25'b00111001_10001101_11000110_0;
      patterns[14736] = 25'b00111001_10001110_11000111_0;
      patterns[14737] = 25'b00111001_10001111_11001000_0;
      patterns[14738] = 25'b00111001_10010000_11001001_0;
      patterns[14739] = 25'b00111001_10010001_11001010_0;
      patterns[14740] = 25'b00111001_10010010_11001011_0;
      patterns[14741] = 25'b00111001_10010011_11001100_0;
      patterns[14742] = 25'b00111001_10010100_11001101_0;
      patterns[14743] = 25'b00111001_10010101_11001110_0;
      patterns[14744] = 25'b00111001_10010110_11001111_0;
      patterns[14745] = 25'b00111001_10010111_11010000_0;
      patterns[14746] = 25'b00111001_10011000_11010001_0;
      patterns[14747] = 25'b00111001_10011001_11010010_0;
      patterns[14748] = 25'b00111001_10011010_11010011_0;
      patterns[14749] = 25'b00111001_10011011_11010100_0;
      patterns[14750] = 25'b00111001_10011100_11010101_0;
      patterns[14751] = 25'b00111001_10011101_11010110_0;
      patterns[14752] = 25'b00111001_10011110_11010111_0;
      patterns[14753] = 25'b00111001_10011111_11011000_0;
      patterns[14754] = 25'b00111001_10100000_11011001_0;
      patterns[14755] = 25'b00111001_10100001_11011010_0;
      patterns[14756] = 25'b00111001_10100010_11011011_0;
      patterns[14757] = 25'b00111001_10100011_11011100_0;
      patterns[14758] = 25'b00111001_10100100_11011101_0;
      patterns[14759] = 25'b00111001_10100101_11011110_0;
      patterns[14760] = 25'b00111001_10100110_11011111_0;
      patterns[14761] = 25'b00111001_10100111_11100000_0;
      patterns[14762] = 25'b00111001_10101000_11100001_0;
      patterns[14763] = 25'b00111001_10101001_11100010_0;
      patterns[14764] = 25'b00111001_10101010_11100011_0;
      patterns[14765] = 25'b00111001_10101011_11100100_0;
      patterns[14766] = 25'b00111001_10101100_11100101_0;
      patterns[14767] = 25'b00111001_10101101_11100110_0;
      patterns[14768] = 25'b00111001_10101110_11100111_0;
      patterns[14769] = 25'b00111001_10101111_11101000_0;
      patterns[14770] = 25'b00111001_10110000_11101001_0;
      patterns[14771] = 25'b00111001_10110001_11101010_0;
      patterns[14772] = 25'b00111001_10110010_11101011_0;
      patterns[14773] = 25'b00111001_10110011_11101100_0;
      patterns[14774] = 25'b00111001_10110100_11101101_0;
      patterns[14775] = 25'b00111001_10110101_11101110_0;
      patterns[14776] = 25'b00111001_10110110_11101111_0;
      patterns[14777] = 25'b00111001_10110111_11110000_0;
      patterns[14778] = 25'b00111001_10111000_11110001_0;
      patterns[14779] = 25'b00111001_10111001_11110010_0;
      patterns[14780] = 25'b00111001_10111010_11110011_0;
      patterns[14781] = 25'b00111001_10111011_11110100_0;
      patterns[14782] = 25'b00111001_10111100_11110101_0;
      patterns[14783] = 25'b00111001_10111101_11110110_0;
      patterns[14784] = 25'b00111001_10111110_11110111_0;
      patterns[14785] = 25'b00111001_10111111_11111000_0;
      patterns[14786] = 25'b00111001_11000000_11111001_0;
      patterns[14787] = 25'b00111001_11000001_11111010_0;
      patterns[14788] = 25'b00111001_11000010_11111011_0;
      patterns[14789] = 25'b00111001_11000011_11111100_0;
      patterns[14790] = 25'b00111001_11000100_11111101_0;
      patterns[14791] = 25'b00111001_11000101_11111110_0;
      patterns[14792] = 25'b00111001_11000110_11111111_0;
      patterns[14793] = 25'b00111001_11000111_00000000_1;
      patterns[14794] = 25'b00111001_11001000_00000001_1;
      patterns[14795] = 25'b00111001_11001001_00000010_1;
      patterns[14796] = 25'b00111001_11001010_00000011_1;
      patterns[14797] = 25'b00111001_11001011_00000100_1;
      patterns[14798] = 25'b00111001_11001100_00000101_1;
      patterns[14799] = 25'b00111001_11001101_00000110_1;
      patterns[14800] = 25'b00111001_11001110_00000111_1;
      patterns[14801] = 25'b00111001_11001111_00001000_1;
      patterns[14802] = 25'b00111001_11010000_00001001_1;
      patterns[14803] = 25'b00111001_11010001_00001010_1;
      patterns[14804] = 25'b00111001_11010010_00001011_1;
      patterns[14805] = 25'b00111001_11010011_00001100_1;
      patterns[14806] = 25'b00111001_11010100_00001101_1;
      patterns[14807] = 25'b00111001_11010101_00001110_1;
      patterns[14808] = 25'b00111001_11010110_00001111_1;
      patterns[14809] = 25'b00111001_11010111_00010000_1;
      patterns[14810] = 25'b00111001_11011000_00010001_1;
      patterns[14811] = 25'b00111001_11011001_00010010_1;
      patterns[14812] = 25'b00111001_11011010_00010011_1;
      patterns[14813] = 25'b00111001_11011011_00010100_1;
      patterns[14814] = 25'b00111001_11011100_00010101_1;
      patterns[14815] = 25'b00111001_11011101_00010110_1;
      patterns[14816] = 25'b00111001_11011110_00010111_1;
      patterns[14817] = 25'b00111001_11011111_00011000_1;
      patterns[14818] = 25'b00111001_11100000_00011001_1;
      patterns[14819] = 25'b00111001_11100001_00011010_1;
      patterns[14820] = 25'b00111001_11100010_00011011_1;
      patterns[14821] = 25'b00111001_11100011_00011100_1;
      patterns[14822] = 25'b00111001_11100100_00011101_1;
      patterns[14823] = 25'b00111001_11100101_00011110_1;
      patterns[14824] = 25'b00111001_11100110_00011111_1;
      patterns[14825] = 25'b00111001_11100111_00100000_1;
      patterns[14826] = 25'b00111001_11101000_00100001_1;
      patterns[14827] = 25'b00111001_11101001_00100010_1;
      patterns[14828] = 25'b00111001_11101010_00100011_1;
      patterns[14829] = 25'b00111001_11101011_00100100_1;
      patterns[14830] = 25'b00111001_11101100_00100101_1;
      patterns[14831] = 25'b00111001_11101101_00100110_1;
      patterns[14832] = 25'b00111001_11101110_00100111_1;
      patterns[14833] = 25'b00111001_11101111_00101000_1;
      patterns[14834] = 25'b00111001_11110000_00101001_1;
      patterns[14835] = 25'b00111001_11110001_00101010_1;
      patterns[14836] = 25'b00111001_11110010_00101011_1;
      patterns[14837] = 25'b00111001_11110011_00101100_1;
      patterns[14838] = 25'b00111001_11110100_00101101_1;
      patterns[14839] = 25'b00111001_11110101_00101110_1;
      patterns[14840] = 25'b00111001_11110110_00101111_1;
      patterns[14841] = 25'b00111001_11110111_00110000_1;
      patterns[14842] = 25'b00111001_11111000_00110001_1;
      patterns[14843] = 25'b00111001_11111001_00110010_1;
      patterns[14844] = 25'b00111001_11111010_00110011_1;
      patterns[14845] = 25'b00111001_11111011_00110100_1;
      patterns[14846] = 25'b00111001_11111100_00110101_1;
      patterns[14847] = 25'b00111001_11111101_00110110_1;
      patterns[14848] = 25'b00111001_11111110_00110111_1;
      patterns[14849] = 25'b00111001_11111111_00111000_1;
      patterns[14850] = 25'b00111010_00000000_00111010_0;
      patterns[14851] = 25'b00111010_00000001_00111011_0;
      patterns[14852] = 25'b00111010_00000010_00111100_0;
      patterns[14853] = 25'b00111010_00000011_00111101_0;
      patterns[14854] = 25'b00111010_00000100_00111110_0;
      patterns[14855] = 25'b00111010_00000101_00111111_0;
      patterns[14856] = 25'b00111010_00000110_01000000_0;
      patterns[14857] = 25'b00111010_00000111_01000001_0;
      patterns[14858] = 25'b00111010_00001000_01000010_0;
      patterns[14859] = 25'b00111010_00001001_01000011_0;
      patterns[14860] = 25'b00111010_00001010_01000100_0;
      patterns[14861] = 25'b00111010_00001011_01000101_0;
      patterns[14862] = 25'b00111010_00001100_01000110_0;
      patterns[14863] = 25'b00111010_00001101_01000111_0;
      patterns[14864] = 25'b00111010_00001110_01001000_0;
      patterns[14865] = 25'b00111010_00001111_01001001_0;
      patterns[14866] = 25'b00111010_00010000_01001010_0;
      patterns[14867] = 25'b00111010_00010001_01001011_0;
      patterns[14868] = 25'b00111010_00010010_01001100_0;
      patterns[14869] = 25'b00111010_00010011_01001101_0;
      patterns[14870] = 25'b00111010_00010100_01001110_0;
      patterns[14871] = 25'b00111010_00010101_01001111_0;
      patterns[14872] = 25'b00111010_00010110_01010000_0;
      patterns[14873] = 25'b00111010_00010111_01010001_0;
      patterns[14874] = 25'b00111010_00011000_01010010_0;
      patterns[14875] = 25'b00111010_00011001_01010011_0;
      patterns[14876] = 25'b00111010_00011010_01010100_0;
      patterns[14877] = 25'b00111010_00011011_01010101_0;
      patterns[14878] = 25'b00111010_00011100_01010110_0;
      patterns[14879] = 25'b00111010_00011101_01010111_0;
      patterns[14880] = 25'b00111010_00011110_01011000_0;
      patterns[14881] = 25'b00111010_00011111_01011001_0;
      patterns[14882] = 25'b00111010_00100000_01011010_0;
      patterns[14883] = 25'b00111010_00100001_01011011_0;
      patterns[14884] = 25'b00111010_00100010_01011100_0;
      patterns[14885] = 25'b00111010_00100011_01011101_0;
      patterns[14886] = 25'b00111010_00100100_01011110_0;
      patterns[14887] = 25'b00111010_00100101_01011111_0;
      patterns[14888] = 25'b00111010_00100110_01100000_0;
      patterns[14889] = 25'b00111010_00100111_01100001_0;
      patterns[14890] = 25'b00111010_00101000_01100010_0;
      patterns[14891] = 25'b00111010_00101001_01100011_0;
      patterns[14892] = 25'b00111010_00101010_01100100_0;
      patterns[14893] = 25'b00111010_00101011_01100101_0;
      patterns[14894] = 25'b00111010_00101100_01100110_0;
      patterns[14895] = 25'b00111010_00101101_01100111_0;
      patterns[14896] = 25'b00111010_00101110_01101000_0;
      patterns[14897] = 25'b00111010_00101111_01101001_0;
      patterns[14898] = 25'b00111010_00110000_01101010_0;
      patterns[14899] = 25'b00111010_00110001_01101011_0;
      patterns[14900] = 25'b00111010_00110010_01101100_0;
      patterns[14901] = 25'b00111010_00110011_01101101_0;
      patterns[14902] = 25'b00111010_00110100_01101110_0;
      patterns[14903] = 25'b00111010_00110101_01101111_0;
      patterns[14904] = 25'b00111010_00110110_01110000_0;
      patterns[14905] = 25'b00111010_00110111_01110001_0;
      patterns[14906] = 25'b00111010_00111000_01110010_0;
      patterns[14907] = 25'b00111010_00111001_01110011_0;
      patterns[14908] = 25'b00111010_00111010_01110100_0;
      patterns[14909] = 25'b00111010_00111011_01110101_0;
      patterns[14910] = 25'b00111010_00111100_01110110_0;
      patterns[14911] = 25'b00111010_00111101_01110111_0;
      patterns[14912] = 25'b00111010_00111110_01111000_0;
      patterns[14913] = 25'b00111010_00111111_01111001_0;
      patterns[14914] = 25'b00111010_01000000_01111010_0;
      patterns[14915] = 25'b00111010_01000001_01111011_0;
      patterns[14916] = 25'b00111010_01000010_01111100_0;
      patterns[14917] = 25'b00111010_01000011_01111101_0;
      patterns[14918] = 25'b00111010_01000100_01111110_0;
      patterns[14919] = 25'b00111010_01000101_01111111_0;
      patterns[14920] = 25'b00111010_01000110_10000000_0;
      patterns[14921] = 25'b00111010_01000111_10000001_0;
      patterns[14922] = 25'b00111010_01001000_10000010_0;
      patterns[14923] = 25'b00111010_01001001_10000011_0;
      patterns[14924] = 25'b00111010_01001010_10000100_0;
      patterns[14925] = 25'b00111010_01001011_10000101_0;
      patterns[14926] = 25'b00111010_01001100_10000110_0;
      patterns[14927] = 25'b00111010_01001101_10000111_0;
      patterns[14928] = 25'b00111010_01001110_10001000_0;
      patterns[14929] = 25'b00111010_01001111_10001001_0;
      patterns[14930] = 25'b00111010_01010000_10001010_0;
      patterns[14931] = 25'b00111010_01010001_10001011_0;
      patterns[14932] = 25'b00111010_01010010_10001100_0;
      patterns[14933] = 25'b00111010_01010011_10001101_0;
      patterns[14934] = 25'b00111010_01010100_10001110_0;
      patterns[14935] = 25'b00111010_01010101_10001111_0;
      patterns[14936] = 25'b00111010_01010110_10010000_0;
      patterns[14937] = 25'b00111010_01010111_10010001_0;
      patterns[14938] = 25'b00111010_01011000_10010010_0;
      patterns[14939] = 25'b00111010_01011001_10010011_0;
      patterns[14940] = 25'b00111010_01011010_10010100_0;
      patterns[14941] = 25'b00111010_01011011_10010101_0;
      patterns[14942] = 25'b00111010_01011100_10010110_0;
      patterns[14943] = 25'b00111010_01011101_10010111_0;
      patterns[14944] = 25'b00111010_01011110_10011000_0;
      patterns[14945] = 25'b00111010_01011111_10011001_0;
      patterns[14946] = 25'b00111010_01100000_10011010_0;
      patterns[14947] = 25'b00111010_01100001_10011011_0;
      patterns[14948] = 25'b00111010_01100010_10011100_0;
      patterns[14949] = 25'b00111010_01100011_10011101_0;
      patterns[14950] = 25'b00111010_01100100_10011110_0;
      patterns[14951] = 25'b00111010_01100101_10011111_0;
      patterns[14952] = 25'b00111010_01100110_10100000_0;
      patterns[14953] = 25'b00111010_01100111_10100001_0;
      patterns[14954] = 25'b00111010_01101000_10100010_0;
      patterns[14955] = 25'b00111010_01101001_10100011_0;
      patterns[14956] = 25'b00111010_01101010_10100100_0;
      patterns[14957] = 25'b00111010_01101011_10100101_0;
      patterns[14958] = 25'b00111010_01101100_10100110_0;
      patterns[14959] = 25'b00111010_01101101_10100111_0;
      patterns[14960] = 25'b00111010_01101110_10101000_0;
      patterns[14961] = 25'b00111010_01101111_10101001_0;
      patterns[14962] = 25'b00111010_01110000_10101010_0;
      patterns[14963] = 25'b00111010_01110001_10101011_0;
      patterns[14964] = 25'b00111010_01110010_10101100_0;
      patterns[14965] = 25'b00111010_01110011_10101101_0;
      patterns[14966] = 25'b00111010_01110100_10101110_0;
      patterns[14967] = 25'b00111010_01110101_10101111_0;
      patterns[14968] = 25'b00111010_01110110_10110000_0;
      patterns[14969] = 25'b00111010_01110111_10110001_0;
      patterns[14970] = 25'b00111010_01111000_10110010_0;
      patterns[14971] = 25'b00111010_01111001_10110011_0;
      patterns[14972] = 25'b00111010_01111010_10110100_0;
      patterns[14973] = 25'b00111010_01111011_10110101_0;
      patterns[14974] = 25'b00111010_01111100_10110110_0;
      patterns[14975] = 25'b00111010_01111101_10110111_0;
      patterns[14976] = 25'b00111010_01111110_10111000_0;
      patterns[14977] = 25'b00111010_01111111_10111001_0;
      patterns[14978] = 25'b00111010_10000000_10111010_0;
      patterns[14979] = 25'b00111010_10000001_10111011_0;
      patterns[14980] = 25'b00111010_10000010_10111100_0;
      patterns[14981] = 25'b00111010_10000011_10111101_0;
      patterns[14982] = 25'b00111010_10000100_10111110_0;
      patterns[14983] = 25'b00111010_10000101_10111111_0;
      patterns[14984] = 25'b00111010_10000110_11000000_0;
      patterns[14985] = 25'b00111010_10000111_11000001_0;
      patterns[14986] = 25'b00111010_10001000_11000010_0;
      patterns[14987] = 25'b00111010_10001001_11000011_0;
      patterns[14988] = 25'b00111010_10001010_11000100_0;
      patterns[14989] = 25'b00111010_10001011_11000101_0;
      patterns[14990] = 25'b00111010_10001100_11000110_0;
      patterns[14991] = 25'b00111010_10001101_11000111_0;
      patterns[14992] = 25'b00111010_10001110_11001000_0;
      patterns[14993] = 25'b00111010_10001111_11001001_0;
      patterns[14994] = 25'b00111010_10010000_11001010_0;
      patterns[14995] = 25'b00111010_10010001_11001011_0;
      patterns[14996] = 25'b00111010_10010010_11001100_0;
      patterns[14997] = 25'b00111010_10010011_11001101_0;
      patterns[14998] = 25'b00111010_10010100_11001110_0;
      patterns[14999] = 25'b00111010_10010101_11001111_0;
      patterns[15000] = 25'b00111010_10010110_11010000_0;
      patterns[15001] = 25'b00111010_10010111_11010001_0;
      patterns[15002] = 25'b00111010_10011000_11010010_0;
      patterns[15003] = 25'b00111010_10011001_11010011_0;
      patterns[15004] = 25'b00111010_10011010_11010100_0;
      patterns[15005] = 25'b00111010_10011011_11010101_0;
      patterns[15006] = 25'b00111010_10011100_11010110_0;
      patterns[15007] = 25'b00111010_10011101_11010111_0;
      patterns[15008] = 25'b00111010_10011110_11011000_0;
      patterns[15009] = 25'b00111010_10011111_11011001_0;
      patterns[15010] = 25'b00111010_10100000_11011010_0;
      patterns[15011] = 25'b00111010_10100001_11011011_0;
      patterns[15012] = 25'b00111010_10100010_11011100_0;
      patterns[15013] = 25'b00111010_10100011_11011101_0;
      patterns[15014] = 25'b00111010_10100100_11011110_0;
      patterns[15015] = 25'b00111010_10100101_11011111_0;
      patterns[15016] = 25'b00111010_10100110_11100000_0;
      patterns[15017] = 25'b00111010_10100111_11100001_0;
      patterns[15018] = 25'b00111010_10101000_11100010_0;
      patterns[15019] = 25'b00111010_10101001_11100011_0;
      patterns[15020] = 25'b00111010_10101010_11100100_0;
      patterns[15021] = 25'b00111010_10101011_11100101_0;
      patterns[15022] = 25'b00111010_10101100_11100110_0;
      patterns[15023] = 25'b00111010_10101101_11100111_0;
      patterns[15024] = 25'b00111010_10101110_11101000_0;
      patterns[15025] = 25'b00111010_10101111_11101001_0;
      patterns[15026] = 25'b00111010_10110000_11101010_0;
      patterns[15027] = 25'b00111010_10110001_11101011_0;
      patterns[15028] = 25'b00111010_10110010_11101100_0;
      patterns[15029] = 25'b00111010_10110011_11101101_0;
      patterns[15030] = 25'b00111010_10110100_11101110_0;
      patterns[15031] = 25'b00111010_10110101_11101111_0;
      patterns[15032] = 25'b00111010_10110110_11110000_0;
      patterns[15033] = 25'b00111010_10110111_11110001_0;
      patterns[15034] = 25'b00111010_10111000_11110010_0;
      patterns[15035] = 25'b00111010_10111001_11110011_0;
      patterns[15036] = 25'b00111010_10111010_11110100_0;
      patterns[15037] = 25'b00111010_10111011_11110101_0;
      patterns[15038] = 25'b00111010_10111100_11110110_0;
      patterns[15039] = 25'b00111010_10111101_11110111_0;
      patterns[15040] = 25'b00111010_10111110_11111000_0;
      patterns[15041] = 25'b00111010_10111111_11111001_0;
      patterns[15042] = 25'b00111010_11000000_11111010_0;
      patterns[15043] = 25'b00111010_11000001_11111011_0;
      patterns[15044] = 25'b00111010_11000010_11111100_0;
      patterns[15045] = 25'b00111010_11000011_11111101_0;
      patterns[15046] = 25'b00111010_11000100_11111110_0;
      patterns[15047] = 25'b00111010_11000101_11111111_0;
      patterns[15048] = 25'b00111010_11000110_00000000_1;
      patterns[15049] = 25'b00111010_11000111_00000001_1;
      patterns[15050] = 25'b00111010_11001000_00000010_1;
      patterns[15051] = 25'b00111010_11001001_00000011_1;
      patterns[15052] = 25'b00111010_11001010_00000100_1;
      patterns[15053] = 25'b00111010_11001011_00000101_1;
      patterns[15054] = 25'b00111010_11001100_00000110_1;
      patterns[15055] = 25'b00111010_11001101_00000111_1;
      patterns[15056] = 25'b00111010_11001110_00001000_1;
      patterns[15057] = 25'b00111010_11001111_00001001_1;
      patterns[15058] = 25'b00111010_11010000_00001010_1;
      patterns[15059] = 25'b00111010_11010001_00001011_1;
      patterns[15060] = 25'b00111010_11010010_00001100_1;
      patterns[15061] = 25'b00111010_11010011_00001101_1;
      patterns[15062] = 25'b00111010_11010100_00001110_1;
      patterns[15063] = 25'b00111010_11010101_00001111_1;
      patterns[15064] = 25'b00111010_11010110_00010000_1;
      patterns[15065] = 25'b00111010_11010111_00010001_1;
      patterns[15066] = 25'b00111010_11011000_00010010_1;
      patterns[15067] = 25'b00111010_11011001_00010011_1;
      patterns[15068] = 25'b00111010_11011010_00010100_1;
      patterns[15069] = 25'b00111010_11011011_00010101_1;
      patterns[15070] = 25'b00111010_11011100_00010110_1;
      patterns[15071] = 25'b00111010_11011101_00010111_1;
      patterns[15072] = 25'b00111010_11011110_00011000_1;
      patterns[15073] = 25'b00111010_11011111_00011001_1;
      patterns[15074] = 25'b00111010_11100000_00011010_1;
      patterns[15075] = 25'b00111010_11100001_00011011_1;
      patterns[15076] = 25'b00111010_11100010_00011100_1;
      patterns[15077] = 25'b00111010_11100011_00011101_1;
      patterns[15078] = 25'b00111010_11100100_00011110_1;
      patterns[15079] = 25'b00111010_11100101_00011111_1;
      patterns[15080] = 25'b00111010_11100110_00100000_1;
      patterns[15081] = 25'b00111010_11100111_00100001_1;
      patterns[15082] = 25'b00111010_11101000_00100010_1;
      patterns[15083] = 25'b00111010_11101001_00100011_1;
      patterns[15084] = 25'b00111010_11101010_00100100_1;
      patterns[15085] = 25'b00111010_11101011_00100101_1;
      patterns[15086] = 25'b00111010_11101100_00100110_1;
      patterns[15087] = 25'b00111010_11101101_00100111_1;
      patterns[15088] = 25'b00111010_11101110_00101000_1;
      patterns[15089] = 25'b00111010_11101111_00101001_1;
      patterns[15090] = 25'b00111010_11110000_00101010_1;
      patterns[15091] = 25'b00111010_11110001_00101011_1;
      patterns[15092] = 25'b00111010_11110010_00101100_1;
      patterns[15093] = 25'b00111010_11110011_00101101_1;
      patterns[15094] = 25'b00111010_11110100_00101110_1;
      patterns[15095] = 25'b00111010_11110101_00101111_1;
      patterns[15096] = 25'b00111010_11110110_00110000_1;
      patterns[15097] = 25'b00111010_11110111_00110001_1;
      patterns[15098] = 25'b00111010_11111000_00110010_1;
      patterns[15099] = 25'b00111010_11111001_00110011_1;
      patterns[15100] = 25'b00111010_11111010_00110100_1;
      patterns[15101] = 25'b00111010_11111011_00110101_1;
      patterns[15102] = 25'b00111010_11111100_00110110_1;
      patterns[15103] = 25'b00111010_11111101_00110111_1;
      patterns[15104] = 25'b00111010_11111110_00111000_1;
      patterns[15105] = 25'b00111010_11111111_00111001_1;
      patterns[15106] = 25'b00111011_00000000_00111011_0;
      patterns[15107] = 25'b00111011_00000001_00111100_0;
      patterns[15108] = 25'b00111011_00000010_00111101_0;
      patterns[15109] = 25'b00111011_00000011_00111110_0;
      patterns[15110] = 25'b00111011_00000100_00111111_0;
      patterns[15111] = 25'b00111011_00000101_01000000_0;
      patterns[15112] = 25'b00111011_00000110_01000001_0;
      patterns[15113] = 25'b00111011_00000111_01000010_0;
      patterns[15114] = 25'b00111011_00001000_01000011_0;
      patterns[15115] = 25'b00111011_00001001_01000100_0;
      patterns[15116] = 25'b00111011_00001010_01000101_0;
      patterns[15117] = 25'b00111011_00001011_01000110_0;
      patterns[15118] = 25'b00111011_00001100_01000111_0;
      patterns[15119] = 25'b00111011_00001101_01001000_0;
      patterns[15120] = 25'b00111011_00001110_01001001_0;
      patterns[15121] = 25'b00111011_00001111_01001010_0;
      patterns[15122] = 25'b00111011_00010000_01001011_0;
      patterns[15123] = 25'b00111011_00010001_01001100_0;
      patterns[15124] = 25'b00111011_00010010_01001101_0;
      patterns[15125] = 25'b00111011_00010011_01001110_0;
      patterns[15126] = 25'b00111011_00010100_01001111_0;
      patterns[15127] = 25'b00111011_00010101_01010000_0;
      patterns[15128] = 25'b00111011_00010110_01010001_0;
      patterns[15129] = 25'b00111011_00010111_01010010_0;
      patterns[15130] = 25'b00111011_00011000_01010011_0;
      patterns[15131] = 25'b00111011_00011001_01010100_0;
      patterns[15132] = 25'b00111011_00011010_01010101_0;
      patterns[15133] = 25'b00111011_00011011_01010110_0;
      patterns[15134] = 25'b00111011_00011100_01010111_0;
      patterns[15135] = 25'b00111011_00011101_01011000_0;
      patterns[15136] = 25'b00111011_00011110_01011001_0;
      patterns[15137] = 25'b00111011_00011111_01011010_0;
      patterns[15138] = 25'b00111011_00100000_01011011_0;
      patterns[15139] = 25'b00111011_00100001_01011100_0;
      patterns[15140] = 25'b00111011_00100010_01011101_0;
      patterns[15141] = 25'b00111011_00100011_01011110_0;
      patterns[15142] = 25'b00111011_00100100_01011111_0;
      patterns[15143] = 25'b00111011_00100101_01100000_0;
      patterns[15144] = 25'b00111011_00100110_01100001_0;
      patterns[15145] = 25'b00111011_00100111_01100010_0;
      patterns[15146] = 25'b00111011_00101000_01100011_0;
      patterns[15147] = 25'b00111011_00101001_01100100_0;
      patterns[15148] = 25'b00111011_00101010_01100101_0;
      patterns[15149] = 25'b00111011_00101011_01100110_0;
      patterns[15150] = 25'b00111011_00101100_01100111_0;
      patterns[15151] = 25'b00111011_00101101_01101000_0;
      patterns[15152] = 25'b00111011_00101110_01101001_0;
      patterns[15153] = 25'b00111011_00101111_01101010_0;
      patterns[15154] = 25'b00111011_00110000_01101011_0;
      patterns[15155] = 25'b00111011_00110001_01101100_0;
      patterns[15156] = 25'b00111011_00110010_01101101_0;
      patterns[15157] = 25'b00111011_00110011_01101110_0;
      patterns[15158] = 25'b00111011_00110100_01101111_0;
      patterns[15159] = 25'b00111011_00110101_01110000_0;
      patterns[15160] = 25'b00111011_00110110_01110001_0;
      patterns[15161] = 25'b00111011_00110111_01110010_0;
      patterns[15162] = 25'b00111011_00111000_01110011_0;
      patterns[15163] = 25'b00111011_00111001_01110100_0;
      patterns[15164] = 25'b00111011_00111010_01110101_0;
      patterns[15165] = 25'b00111011_00111011_01110110_0;
      patterns[15166] = 25'b00111011_00111100_01110111_0;
      patterns[15167] = 25'b00111011_00111101_01111000_0;
      patterns[15168] = 25'b00111011_00111110_01111001_0;
      patterns[15169] = 25'b00111011_00111111_01111010_0;
      patterns[15170] = 25'b00111011_01000000_01111011_0;
      patterns[15171] = 25'b00111011_01000001_01111100_0;
      patterns[15172] = 25'b00111011_01000010_01111101_0;
      patterns[15173] = 25'b00111011_01000011_01111110_0;
      patterns[15174] = 25'b00111011_01000100_01111111_0;
      patterns[15175] = 25'b00111011_01000101_10000000_0;
      patterns[15176] = 25'b00111011_01000110_10000001_0;
      patterns[15177] = 25'b00111011_01000111_10000010_0;
      patterns[15178] = 25'b00111011_01001000_10000011_0;
      patterns[15179] = 25'b00111011_01001001_10000100_0;
      patterns[15180] = 25'b00111011_01001010_10000101_0;
      patterns[15181] = 25'b00111011_01001011_10000110_0;
      patterns[15182] = 25'b00111011_01001100_10000111_0;
      patterns[15183] = 25'b00111011_01001101_10001000_0;
      patterns[15184] = 25'b00111011_01001110_10001001_0;
      patterns[15185] = 25'b00111011_01001111_10001010_0;
      patterns[15186] = 25'b00111011_01010000_10001011_0;
      patterns[15187] = 25'b00111011_01010001_10001100_0;
      patterns[15188] = 25'b00111011_01010010_10001101_0;
      patterns[15189] = 25'b00111011_01010011_10001110_0;
      patterns[15190] = 25'b00111011_01010100_10001111_0;
      patterns[15191] = 25'b00111011_01010101_10010000_0;
      patterns[15192] = 25'b00111011_01010110_10010001_0;
      patterns[15193] = 25'b00111011_01010111_10010010_0;
      patterns[15194] = 25'b00111011_01011000_10010011_0;
      patterns[15195] = 25'b00111011_01011001_10010100_0;
      patterns[15196] = 25'b00111011_01011010_10010101_0;
      patterns[15197] = 25'b00111011_01011011_10010110_0;
      patterns[15198] = 25'b00111011_01011100_10010111_0;
      patterns[15199] = 25'b00111011_01011101_10011000_0;
      patterns[15200] = 25'b00111011_01011110_10011001_0;
      patterns[15201] = 25'b00111011_01011111_10011010_0;
      patterns[15202] = 25'b00111011_01100000_10011011_0;
      patterns[15203] = 25'b00111011_01100001_10011100_0;
      patterns[15204] = 25'b00111011_01100010_10011101_0;
      patterns[15205] = 25'b00111011_01100011_10011110_0;
      patterns[15206] = 25'b00111011_01100100_10011111_0;
      patterns[15207] = 25'b00111011_01100101_10100000_0;
      patterns[15208] = 25'b00111011_01100110_10100001_0;
      patterns[15209] = 25'b00111011_01100111_10100010_0;
      patterns[15210] = 25'b00111011_01101000_10100011_0;
      patterns[15211] = 25'b00111011_01101001_10100100_0;
      patterns[15212] = 25'b00111011_01101010_10100101_0;
      patterns[15213] = 25'b00111011_01101011_10100110_0;
      patterns[15214] = 25'b00111011_01101100_10100111_0;
      patterns[15215] = 25'b00111011_01101101_10101000_0;
      patterns[15216] = 25'b00111011_01101110_10101001_0;
      patterns[15217] = 25'b00111011_01101111_10101010_0;
      patterns[15218] = 25'b00111011_01110000_10101011_0;
      patterns[15219] = 25'b00111011_01110001_10101100_0;
      patterns[15220] = 25'b00111011_01110010_10101101_0;
      patterns[15221] = 25'b00111011_01110011_10101110_0;
      patterns[15222] = 25'b00111011_01110100_10101111_0;
      patterns[15223] = 25'b00111011_01110101_10110000_0;
      patterns[15224] = 25'b00111011_01110110_10110001_0;
      patterns[15225] = 25'b00111011_01110111_10110010_0;
      patterns[15226] = 25'b00111011_01111000_10110011_0;
      patterns[15227] = 25'b00111011_01111001_10110100_0;
      patterns[15228] = 25'b00111011_01111010_10110101_0;
      patterns[15229] = 25'b00111011_01111011_10110110_0;
      patterns[15230] = 25'b00111011_01111100_10110111_0;
      patterns[15231] = 25'b00111011_01111101_10111000_0;
      patterns[15232] = 25'b00111011_01111110_10111001_0;
      patterns[15233] = 25'b00111011_01111111_10111010_0;
      patterns[15234] = 25'b00111011_10000000_10111011_0;
      patterns[15235] = 25'b00111011_10000001_10111100_0;
      patterns[15236] = 25'b00111011_10000010_10111101_0;
      patterns[15237] = 25'b00111011_10000011_10111110_0;
      patterns[15238] = 25'b00111011_10000100_10111111_0;
      patterns[15239] = 25'b00111011_10000101_11000000_0;
      patterns[15240] = 25'b00111011_10000110_11000001_0;
      patterns[15241] = 25'b00111011_10000111_11000010_0;
      patterns[15242] = 25'b00111011_10001000_11000011_0;
      patterns[15243] = 25'b00111011_10001001_11000100_0;
      patterns[15244] = 25'b00111011_10001010_11000101_0;
      patterns[15245] = 25'b00111011_10001011_11000110_0;
      patterns[15246] = 25'b00111011_10001100_11000111_0;
      patterns[15247] = 25'b00111011_10001101_11001000_0;
      patterns[15248] = 25'b00111011_10001110_11001001_0;
      patterns[15249] = 25'b00111011_10001111_11001010_0;
      patterns[15250] = 25'b00111011_10010000_11001011_0;
      patterns[15251] = 25'b00111011_10010001_11001100_0;
      patterns[15252] = 25'b00111011_10010010_11001101_0;
      patterns[15253] = 25'b00111011_10010011_11001110_0;
      patterns[15254] = 25'b00111011_10010100_11001111_0;
      patterns[15255] = 25'b00111011_10010101_11010000_0;
      patterns[15256] = 25'b00111011_10010110_11010001_0;
      patterns[15257] = 25'b00111011_10010111_11010010_0;
      patterns[15258] = 25'b00111011_10011000_11010011_0;
      patterns[15259] = 25'b00111011_10011001_11010100_0;
      patterns[15260] = 25'b00111011_10011010_11010101_0;
      patterns[15261] = 25'b00111011_10011011_11010110_0;
      patterns[15262] = 25'b00111011_10011100_11010111_0;
      patterns[15263] = 25'b00111011_10011101_11011000_0;
      patterns[15264] = 25'b00111011_10011110_11011001_0;
      patterns[15265] = 25'b00111011_10011111_11011010_0;
      patterns[15266] = 25'b00111011_10100000_11011011_0;
      patterns[15267] = 25'b00111011_10100001_11011100_0;
      patterns[15268] = 25'b00111011_10100010_11011101_0;
      patterns[15269] = 25'b00111011_10100011_11011110_0;
      patterns[15270] = 25'b00111011_10100100_11011111_0;
      patterns[15271] = 25'b00111011_10100101_11100000_0;
      patterns[15272] = 25'b00111011_10100110_11100001_0;
      patterns[15273] = 25'b00111011_10100111_11100010_0;
      patterns[15274] = 25'b00111011_10101000_11100011_0;
      patterns[15275] = 25'b00111011_10101001_11100100_0;
      patterns[15276] = 25'b00111011_10101010_11100101_0;
      patterns[15277] = 25'b00111011_10101011_11100110_0;
      patterns[15278] = 25'b00111011_10101100_11100111_0;
      patterns[15279] = 25'b00111011_10101101_11101000_0;
      patterns[15280] = 25'b00111011_10101110_11101001_0;
      patterns[15281] = 25'b00111011_10101111_11101010_0;
      patterns[15282] = 25'b00111011_10110000_11101011_0;
      patterns[15283] = 25'b00111011_10110001_11101100_0;
      patterns[15284] = 25'b00111011_10110010_11101101_0;
      patterns[15285] = 25'b00111011_10110011_11101110_0;
      patterns[15286] = 25'b00111011_10110100_11101111_0;
      patterns[15287] = 25'b00111011_10110101_11110000_0;
      patterns[15288] = 25'b00111011_10110110_11110001_0;
      patterns[15289] = 25'b00111011_10110111_11110010_0;
      patterns[15290] = 25'b00111011_10111000_11110011_0;
      patterns[15291] = 25'b00111011_10111001_11110100_0;
      patterns[15292] = 25'b00111011_10111010_11110101_0;
      patterns[15293] = 25'b00111011_10111011_11110110_0;
      patterns[15294] = 25'b00111011_10111100_11110111_0;
      patterns[15295] = 25'b00111011_10111101_11111000_0;
      patterns[15296] = 25'b00111011_10111110_11111001_0;
      patterns[15297] = 25'b00111011_10111111_11111010_0;
      patterns[15298] = 25'b00111011_11000000_11111011_0;
      patterns[15299] = 25'b00111011_11000001_11111100_0;
      patterns[15300] = 25'b00111011_11000010_11111101_0;
      patterns[15301] = 25'b00111011_11000011_11111110_0;
      patterns[15302] = 25'b00111011_11000100_11111111_0;
      patterns[15303] = 25'b00111011_11000101_00000000_1;
      patterns[15304] = 25'b00111011_11000110_00000001_1;
      patterns[15305] = 25'b00111011_11000111_00000010_1;
      patterns[15306] = 25'b00111011_11001000_00000011_1;
      patterns[15307] = 25'b00111011_11001001_00000100_1;
      patterns[15308] = 25'b00111011_11001010_00000101_1;
      patterns[15309] = 25'b00111011_11001011_00000110_1;
      patterns[15310] = 25'b00111011_11001100_00000111_1;
      patterns[15311] = 25'b00111011_11001101_00001000_1;
      patterns[15312] = 25'b00111011_11001110_00001001_1;
      patterns[15313] = 25'b00111011_11001111_00001010_1;
      patterns[15314] = 25'b00111011_11010000_00001011_1;
      patterns[15315] = 25'b00111011_11010001_00001100_1;
      patterns[15316] = 25'b00111011_11010010_00001101_1;
      patterns[15317] = 25'b00111011_11010011_00001110_1;
      patterns[15318] = 25'b00111011_11010100_00001111_1;
      patterns[15319] = 25'b00111011_11010101_00010000_1;
      patterns[15320] = 25'b00111011_11010110_00010001_1;
      patterns[15321] = 25'b00111011_11010111_00010010_1;
      patterns[15322] = 25'b00111011_11011000_00010011_1;
      patterns[15323] = 25'b00111011_11011001_00010100_1;
      patterns[15324] = 25'b00111011_11011010_00010101_1;
      patterns[15325] = 25'b00111011_11011011_00010110_1;
      patterns[15326] = 25'b00111011_11011100_00010111_1;
      patterns[15327] = 25'b00111011_11011101_00011000_1;
      patterns[15328] = 25'b00111011_11011110_00011001_1;
      patterns[15329] = 25'b00111011_11011111_00011010_1;
      patterns[15330] = 25'b00111011_11100000_00011011_1;
      patterns[15331] = 25'b00111011_11100001_00011100_1;
      patterns[15332] = 25'b00111011_11100010_00011101_1;
      patterns[15333] = 25'b00111011_11100011_00011110_1;
      patterns[15334] = 25'b00111011_11100100_00011111_1;
      patterns[15335] = 25'b00111011_11100101_00100000_1;
      patterns[15336] = 25'b00111011_11100110_00100001_1;
      patterns[15337] = 25'b00111011_11100111_00100010_1;
      patterns[15338] = 25'b00111011_11101000_00100011_1;
      patterns[15339] = 25'b00111011_11101001_00100100_1;
      patterns[15340] = 25'b00111011_11101010_00100101_1;
      patterns[15341] = 25'b00111011_11101011_00100110_1;
      patterns[15342] = 25'b00111011_11101100_00100111_1;
      patterns[15343] = 25'b00111011_11101101_00101000_1;
      patterns[15344] = 25'b00111011_11101110_00101001_1;
      patterns[15345] = 25'b00111011_11101111_00101010_1;
      patterns[15346] = 25'b00111011_11110000_00101011_1;
      patterns[15347] = 25'b00111011_11110001_00101100_1;
      patterns[15348] = 25'b00111011_11110010_00101101_1;
      patterns[15349] = 25'b00111011_11110011_00101110_1;
      patterns[15350] = 25'b00111011_11110100_00101111_1;
      patterns[15351] = 25'b00111011_11110101_00110000_1;
      patterns[15352] = 25'b00111011_11110110_00110001_1;
      patterns[15353] = 25'b00111011_11110111_00110010_1;
      patterns[15354] = 25'b00111011_11111000_00110011_1;
      patterns[15355] = 25'b00111011_11111001_00110100_1;
      patterns[15356] = 25'b00111011_11111010_00110101_1;
      patterns[15357] = 25'b00111011_11111011_00110110_1;
      patterns[15358] = 25'b00111011_11111100_00110111_1;
      patterns[15359] = 25'b00111011_11111101_00111000_1;
      patterns[15360] = 25'b00111011_11111110_00111001_1;
      patterns[15361] = 25'b00111011_11111111_00111010_1;
      patterns[15362] = 25'b00111100_00000000_00111100_0;
      patterns[15363] = 25'b00111100_00000001_00111101_0;
      patterns[15364] = 25'b00111100_00000010_00111110_0;
      patterns[15365] = 25'b00111100_00000011_00111111_0;
      patterns[15366] = 25'b00111100_00000100_01000000_0;
      patterns[15367] = 25'b00111100_00000101_01000001_0;
      patterns[15368] = 25'b00111100_00000110_01000010_0;
      patterns[15369] = 25'b00111100_00000111_01000011_0;
      patterns[15370] = 25'b00111100_00001000_01000100_0;
      patterns[15371] = 25'b00111100_00001001_01000101_0;
      patterns[15372] = 25'b00111100_00001010_01000110_0;
      patterns[15373] = 25'b00111100_00001011_01000111_0;
      patterns[15374] = 25'b00111100_00001100_01001000_0;
      patterns[15375] = 25'b00111100_00001101_01001001_0;
      patterns[15376] = 25'b00111100_00001110_01001010_0;
      patterns[15377] = 25'b00111100_00001111_01001011_0;
      patterns[15378] = 25'b00111100_00010000_01001100_0;
      patterns[15379] = 25'b00111100_00010001_01001101_0;
      patterns[15380] = 25'b00111100_00010010_01001110_0;
      patterns[15381] = 25'b00111100_00010011_01001111_0;
      patterns[15382] = 25'b00111100_00010100_01010000_0;
      patterns[15383] = 25'b00111100_00010101_01010001_0;
      patterns[15384] = 25'b00111100_00010110_01010010_0;
      patterns[15385] = 25'b00111100_00010111_01010011_0;
      patterns[15386] = 25'b00111100_00011000_01010100_0;
      patterns[15387] = 25'b00111100_00011001_01010101_0;
      patterns[15388] = 25'b00111100_00011010_01010110_0;
      patterns[15389] = 25'b00111100_00011011_01010111_0;
      patterns[15390] = 25'b00111100_00011100_01011000_0;
      patterns[15391] = 25'b00111100_00011101_01011001_0;
      patterns[15392] = 25'b00111100_00011110_01011010_0;
      patterns[15393] = 25'b00111100_00011111_01011011_0;
      patterns[15394] = 25'b00111100_00100000_01011100_0;
      patterns[15395] = 25'b00111100_00100001_01011101_0;
      patterns[15396] = 25'b00111100_00100010_01011110_0;
      patterns[15397] = 25'b00111100_00100011_01011111_0;
      patterns[15398] = 25'b00111100_00100100_01100000_0;
      patterns[15399] = 25'b00111100_00100101_01100001_0;
      patterns[15400] = 25'b00111100_00100110_01100010_0;
      patterns[15401] = 25'b00111100_00100111_01100011_0;
      patterns[15402] = 25'b00111100_00101000_01100100_0;
      patterns[15403] = 25'b00111100_00101001_01100101_0;
      patterns[15404] = 25'b00111100_00101010_01100110_0;
      patterns[15405] = 25'b00111100_00101011_01100111_0;
      patterns[15406] = 25'b00111100_00101100_01101000_0;
      patterns[15407] = 25'b00111100_00101101_01101001_0;
      patterns[15408] = 25'b00111100_00101110_01101010_0;
      patterns[15409] = 25'b00111100_00101111_01101011_0;
      patterns[15410] = 25'b00111100_00110000_01101100_0;
      patterns[15411] = 25'b00111100_00110001_01101101_0;
      patterns[15412] = 25'b00111100_00110010_01101110_0;
      patterns[15413] = 25'b00111100_00110011_01101111_0;
      patterns[15414] = 25'b00111100_00110100_01110000_0;
      patterns[15415] = 25'b00111100_00110101_01110001_0;
      patterns[15416] = 25'b00111100_00110110_01110010_0;
      patterns[15417] = 25'b00111100_00110111_01110011_0;
      patterns[15418] = 25'b00111100_00111000_01110100_0;
      patterns[15419] = 25'b00111100_00111001_01110101_0;
      patterns[15420] = 25'b00111100_00111010_01110110_0;
      patterns[15421] = 25'b00111100_00111011_01110111_0;
      patterns[15422] = 25'b00111100_00111100_01111000_0;
      patterns[15423] = 25'b00111100_00111101_01111001_0;
      patterns[15424] = 25'b00111100_00111110_01111010_0;
      patterns[15425] = 25'b00111100_00111111_01111011_0;
      patterns[15426] = 25'b00111100_01000000_01111100_0;
      patterns[15427] = 25'b00111100_01000001_01111101_0;
      patterns[15428] = 25'b00111100_01000010_01111110_0;
      patterns[15429] = 25'b00111100_01000011_01111111_0;
      patterns[15430] = 25'b00111100_01000100_10000000_0;
      patterns[15431] = 25'b00111100_01000101_10000001_0;
      patterns[15432] = 25'b00111100_01000110_10000010_0;
      patterns[15433] = 25'b00111100_01000111_10000011_0;
      patterns[15434] = 25'b00111100_01001000_10000100_0;
      patterns[15435] = 25'b00111100_01001001_10000101_0;
      patterns[15436] = 25'b00111100_01001010_10000110_0;
      patterns[15437] = 25'b00111100_01001011_10000111_0;
      patterns[15438] = 25'b00111100_01001100_10001000_0;
      patterns[15439] = 25'b00111100_01001101_10001001_0;
      patterns[15440] = 25'b00111100_01001110_10001010_0;
      patterns[15441] = 25'b00111100_01001111_10001011_0;
      patterns[15442] = 25'b00111100_01010000_10001100_0;
      patterns[15443] = 25'b00111100_01010001_10001101_0;
      patterns[15444] = 25'b00111100_01010010_10001110_0;
      patterns[15445] = 25'b00111100_01010011_10001111_0;
      patterns[15446] = 25'b00111100_01010100_10010000_0;
      patterns[15447] = 25'b00111100_01010101_10010001_0;
      patterns[15448] = 25'b00111100_01010110_10010010_0;
      patterns[15449] = 25'b00111100_01010111_10010011_0;
      patterns[15450] = 25'b00111100_01011000_10010100_0;
      patterns[15451] = 25'b00111100_01011001_10010101_0;
      patterns[15452] = 25'b00111100_01011010_10010110_0;
      patterns[15453] = 25'b00111100_01011011_10010111_0;
      patterns[15454] = 25'b00111100_01011100_10011000_0;
      patterns[15455] = 25'b00111100_01011101_10011001_0;
      patterns[15456] = 25'b00111100_01011110_10011010_0;
      patterns[15457] = 25'b00111100_01011111_10011011_0;
      patterns[15458] = 25'b00111100_01100000_10011100_0;
      patterns[15459] = 25'b00111100_01100001_10011101_0;
      patterns[15460] = 25'b00111100_01100010_10011110_0;
      patterns[15461] = 25'b00111100_01100011_10011111_0;
      patterns[15462] = 25'b00111100_01100100_10100000_0;
      patterns[15463] = 25'b00111100_01100101_10100001_0;
      patterns[15464] = 25'b00111100_01100110_10100010_0;
      patterns[15465] = 25'b00111100_01100111_10100011_0;
      patterns[15466] = 25'b00111100_01101000_10100100_0;
      patterns[15467] = 25'b00111100_01101001_10100101_0;
      patterns[15468] = 25'b00111100_01101010_10100110_0;
      patterns[15469] = 25'b00111100_01101011_10100111_0;
      patterns[15470] = 25'b00111100_01101100_10101000_0;
      patterns[15471] = 25'b00111100_01101101_10101001_0;
      patterns[15472] = 25'b00111100_01101110_10101010_0;
      patterns[15473] = 25'b00111100_01101111_10101011_0;
      patterns[15474] = 25'b00111100_01110000_10101100_0;
      patterns[15475] = 25'b00111100_01110001_10101101_0;
      patterns[15476] = 25'b00111100_01110010_10101110_0;
      patterns[15477] = 25'b00111100_01110011_10101111_0;
      patterns[15478] = 25'b00111100_01110100_10110000_0;
      patterns[15479] = 25'b00111100_01110101_10110001_0;
      patterns[15480] = 25'b00111100_01110110_10110010_0;
      patterns[15481] = 25'b00111100_01110111_10110011_0;
      patterns[15482] = 25'b00111100_01111000_10110100_0;
      patterns[15483] = 25'b00111100_01111001_10110101_0;
      patterns[15484] = 25'b00111100_01111010_10110110_0;
      patterns[15485] = 25'b00111100_01111011_10110111_0;
      patterns[15486] = 25'b00111100_01111100_10111000_0;
      patterns[15487] = 25'b00111100_01111101_10111001_0;
      patterns[15488] = 25'b00111100_01111110_10111010_0;
      patterns[15489] = 25'b00111100_01111111_10111011_0;
      patterns[15490] = 25'b00111100_10000000_10111100_0;
      patterns[15491] = 25'b00111100_10000001_10111101_0;
      patterns[15492] = 25'b00111100_10000010_10111110_0;
      patterns[15493] = 25'b00111100_10000011_10111111_0;
      patterns[15494] = 25'b00111100_10000100_11000000_0;
      patterns[15495] = 25'b00111100_10000101_11000001_0;
      patterns[15496] = 25'b00111100_10000110_11000010_0;
      patterns[15497] = 25'b00111100_10000111_11000011_0;
      patterns[15498] = 25'b00111100_10001000_11000100_0;
      patterns[15499] = 25'b00111100_10001001_11000101_0;
      patterns[15500] = 25'b00111100_10001010_11000110_0;
      patterns[15501] = 25'b00111100_10001011_11000111_0;
      patterns[15502] = 25'b00111100_10001100_11001000_0;
      patterns[15503] = 25'b00111100_10001101_11001001_0;
      patterns[15504] = 25'b00111100_10001110_11001010_0;
      patterns[15505] = 25'b00111100_10001111_11001011_0;
      patterns[15506] = 25'b00111100_10010000_11001100_0;
      patterns[15507] = 25'b00111100_10010001_11001101_0;
      patterns[15508] = 25'b00111100_10010010_11001110_0;
      patterns[15509] = 25'b00111100_10010011_11001111_0;
      patterns[15510] = 25'b00111100_10010100_11010000_0;
      patterns[15511] = 25'b00111100_10010101_11010001_0;
      patterns[15512] = 25'b00111100_10010110_11010010_0;
      patterns[15513] = 25'b00111100_10010111_11010011_0;
      patterns[15514] = 25'b00111100_10011000_11010100_0;
      patterns[15515] = 25'b00111100_10011001_11010101_0;
      patterns[15516] = 25'b00111100_10011010_11010110_0;
      patterns[15517] = 25'b00111100_10011011_11010111_0;
      patterns[15518] = 25'b00111100_10011100_11011000_0;
      patterns[15519] = 25'b00111100_10011101_11011001_0;
      patterns[15520] = 25'b00111100_10011110_11011010_0;
      patterns[15521] = 25'b00111100_10011111_11011011_0;
      patterns[15522] = 25'b00111100_10100000_11011100_0;
      patterns[15523] = 25'b00111100_10100001_11011101_0;
      patterns[15524] = 25'b00111100_10100010_11011110_0;
      patterns[15525] = 25'b00111100_10100011_11011111_0;
      patterns[15526] = 25'b00111100_10100100_11100000_0;
      patterns[15527] = 25'b00111100_10100101_11100001_0;
      patterns[15528] = 25'b00111100_10100110_11100010_0;
      patterns[15529] = 25'b00111100_10100111_11100011_0;
      patterns[15530] = 25'b00111100_10101000_11100100_0;
      patterns[15531] = 25'b00111100_10101001_11100101_0;
      patterns[15532] = 25'b00111100_10101010_11100110_0;
      patterns[15533] = 25'b00111100_10101011_11100111_0;
      patterns[15534] = 25'b00111100_10101100_11101000_0;
      patterns[15535] = 25'b00111100_10101101_11101001_0;
      patterns[15536] = 25'b00111100_10101110_11101010_0;
      patterns[15537] = 25'b00111100_10101111_11101011_0;
      patterns[15538] = 25'b00111100_10110000_11101100_0;
      patterns[15539] = 25'b00111100_10110001_11101101_0;
      patterns[15540] = 25'b00111100_10110010_11101110_0;
      patterns[15541] = 25'b00111100_10110011_11101111_0;
      patterns[15542] = 25'b00111100_10110100_11110000_0;
      patterns[15543] = 25'b00111100_10110101_11110001_0;
      patterns[15544] = 25'b00111100_10110110_11110010_0;
      patterns[15545] = 25'b00111100_10110111_11110011_0;
      patterns[15546] = 25'b00111100_10111000_11110100_0;
      patterns[15547] = 25'b00111100_10111001_11110101_0;
      patterns[15548] = 25'b00111100_10111010_11110110_0;
      patterns[15549] = 25'b00111100_10111011_11110111_0;
      patterns[15550] = 25'b00111100_10111100_11111000_0;
      patterns[15551] = 25'b00111100_10111101_11111001_0;
      patterns[15552] = 25'b00111100_10111110_11111010_0;
      patterns[15553] = 25'b00111100_10111111_11111011_0;
      patterns[15554] = 25'b00111100_11000000_11111100_0;
      patterns[15555] = 25'b00111100_11000001_11111101_0;
      patterns[15556] = 25'b00111100_11000010_11111110_0;
      patterns[15557] = 25'b00111100_11000011_11111111_0;
      patterns[15558] = 25'b00111100_11000100_00000000_1;
      patterns[15559] = 25'b00111100_11000101_00000001_1;
      patterns[15560] = 25'b00111100_11000110_00000010_1;
      patterns[15561] = 25'b00111100_11000111_00000011_1;
      patterns[15562] = 25'b00111100_11001000_00000100_1;
      patterns[15563] = 25'b00111100_11001001_00000101_1;
      patterns[15564] = 25'b00111100_11001010_00000110_1;
      patterns[15565] = 25'b00111100_11001011_00000111_1;
      patterns[15566] = 25'b00111100_11001100_00001000_1;
      patterns[15567] = 25'b00111100_11001101_00001001_1;
      patterns[15568] = 25'b00111100_11001110_00001010_1;
      patterns[15569] = 25'b00111100_11001111_00001011_1;
      patterns[15570] = 25'b00111100_11010000_00001100_1;
      patterns[15571] = 25'b00111100_11010001_00001101_1;
      patterns[15572] = 25'b00111100_11010010_00001110_1;
      patterns[15573] = 25'b00111100_11010011_00001111_1;
      patterns[15574] = 25'b00111100_11010100_00010000_1;
      patterns[15575] = 25'b00111100_11010101_00010001_1;
      patterns[15576] = 25'b00111100_11010110_00010010_1;
      patterns[15577] = 25'b00111100_11010111_00010011_1;
      patterns[15578] = 25'b00111100_11011000_00010100_1;
      patterns[15579] = 25'b00111100_11011001_00010101_1;
      patterns[15580] = 25'b00111100_11011010_00010110_1;
      patterns[15581] = 25'b00111100_11011011_00010111_1;
      patterns[15582] = 25'b00111100_11011100_00011000_1;
      patterns[15583] = 25'b00111100_11011101_00011001_1;
      patterns[15584] = 25'b00111100_11011110_00011010_1;
      patterns[15585] = 25'b00111100_11011111_00011011_1;
      patterns[15586] = 25'b00111100_11100000_00011100_1;
      patterns[15587] = 25'b00111100_11100001_00011101_1;
      patterns[15588] = 25'b00111100_11100010_00011110_1;
      patterns[15589] = 25'b00111100_11100011_00011111_1;
      patterns[15590] = 25'b00111100_11100100_00100000_1;
      patterns[15591] = 25'b00111100_11100101_00100001_1;
      patterns[15592] = 25'b00111100_11100110_00100010_1;
      patterns[15593] = 25'b00111100_11100111_00100011_1;
      patterns[15594] = 25'b00111100_11101000_00100100_1;
      patterns[15595] = 25'b00111100_11101001_00100101_1;
      patterns[15596] = 25'b00111100_11101010_00100110_1;
      patterns[15597] = 25'b00111100_11101011_00100111_1;
      patterns[15598] = 25'b00111100_11101100_00101000_1;
      patterns[15599] = 25'b00111100_11101101_00101001_1;
      patterns[15600] = 25'b00111100_11101110_00101010_1;
      patterns[15601] = 25'b00111100_11101111_00101011_1;
      patterns[15602] = 25'b00111100_11110000_00101100_1;
      patterns[15603] = 25'b00111100_11110001_00101101_1;
      patterns[15604] = 25'b00111100_11110010_00101110_1;
      patterns[15605] = 25'b00111100_11110011_00101111_1;
      patterns[15606] = 25'b00111100_11110100_00110000_1;
      patterns[15607] = 25'b00111100_11110101_00110001_1;
      patterns[15608] = 25'b00111100_11110110_00110010_1;
      patterns[15609] = 25'b00111100_11110111_00110011_1;
      patterns[15610] = 25'b00111100_11111000_00110100_1;
      patterns[15611] = 25'b00111100_11111001_00110101_1;
      patterns[15612] = 25'b00111100_11111010_00110110_1;
      patterns[15613] = 25'b00111100_11111011_00110111_1;
      patterns[15614] = 25'b00111100_11111100_00111000_1;
      patterns[15615] = 25'b00111100_11111101_00111001_1;
      patterns[15616] = 25'b00111100_11111110_00111010_1;
      patterns[15617] = 25'b00111100_11111111_00111011_1;
      patterns[15618] = 25'b00111101_00000000_00111101_0;
      patterns[15619] = 25'b00111101_00000001_00111110_0;
      patterns[15620] = 25'b00111101_00000010_00111111_0;
      patterns[15621] = 25'b00111101_00000011_01000000_0;
      patterns[15622] = 25'b00111101_00000100_01000001_0;
      patterns[15623] = 25'b00111101_00000101_01000010_0;
      patterns[15624] = 25'b00111101_00000110_01000011_0;
      patterns[15625] = 25'b00111101_00000111_01000100_0;
      patterns[15626] = 25'b00111101_00001000_01000101_0;
      patterns[15627] = 25'b00111101_00001001_01000110_0;
      patterns[15628] = 25'b00111101_00001010_01000111_0;
      patterns[15629] = 25'b00111101_00001011_01001000_0;
      patterns[15630] = 25'b00111101_00001100_01001001_0;
      patterns[15631] = 25'b00111101_00001101_01001010_0;
      patterns[15632] = 25'b00111101_00001110_01001011_0;
      patterns[15633] = 25'b00111101_00001111_01001100_0;
      patterns[15634] = 25'b00111101_00010000_01001101_0;
      patterns[15635] = 25'b00111101_00010001_01001110_0;
      patterns[15636] = 25'b00111101_00010010_01001111_0;
      patterns[15637] = 25'b00111101_00010011_01010000_0;
      patterns[15638] = 25'b00111101_00010100_01010001_0;
      patterns[15639] = 25'b00111101_00010101_01010010_0;
      patterns[15640] = 25'b00111101_00010110_01010011_0;
      patterns[15641] = 25'b00111101_00010111_01010100_0;
      patterns[15642] = 25'b00111101_00011000_01010101_0;
      patterns[15643] = 25'b00111101_00011001_01010110_0;
      patterns[15644] = 25'b00111101_00011010_01010111_0;
      patterns[15645] = 25'b00111101_00011011_01011000_0;
      patterns[15646] = 25'b00111101_00011100_01011001_0;
      patterns[15647] = 25'b00111101_00011101_01011010_0;
      patterns[15648] = 25'b00111101_00011110_01011011_0;
      patterns[15649] = 25'b00111101_00011111_01011100_0;
      patterns[15650] = 25'b00111101_00100000_01011101_0;
      patterns[15651] = 25'b00111101_00100001_01011110_0;
      patterns[15652] = 25'b00111101_00100010_01011111_0;
      patterns[15653] = 25'b00111101_00100011_01100000_0;
      patterns[15654] = 25'b00111101_00100100_01100001_0;
      patterns[15655] = 25'b00111101_00100101_01100010_0;
      patterns[15656] = 25'b00111101_00100110_01100011_0;
      patterns[15657] = 25'b00111101_00100111_01100100_0;
      patterns[15658] = 25'b00111101_00101000_01100101_0;
      patterns[15659] = 25'b00111101_00101001_01100110_0;
      patterns[15660] = 25'b00111101_00101010_01100111_0;
      patterns[15661] = 25'b00111101_00101011_01101000_0;
      patterns[15662] = 25'b00111101_00101100_01101001_0;
      patterns[15663] = 25'b00111101_00101101_01101010_0;
      patterns[15664] = 25'b00111101_00101110_01101011_0;
      patterns[15665] = 25'b00111101_00101111_01101100_0;
      patterns[15666] = 25'b00111101_00110000_01101101_0;
      patterns[15667] = 25'b00111101_00110001_01101110_0;
      patterns[15668] = 25'b00111101_00110010_01101111_0;
      patterns[15669] = 25'b00111101_00110011_01110000_0;
      patterns[15670] = 25'b00111101_00110100_01110001_0;
      patterns[15671] = 25'b00111101_00110101_01110010_0;
      patterns[15672] = 25'b00111101_00110110_01110011_0;
      patterns[15673] = 25'b00111101_00110111_01110100_0;
      patterns[15674] = 25'b00111101_00111000_01110101_0;
      patterns[15675] = 25'b00111101_00111001_01110110_0;
      patterns[15676] = 25'b00111101_00111010_01110111_0;
      patterns[15677] = 25'b00111101_00111011_01111000_0;
      patterns[15678] = 25'b00111101_00111100_01111001_0;
      patterns[15679] = 25'b00111101_00111101_01111010_0;
      patterns[15680] = 25'b00111101_00111110_01111011_0;
      patterns[15681] = 25'b00111101_00111111_01111100_0;
      patterns[15682] = 25'b00111101_01000000_01111101_0;
      patterns[15683] = 25'b00111101_01000001_01111110_0;
      patterns[15684] = 25'b00111101_01000010_01111111_0;
      patterns[15685] = 25'b00111101_01000011_10000000_0;
      patterns[15686] = 25'b00111101_01000100_10000001_0;
      patterns[15687] = 25'b00111101_01000101_10000010_0;
      patterns[15688] = 25'b00111101_01000110_10000011_0;
      patterns[15689] = 25'b00111101_01000111_10000100_0;
      patterns[15690] = 25'b00111101_01001000_10000101_0;
      patterns[15691] = 25'b00111101_01001001_10000110_0;
      patterns[15692] = 25'b00111101_01001010_10000111_0;
      patterns[15693] = 25'b00111101_01001011_10001000_0;
      patterns[15694] = 25'b00111101_01001100_10001001_0;
      patterns[15695] = 25'b00111101_01001101_10001010_0;
      patterns[15696] = 25'b00111101_01001110_10001011_0;
      patterns[15697] = 25'b00111101_01001111_10001100_0;
      patterns[15698] = 25'b00111101_01010000_10001101_0;
      patterns[15699] = 25'b00111101_01010001_10001110_0;
      patterns[15700] = 25'b00111101_01010010_10001111_0;
      patterns[15701] = 25'b00111101_01010011_10010000_0;
      patterns[15702] = 25'b00111101_01010100_10010001_0;
      patterns[15703] = 25'b00111101_01010101_10010010_0;
      patterns[15704] = 25'b00111101_01010110_10010011_0;
      patterns[15705] = 25'b00111101_01010111_10010100_0;
      patterns[15706] = 25'b00111101_01011000_10010101_0;
      patterns[15707] = 25'b00111101_01011001_10010110_0;
      patterns[15708] = 25'b00111101_01011010_10010111_0;
      patterns[15709] = 25'b00111101_01011011_10011000_0;
      patterns[15710] = 25'b00111101_01011100_10011001_0;
      patterns[15711] = 25'b00111101_01011101_10011010_0;
      patterns[15712] = 25'b00111101_01011110_10011011_0;
      patterns[15713] = 25'b00111101_01011111_10011100_0;
      patterns[15714] = 25'b00111101_01100000_10011101_0;
      patterns[15715] = 25'b00111101_01100001_10011110_0;
      patterns[15716] = 25'b00111101_01100010_10011111_0;
      patterns[15717] = 25'b00111101_01100011_10100000_0;
      patterns[15718] = 25'b00111101_01100100_10100001_0;
      patterns[15719] = 25'b00111101_01100101_10100010_0;
      patterns[15720] = 25'b00111101_01100110_10100011_0;
      patterns[15721] = 25'b00111101_01100111_10100100_0;
      patterns[15722] = 25'b00111101_01101000_10100101_0;
      patterns[15723] = 25'b00111101_01101001_10100110_0;
      patterns[15724] = 25'b00111101_01101010_10100111_0;
      patterns[15725] = 25'b00111101_01101011_10101000_0;
      patterns[15726] = 25'b00111101_01101100_10101001_0;
      patterns[15727] = 25'b00111101_01101101_10101010_0;
      patterns[15728] = 25'b00111101_01101110_10101011_0;
      patterns[15729] = 25'b00111101_01101111_10101100_0;
      patterns[15730] = 25'b00111101_01110000_10101101_0;
      patterns[15731] = 25'b00111101_01110001_10101110_0;
      patterns[15732] = 25'b00111101_01110010_10101111_0;
      patterns[15733] = 25'b00111101_01110011_10110000_0;
      patterns[15734] = 25'b00111101_01110100_10110001_0;
      patterns[15735] = 25'b00111101_01110101_10110010_0;
      patterns[15736] = 25'b00111101_01110110_10110011_0;
      patterns[15737] = 25'b00111101_01110111_10110100_0;
      patterns[15738] = 25'b00111101_01111000_10110101_0;
      patterns[15739] = 25'b00111101_01111001_10110110_0;
      patterns[15740] = 25'b00111101_01111010_10110111_0;
      patterns[15741] = 25'b00111101_01111011_10111000_0;
      patterns[15742] = 25'b00111101_01111100_10111001_0;
      patterns[15743] = 25'b00111101_01111101_10111010_0;
      patterns[15744] = 25'b00111101_01111110_10111011_0;
      patterns[15745] = 25'b00111101_01111111_10111100_0;
      patterns[15746] = 25'b00111101_10000000_10111101_0;
      patterns[15747] = 25'b00111101_10000001_10111110_0;
      patterns[15748] = 25'b00111101_10000010_10111111_0;
      patterns[15749] = 25'b00111101_10000011_11000000_0;
      patterns[15750] = 25'b00111101_10000100_11000001_0;
      patterns[15751] = 25'b00111101_10000101_11000010_0;
      patterns[15752] = 25'b00111101_10000110_11000011_0;
      patterns[15753] = 25'b00111101_10000111_11000100_0;
      patterns[15754] = 25'b00111101_10001000_11000101_0;
      patterns[15755] = 25'b00111101_10001001_11000110_0;
      patterns[15756] = 25'b00111101_10001010_11000111_0;
      patterns[15757] = 25'b00111101_10001011_11001000_0;
      patterns[15758] = 25'b00111101_10001100_11001001_0;
      patterns[15759] = 25'b00111101_10001101_11001010_0;
      patterns[15760] = 25'b00111101_10001110_11001011_0;
      patterns[15761] = 25'b00111101_10001111_11001100_0;
      patterns[15762] = 25'b00111101_10010000_11001101_0;
      patterns[15763] = 25'b00111101_10010001_11001110_0;
      patterns[15764] = 25'b00111101_10010010_11001111_0;
      patterns[15765] = 25'b00111101_10010011_11010000_0;
      patterns[15766] = 25'b00111101_10010100_11010001_0;
      patterns[15767] = 25'b00111101_10010101_11010010_0;
      patterns[15768] = 25'b00111101_10010110_11010011_0;
      patterns[15769] = 25'b00111101_10010111_11010100_0;
      patterns[15770] = 25'b00111101_10011000_11010101_0;
      patterns[15771] = 25'b00111101_10011001_11010110_0;
      patterns[15772] = 25'b00111101_10011010_11010111_0;
      patterns[15773] = 25'b00111101_10011011_11011000_0;
      patterns[15774] = 25'b00111101_10011100_11011001_0;
      patterns[15775] = 25'b00111101_10011101_11011010_0;
      patterns[15776] = 25'b00111101_10011110_11011011_0;
      patterns[15777] = 25'b00111101_10011111_11011100_0;
      patterns[15778] = 25'b00111101_10100000_11011101_0;
      patterns[15779] = 25'b00111101_10100001_11011110_0;
      patterns[15780] = 25'b00111101_10100010_11011111_0;
      patterns[15781] = 25'b00111101_10100011_11100000_0;
      patterns[15782] = 25'b00111101_10100100_11100001_0;
      patterns[15783] = 25'b00111101_10100101_11100010_0;
      patterns[15784] = 25'b00111101_10100110_11100011_0;
      patterns[15785] = 25'b00111101_10100111_11100100_0;
      patterns[15786] = 25'b00111101_10101000_11100101_0;
      patterns[15787] = 25'b00111101_10101001_11100110_0;
      patterns[15788] = 25'b00111101_10101010_11100111_0;
      patterns[15789] = 25'b00111101_10101011_11101000_0;
      patterns[15790] = 25'b00111101_10101100_11101001_0;
      patterns[15791] = 25'b00111101_10101101_11101010_0;
      patterns[15792] = 25'b00111101_10101110_11101011_0;
      patterns[15793] = 25'b00111101_10101111_11101100_0;
      patterns[15794] = 25'b00111101_10110000_11101101_0;
      patterns[15795] = 25'b00111101_10110001_11101110_0;
      patterns[15796] = 25'b00111101_10110010_11101111_0;
      patterns[15797] = 25'b00111101_10110011_11110000_0;
      patterns[15798] = 25'b00111101_10110100_11110001_0;
      patterns[15799] = 25'b00111101_10110101_11110010_0;
      patterns[15800] = 25'b00111101_10110110_11110011_0;
      patterns[15801] = 25'b00111101_10110111_11110100_0;
      patterns[15802] = 25'b00111101_10111000_11110101_0;
      patterns[15803] = 25'b00111101_10111001_11110110_0;
      patterns[15804] = 25'b00111101_10111010_11110111_0;
      patterns[15805] = 25'b00111101_10111011_11111000_0;
      patterns[15806] = 25'b00111101_10111100_11111001_0;
      patterns[15807] = 25'b00111101_10111101_11111010_0;
      patterns[15808] = 25'b00111101_10111110_11111011_0;
      patterns[15809] = 25'b00111101_10111111_11111100_0;
      patterns[15810] = 25'b00111101_11000000_11111101_0;
      patterns[15811] = 25'b00111101_11000001_11111110_0;
      patterns[15812] = 25'b00111101_11000010_11111111_0;
      patterns[15813] = 25'b00111101_11000011_00000000_1;
      patterns[15814] = 25'b00111101_11000100_00000001_1;
      patterns[15815] = 25'b00111101_11000101_00000010_1;
      patterns[15816] = 25'b00111101_11000110_00000011_1;
      patterns[15817] = 25'b00111101_11000111_00000100_1;
      patterns[15818] = 25'b00111101_11001000_00000101_1;
      patterns[15819] = 25'b00111101_11001001_00000110_1;
      patterns[15820] = 25'b00111101_11001010_00000111_1;
      patterns[15821] = 25'b00111101_11001011_00001000_1;
      patterns[15822] = 25'b00111101_11001100_00001001_1;
      patterns[15823] = 25'b00111101_11001101_00001010_1;
      patterns[15824] = 25'b00111101_11001110_00001011_1;
      patterns[15825] = 25'b00111101_11001111_00001100_1;
      patterns[15826] = 25'b00111101_11010000_00001101_1;
      patterns[15827] = 25'b00111101_11010001_00001110_1;
      patterns[15828] = 25'b00111101_11010010_00001111_1;
      patterns[15829] = 25'b00111101_11010011_00010000_1;
      patterns[15830] = 25'b00111101_11010100_00010001_1;
      patterns[15831] = 25'b00111101_11010101_00010010_1;
      patterns[15832] = 25'b00111101_11010110_00010011_1;
      patterns[15833] = 25'b00111101_11010111_00010100_1;
      patterns[15834] = 25'b00111101_11011000_00010101_1;
      patterns[15835] = 25'b00111101_11011001_00010110_1;
      patterns[15836] = 25'b00111101_11011010_00010111_1;
      patterns[15837] = 25'b00111101_11011011_00011000_1;
      patterns[15838] = 25'b00111101_11011100_00011001_1;
      patterns[15839] = 25'b00111101_11011101_00011010_1;
      patterns[15840] = 25'b00111101_11011110_00011011_1;
      patterns[15841] = 25'b00111101_11011111_00011100_1;
      patterns[15842] = 25'b00111101_11100000_00011101_1;
      patterns[15843] = 25'b00111101_11100001_00011110_1;
      patterns[15844] = 25'b00111101_11100010_00011111_1;
      patterns[15845] = 25'b00111101_11100011_00100000_1;
      patterns[15846] = 25'b00111101_11100100_00100001_1;
      patterns[15847] = 25'b00111101_11100101_00100010_1;
      patterns[15848] = 25'b00111101_11100110_00100011_1;
      patterns[15849] = 25'b00111101_11100111_00100100_1;
      patterns[15850] = 25'b00111101_11101000_00100101_1;
      patterns[15851] = 25'b00111101_11101001_00100110_1;
      patterns[15852] = 25'b00111101_11101010_00100111_1;
      patterns[15853] = 25'b00111101_11101011_00101000_1;
      patterns[15854] = 25'b00111101_11101100_00101001_1;
      patterns[15855] = 25'b00111101_11101101_00101010_1;
      patterns[15856] = 25'b00111101_11101110_00101011_1;
      patterns[15857] = 25'b00111101_11101111_00101100_1;
      patterns[15858] = 25'b00111101_11110000_00101101_1;
      patterns[15859] = 25'b00111101_11110001_00101110_1;
      patterns[15860] = 25'b00111101_11110010_00101111_1;
      patterns[15861] = 25'b00111101_11110011_00110000_1;
      patterns[15862] = 25'b00111101_11110100_00110001_1;
      patterns[15863] = 25'b00111101_11110101_00110010_1;
      patterns[15864] = 25'b00111101_11110110_00110011_1;
      patterns[15865] = 25'b00111101_11110111_00110100_1;
      patterns[15866] = 25'b00111101_11111000_00110101_1;
      patterns[15867] = 25'b00111101_11111001_00110110_1;
      patterns[15868] = 25'b00111101_11111010_00110111_1;
      patterns[15869] = 25'b00111101_11111011_00111000_1;
      patterns[15870] = 25'b00111101_11111100_00111001_1;
      patterns[15871] = 25'b00111101_11111101_00111010_1;
      patterns[15872] = 25'b00111101_11111110_00111011_1;
      patterns[15873] = 25'b00111101_11111111_00111100_1;
      patterns[15874] = 25'b00111110_00000000_00111110_0;
      patterns[15875] = 25'b00111110_00000001_00111111_0;
      patterns[15876] = 25'b00111110_00000010_01000000_0;
      patterns[15877] = 25'b00111110_00000011_01000001_0;
      patterns[15878] = 25'b00111110_00000100_01000010_0;
      patterns[15879] = 25'b00111110_00000101_01000011_0;
      patterns[15880] = 25'b00111110_00000110_01000100_0;
      patterns[15881] = 25'b00111110_00000111_01000101_0;
      patterns[15882] = 25'b00111110_00001000_01000110_0;
      patterns[15883] = 25'b00111110_00001001_01000111_0;
      patterns[15884] = 25'b00111110_00001010_01001000_0;
      patterns[15885] = 25'b00111110_00001011_01001001_0;
      patterns[15886] = 25'b00111110_00001100_01001010_0;
      patterns[15887] = 25'b00111110_00001101_01001011_0;
      patterns[15888] = 25'b00111110_00001110_01001100_0;
      patterns[15889] = 25'b00111110_00001111_01001101_0;
      patterns[15890] = 25'b00111110_00010000_01001110_0;
      patterns[15891] = 25'b00111110_00010001_01001111_0;
      patterns[15892] = 25'b00111110_00010010_01010000_0;
      patterns[15893] = 25'b00111110_00010011_01010001_0;
      patterns[15894] = 25'b00111110_00010100_01010010_0;
      patterns[15895] = 25'b00111110_00010101_01010011_0;
      patterns[15896] = 25'b00111110_00010110_01010100_0;
      patterns[15897] = 25'b00111110_00010111_01010101_0;
      patterns[15898] = 25'b00111110_00011000_01010110_0;
      patterns[15899] = 25'b00111110_00011001_01010111_0;
      patterns[15900] = 25'b00111110_00011010_01011000_0;
      patterns[15901] = 25'b00111110_00011011_01011001_0;
      patterns[15902] = 25'b00111110_00011100_01011010_0;
      patterns[15903] = 25'b00111110_00011101_01011011_0;
      patterns[15904] = 25'b00111110_00011110_01011100_0;
      patterns[15905] = 25'b00111110_00011111_01011101_0;
      patterns[15906] = 25'b00111110_00100000_01011110_0;
      patterns[15907] = 25'b00111110_00100001_01011111_0;
      patterns[15908] = 25'b00111110_00100010_01100000_0;
      patterns[15909] = 25'b00111110_00100011_01100001_0;
      patterns[15910] = 25'b00111110_00100100_01100010_0;
      patterns[15911] = 25'b00111110_00100101_01100011_0;
      patterns[15912] = 25'b00111110_00100110_01100100_0;
      patterns[15913] = 25'b00111110_00100111_01100101_0;
      patterns[15914] = 25'b00111110_00101000_01100110_0;
      patterns[15915] = 25'b00111110_00101001_01100111_0;
      patterns[15916] = 25'b00111110_00101010_01101000_0;
      patterns[15917] = 25'b00111110_00101011_01101001_0;
      patterns[15918] = 25'b00111110_00101100_01101010_0;
      patterns[15919] = 25'b00111110_00101101_01101011_0;
      patterns[15920] = 25'b00111110_00101110_01101100_0;
      patterns[15921] = 25'b00111110_00101111_01101101_0;
      patterns[15922] = 25'b00111110_00110000_01101110_0;
      patterns[15923] = 25'b00111110_00110001_01101111_0;
      patterns[15924] = 25'b00111110_00110010_01110000_0;
      patterns[15925] = 25'b00111110_00110011_01110001_0;
      patterns[15926] = 25'b00111110_00110100_01110010_0;
      patterns[15927] = 25'b00111110_00110101_01110011_0;
      patterns[15928] = 25'b00111110_00110110_01110100_0;
      patterns[15929] = 25'b00111110_00110111_01110101_0;
      patterns[15930] = 25'b00111110_00111000_01110110_0;
      patterns[15931] = 25'b00111110_00111001_01110111_0;
      patterns[15932] = 25'b00111110_00111010_01111000_0;
      patterns[15933] = 25'b00111110_00111011_01111001_0;
      patterns[15934] = 25'b00111110_00111100_01111010_0;
      patterns[15935] = 25'b00111110_00111101_01111011_0;
      patterns[15936] = 25'b00111110_00111110_01111100_0;
      patterns[15937] = 25'b00111110_00111111_01111101_0;
      patterns[15938] = 25'b00111110_01000000_01111110_0;
      patterns[15939] = 25'b00111110_01000001_01111111_0;
      patterns[15940] = 25'b00111110_01000010_10000000_0;
      patterns[15941] = 25'b00111110_01000011_10000001_0;
      patterns[15942] = 25'b00111110_01000100_10000010_0;
      patterns[15943] = 25'b00111110_01000101_10000011_0;
      patterns[15944] = 25'b00111110_01000110_10000100_0;
      patterns[15945] = 25'b00111110_01000111_10000101_0;
      patterns[15946] = 25'b00111110_01001000_10000110_0;
      patterns[15947] = 25'b00111110_01001001_10000111_0;
      patterns[15948] = 25'b00111110_01001010_10001000_0;
      patterns[15949] = 25'b00111110_01001011_10001001_0;
      patterns[15950] = 25'b00111110_01001100_10001010_0;
      patterns[15951] = 25'b00111110_01001101_10001011_0;
      patterns[15952] = 25'b00111110_01001110_10001100_0;
      patterns[15953] = 25'b00111110_01001111_10001101_0;
      patterns[15954] = 25'b00111110_01010000_10001110_0;
      patterns[15955] = 25'b00111110_01010001_10001111_0;
      patterns[15956] = 25'b00111110_01010010_10010000_0;
      patterns[15957] = 25'b00111110_01010011_10010001_0;
      patterns[15958] = 25'b00111110_01010100_10010010_0;
      patterns[15959] = 25'b00111110_01010101_10010011_0;
      patterns[15960] = 25'b00111110_01010110_10010100_0;
      patterns[15961] = 25'b00111110_01010111_10010101_0;
      patterns[15962] = 25'b00111110_01011000_10010110_0;
      patterns[15963] = 25'b00111110_01011001_10010111_0;
      patterns[15964] = 25'b00111110_01011010_10011000_0;
      patterns[15965] = 25'b00111110_01011011_10011001_0;
      patterns[15966] = 25'b00111110_01011100_10011010_0;
      patterns[15967] = 25'b00111110_01011101_10011011_0;
      patterns[15968] = 25'b00111110_01011110_10011100_0;
      patterns[15969] = 25'b00111110_01011111_10011101_0;
      patterns[15970] = 25'b00111110_01100000_10011110_0;
      patterns[15971] = 25'b00111110_01100001_10011111_0;
      patterns[15972] = 25'b00111110_01100010_10100000_0;
      patterns[15973] = 25'b00111110_01100011_10100001_0;
      patterns[15974] = 25'b00111110_01100100_10100010_0;
      patterns[15975] = 25'b00111110_01100101_10100011_0;
      patterns[15976] = 25'b00111110_01100110_10100100_0;
      patterns[15977] = 25'b00111110_01100111_10100101_0;
      patterns[15978] = 25'b00111110_01101000_10100110_0;
      patterns[15979] = 25'b00111110_01101001_10100111_0;
      patterns[15980] = 25'b00111110_01101010_10101000_0;
      patterns[15981] = 25'b00111110_01101011_10101001_0;
      patterns[15982] = 25'b00111110_01101100_10101010_0;
      patterns[15983] = 25'b00111110_01101101_10101011_0;
      patterns[15984] = 25'b00111110_01101110_10101100_0;
      patterns[15985] = 25'b00111110_01101111_10101101_0;
      patterns[15986] = 25'b00111110_01110000_10101110_0;
      patterns[15987] = 25'b00111110_01110001_10101111_0;
      patterns[15988] = 25'b00111110_01110010_10110000_0;
      patterns[15989] = 25'b00111110_01110011_10110001_0;
      patterns[15990] = 25'b00111110_01110100_10110010_0;
      patterns[15991] = 25'b00111110_01110101_10110011_0;
      patterns[15992] = 25'b00111110_01110110_10110100_0;
      patterns[15993] = 25'b00111110_01110111_10110101_0;
      patterns[15994] = 25'b00111110_01111000_10110110_0;
      patterns[15995] = 25'b00111110_01111001_10110111_0;
      patterns[15996] = 25'b00111110_01111010_10111000_0;
      patterns[15997] = 25'b00111110_01111011_10111001_0;
      patterns[15998] = 25'b00111110_01111100_10111010_0;
      patterns[15999] = 25'b00111110_01111101_10111011_0;
      patterns[16000] = 25'b00111110_01111110_10111100_0;
      patterns[16001] = 25'b00111110_01111111_10111101_0;
      patterns[16002] = 25'b00111110_10000000_10111110_0;
      patterns[16003] = 25'b00111110_10000001_10111111_0;
      patterns[16004] = 25'b00111110_10000010_11000000_0;
      patterns[16005] = 25'b00111110_10000011_11000001_0;
      patterns[16006] = 25'b00111110_10000100_11000010_0;
      patterns[16007] = 25'b00111110_10000101_11000011_0;
      patterns[16008] = 25'b00111110_10000110_11000100_0;
      patterns[16009] = 25'b00111110_10000111_11000101_0;
      patterns[16010] = 25'b00111110_10001000_11000110_0;
      patterns[16011] = 25'b00111110_10001001_11000111_0;
      patterns[16012] = 25'b00111110_10001010_11001000_0;
      patterns[16013] = 25'b00111110_10001011_11001001_0;
      patterns[16014] = 25'b00111110_10001100_11001010_0;
      patterns[16015] = 25'b00111110_10001101_11001011_0;
      patterns[16016] = 25'b00111110_10001110_11001100_0;
      patterns[16017] = 25'b00111110_10001111_11001101_0;
      patterns[16018] = 25'b00111110_10010000_11001110_0;
      patterns[16019] = 25'b00111110_10010001_11001111_0;
      patterns[16020] = 25'b00111110_10010010_11010000_0;
      patterns[16021] = 25'b00111110_10010011_11010001_0;
      patterns[16022] = 25'b00111110_10010100_11010010_0;
      patterns[16023] = 25'b00111110_10010101_11010011_0;
      patterns[16024] = 25'b00111110_10010110_11010100_0;
      patterns[16025] = 25'b00111110_10010111_11010101_0;
      patterns[16026] = 25'b00111110_10011000_11010110_0;
      patterns[16027] = 25'b00111110_10011001_11010111_0;
      patterns[16028] = 25'b00111110_10011010_11011000_0;
      patterns[16029] = 25'b00111110_10011011_11011001_0;
      patterns[16030] = 25'b00111110_10011100_11011010_0;
      patterns[16031] = 25'b00111110_10011101_11011011_0;
      patterns[16032] = 25'b00111110_10011110_11011100_0;
      patterns[16033] = 25'b00111110_10011111_11011101_0;
      patterns[16034] = 25'b00111110_10100000_11011110_0;
      patterns[16035] = 25'b00111110_10100001_11011111_0;
      patterns[16036] = 25'b00111110_10100010_11100000_0;
      patterns[16037] = 25'b00111110_10100011_11100001_0;
      patterns[16038] = 25'b00111110_10100100_11100010_0;
      patterns[16039] = 25'b00111110_10100101_11100011_0;
      patterns[16040] = 25'b00111110_10100110_11100100_0;
      patterns[16041] = 25'b00111110_10100111_11100101_0;
      patterns[16042] = 25'b00111110_10101000_11100110_0;
      patterns[16043] = 25'b00111110_10101001_11100111_0;
      patterns[16044] = 25'b00111110_10101010_11101000_0;
      patterns[16045] = 25'b00111110_10101011_11101001_0;
      patterns[16046] = 25'b00111110_10101100_11101010_0;
      patterns[16047] = 25'b00111110_10101101_11101011_0;
      patterns[16048] = 25'b00111110_10101110_11101100_0;
      patterns[16049] = 25'b00111110_10101111_11101101_0;
      patterns[16050] = 25'b00111110_10110000_11101110_0;
      patterns[16051] = 25'b00111110_10110001_11101111_0;
      patterns[16052] = 25'b00111110_10110010_11110000_0;
      patterns[16053] = 25'b00111110_10110011_11110001_0;
      patterns[16054] = 25'b00111110_10110100_11110010_0;
      patterns[16055] = 25'b00111110_10110101_11110011_0;
      patterns[16056] = 25'b00111110_10110110_11110100_0;
      patterns[16057] = 25'b00111110_10110111_11110101_0;
      patterns[16058] = 25'b00111110_10111000_11110110_0;
      patterns[16059] = 25'b00111110_10111001_11110111_0;
      patterns[16060] = 25'b00111110_10111010_11111000_0;
      patterns[16061] = 25'b00111110_10111011_11111001_0;
      patterns[16062] = 25'b00111110_10111100_11111010_0;
      patterns[16063] = 25'b00111110_10111101_11111011_0;
      patterns[16064] = 25'b00111110_10111110_11111100_0;
      patterns[16065] = 25'b00111110_10111111_11111101_0;
      patterns[16066] = 25'b00111110_11000000_11111110_0;
      patterns[16067] = 25'b00111110_11000001_11111111_0;
      patterns[16068] = 25'b00111110_11000010_00000000_1;
      patterns[16069] = 25'b00111110_11000011_00000001_1;
      patterns[16070] = 25'b00111110_11000100_00000010_1;
      patterns[16071] = 25'b00111110_11000101_00000011_1;
      patterns[16072] = 25'b00111110_11000110_00000100_1;
      patterns[16073] = 25'b00111110_11000111_00000101_1;
      patterns[16074] = 25'b00111110_11001000_00000110_1;
      patterns[16075] = 25'b00111110_11001001_00000111_1;
      patterns[16076] = 25'b00111110_11001010_00001000_1;
      patterns[16077] = 25'b00111110_11001011_00001001_1;
      patterns[16078] = 25'b00111110_11001100_00001010_1;
      patterns[16079] = 25'b00111110_11001101_00001011_1;
      patterns[16080] = 25'b00111110_11001110_00001100_1;
      patterns[16081] = 25'b00111110_11001111_00001101_1;
      patterns[16082] = 25'b00111110_11010000_00001110_1;
      patterns[16083] = 25'b00111110_11010001_00001111_1;
      patterns[16084] = 25'b00111110_11010010_00010000_1;
      patterns[16085] = 25'b00111110_11010011_00010001_1;
      patterns[16086] = 25'b00111110_11010100_00010010_1;
      patterns[16087] = 25'b00111110_11010101_00010011_1;
      patterns[16088] = 25'b00111110_11010110_00010100_1;
      patterns[16089] = 25'b00111110_11010111_00010101_1;
      patterns[16090] = 25'b00111110_11011000_00010110_1;
      patterns[16091] = 25'b00111110_11011001_00010111_1;
      patterns[16092] = 25'b00111110_11011010_00011000_1;
      patterns[16093] = 25'b00111110_11011011_00011001_1;
      patterns[16094] = 25'b00111110_11011100_00011010_1;
      patterns[16095] = 25'b00111110_11011101_00011011_1;
      patterns[16096] = 25'b00111110_11011110_00011100_1;
      patterns[16097] = 25'b00111110_11011111_00011101_1;
      patterns[16098] = 25'b00111110_11100000_00011110_1;
      patterns[16099] = 25'b00111110_11100001_00011111_1;
      patterns[16100] = 25'b00111110_11100010_00100000_1;
      patterns[16101] = 25'b00111110_11100011_00100001_1;
      patterns[16102] = 25'b00111110_11100100_00100010_1;
      patterns[16103] = 25'b00111110_11100101_00100011_1;
      patterns[16104] = 25'b00111110_11100110_00100100_1;
      patterns[16105] = 25'b00111110_11100111_00100101_1;
      patterns[16106] = 25'b00111110_11101000_00100110_1;
      patterns[16107] = 25'b00111110_11101001_00100111_1;
      patterns[16108] = 25'b00111110_11101010_00101000_1;
      patterns[16109] = 25'b00111110_11101011_00101001_1;
      patterns[16110] = 25'b00111110_11101100_00101010_1;
      patterns[16111] = 25'b00111110_11101101_00101011_1;
      patterns[16112] = 25'b00111110_11101110_00101100_1;
      patterns[16113] = 25'b00111110_11101111_00101101_1;
      patterns[16114] = 25'b00111110_11110000_00101110_1;
      patterns[16115] = 25'b00111110_11110001_00101111_1;
      patterns[16116] = 25'b00111110_11110010_00110000_1;
      patterns[16117] = 25'b00111110_11110011_00110001_1;
      patterns[16118] = 25'b00111110_11110100_00110010_1;
      patterns[16119] = 25'b00111110_11110101_00110011_1;
      patterns[16120] = 25'b00111110_11110110_00110100_1;
      patterns[16121] = 25'b00111110_11110111_00110101_1;
      patterns[16122] = 25'b00111110_11111000_00110110_1;
      patterns[16123] = 25'b00111110_11111001_00110111_1;
      patterns[16124] = 25'b00111110_11111010_00111000_1;
      patterns[16125] = 25'b00111110_11111011_00111001_1;
      patterns[16126] = 25'b00111110_11111100_00111010_1;
      patterns[16127] = 25'b00111110_11111101_00111011_1;
      patterns[16128] = 25'b00111110_11111110_00111100_1;
      patterns[16129] = 25'b00111110_11111111_00111101_1;
      patterns[16130] = 25'b00111111_00000000_00111111_0;
      patterns[16131] = 25'b00111111_00000001_01000000_0;
      patterns[16132] = 25'b00111111_00000010_01000001_0;
      patterns[16133] = 25'b00111111_00000011_01000010_0;
      patterns[16134] = 25'b00111111_00000100_01000011_0;
      patterns[16135] = 25'b00111111_00000101_01000100_0;
      patterns[16136] = 25'b00111111_00000110_01000101_0;
      patterns[16137] = 25'b00111111_00000111_01000110_0;
      patterns[16138] = 25'b00111111_00001000_01000111_0;
      patterns[16139] = 25'b00111111_00001001_01001000_0;
      patterns[16140] = 25'b00111111_00001010_01001001_0;
      patterns[16141] = 25'b00111111_00001011_01001010_0;
      patterns[16142] = 25'b00111111_00001100_01001011_0;
      patterns[16143] = 25'b00111111_00001101_01001100_0;
      patterns[16144] = 25'b00111111_00001110_01001101_0;
      patterns[16145] = 25'b00111111_00001111_01001110_0;
      patterns[16146] = 25'b00111111_00010000_01001111_0;
      patterns[16147] = 25'b00111111_00010001_01010000_0;
      patterns[16148] = 25'b00111111_00010010_01010001_0;
      patterns[16149] = 25'b00111111_00010011_01010010_0;
      patterns[16150] = 25'b00111111_00010100_01010011_0;
      patterns[16151] = 25'b00111111_00010101_01010100_0;
      patterns[16152] = 25'b00111111_00010110_01010101_0;
      patterns[16153] = 25'b00111111_00010111_01010110_0;
      patterns[16154] = 25'b00111111_00011000_01010111_0;
      patterns[16155] = 25'b00111111_00011001_01011000_0;
      patterns[16156] = 25'b00111111_00011010_01011001_0;
      patterns[16157] = 25'b00111111_00011011_01011010_0;
      patterns[16158] = 25'b00111111_00011100_01011011_0;
      patterns[16159] = 25'b00111111_00011101_01011100_0;
      patterns[16160] = 25'b00111111_00011110_01011101_0;
      patterns[16161] = 25'b00111111_00011111_01011110_0;
      patterns[16162] = 25'b00111111_00100000_01011111_0;
      patterns[16163] = 25'b00111111_00100001_01100000_0;
      patterns[16164] = 25'b00111111_00100010_01100001_0;
      patterns[16165] = 25'b00111111_00100011_01100010_0;
      patterns[16166] = 25'b00111111_00100100_01100011_0;
      patterns[16167] = 25'b00111111_00100101_01100100_0;
      patterns[16168] = 25'b00111111_00100110_01100101_0;
      patterns[16169] = 25'b00111111_00100111_01100110_0;
      patterns[16170] = 25'b00111111_00101000_01100111_0;
      patterns[16171] = 25'b00111111_00101001_01101000_0;
      patterns[16172] = 25'b00111111_00101010_01101001_0;
      patterns[16173] = 25'b00111111_00101011_01101010_0;
      patterns[16174] = 25'b00111111_00101100_01101011_0;
      patterns[16175] = 25'b00111111_00101101_01101100_0;
      patterns[16176] = 25'b00111111_00101110_01101101_0;
      patterns[16177] = 25'b00111111_00101111_01101110_0;
      patterns[16178] = 25'b00111111_00110000_01101111_0;
      patterns[16179] = 25'b00111111_00110001_01110000_0;
      patterns[16180] = 25'b00111111_00110010_01110001_0;
      patterns[16181] = 25'b00111111_00110011_01110010_0;
      patterns[16182] = 25'b00111111_00110100_01110011_0;
      patterns[16183] = 25'b00111111_00110101_01110100_0;
      patterns[16184] = 25'b00111111_00110110_01110101_0;
      patterns[16185] = 25'b00111111_00110111_01110110_0;
      patterns[16186] = 25'b00111111_00111000_01110111_0;
      patterns[16187] = 25'b00111111_00111001_01111000_0;
      patterns[16188] = 25'b00111111_00111010_01111001_0;
      patterns[16189] = 25'b00111111_00111011_01111010_0;
      patterns[16190] = 25'b00111111_00111100_01111011_0;
      patterns[16191] = 25'b00111111_00111101_01111100_0;
      patterns[16192] = 25'b00111111_00111110_01111101_0;
      patterns[16193] = 25'b00111111_00111111_01111110_0;
      patterns[16194] = 25'b00111111_01000000_01111111_0;
      patterns[16195] = 25'b00111111_01000001_10000000_0;
      patterns[16196] = 25'b00111111_01000010_10000001_0;
      patterns[16197] = 25'b00111111_01000011_10000010_0;
      patterns[16198] = 25'b00111111_01000100_10000011_0;
      patterns[16199] = 25'b00111111_01000101_10000100_0;
      patterns[16200] = 25'b00111111_01000110_10000101_0;
      patterns[16201] = 25'b00111111_01000111_10000110_0;
      patterns[16202] = 25'b00111111_01001000_10000111_0;
      patterns[16203] = 25'b00111111_01001001_10001000_0;
      patterns[16204] = 25'b00111111_01001010_10001001_0;
      patterns[16205] = 25'b00111111_01001011_10001010_0;
      patterns[16206] = 25'b00111111_01001100_10001011_0;
      patterns[16207] = 25'b00111111_01001101_10001100_0;
      patterns[16208] = 25'b00111111_01001110_10001101_0;
      patterns[16209] = 25'b00111111_01001111_10001110_0;
      patterns[16210] = 25'b00111111_01010000_10001111_0;
      patterns[16211] = 25'b00111111_01010001_10010000_0;
      patterns[16212] = 25'b00111111_01010010_10010001_0;
      patterns[16213] = 25'b00111111_01010011_10010010_0;
      patterns[16214] = 25'b00111111_01010100_10010011_0;
      patterns[16215] = 25'b00111111_01010101_10010100_0;
      patterns[16216] = 25'b00111111_01010110_10010101_0;
      patterns[16217] = 25'b00111111_01010111_10010110_0;
      patterns[16218] = 25'b00111111_01011000_10010111_0;
      patterns[16219] = 25'b00111111_01011001_10011000_0;
      patterns[16220] = 25'b00111111_01011010_10011001_0;
      patterns[16221] = 25'b00111111_01011011_10011010_0;
      patterns[16222] = 25'b00111111_01011100_10011011_0;
      patterns[16223] = 25'b00111111_01011101_10011100_0;
      patterns[16224] = 25'b00111111_01011110_10011101_0;
      patterns[16225] = 25'b00111111_01011111_10011110_0;
      patterns[16226] = 25'b00111111_01100000_10011111_0;
      patterns[16227] = 25'b00111111_01100001_10100000_0;
      patterns[16228] = 25'b00111111_01100010_10100001_0;
      patterns[16229] = 25'b00111111_01100011_10100010_0;
      patterns[16230] = 25'b00111111_01100100_10100011_0;
      patterns[16231] = 25'b00111111_01100101_10100100_0;
      patterns[16232] = 25'b00111111_01100110_10100101_0;
      patterns[16233] = 25'b00111111_01100111_10100110_0;
      patterns[16234] = 25'b00111111_01101000_10100111_0;
      patterns[16235] = 25'b00111111_01101001_10101000_0;
      patterns[16236] = 25'b00111111_01101010_10101001_0;
      patterns[16237] = 25'b00111111_01101011_10101010_0;
      patterns[16238] = 25'b00111111_01101100_10101011_0;
      patterns[16239] = 25'b00111111_01101101_10101100_0;
      patterns[16240] = 25'b00111111_01101110_10101101_0;
      patterns[16241] = 25'b00111111_01101111_10101110_0;
      patterns[16242] = 25'b00111111_01110000_10101111_0;
      patterns[16243] = 25'b00111111_01110001_10110000_0;
      patterns[16244] = 25'b00111111_01110010_10110001_0;
      patterns[16245] = 25'b00111111_01110011_10110010_0;
      patterns[16246] = 25'b00111111_01110100_10110011_0;
      patterns[16247] = 25'b00111111_01110101_10110100_0;
      patterns[16248] = 25'b00111111_01110110_10110101_0;
      patterns[16249] = 25'b00111111_01110111_10110110_0;
      patterns[16250] = 25'b00111111_01111000_10110111_0;
      patterns[16251] = 25'b00111111_01111001_10111000_0;
      patterns[16252] = 25'b00111111_01111010_10111001_0;
      patterns[16253] = 25'b00111111_01111011_10111010_0;
      patterns[16254] = 25'b00111111_01111100_10111011_0;
      patterns[16255] = 25'b00111111_01111101_10111100_0;
      patterns[16256] = 25'b00111111_01111110_10111101_0;
      patterns[16257] = 25'b00111111_01111111_10111110_0;
      patterns[16258] = 25'b00111111_10000000_10111111_0;
      patterns[16259] = 25'b00111111_10000001_11000000_0;
      patterns[16260] = 25'b00111111_10000010_11000001_0;
      patterns[16261] = 25'b00111111_10000011_11000010_0;
      patterns[16262] = 25'b00111111_10000100_11000011_0;
      patterns[16263] = 25'b00111111_10000101_11000100_0;
      patterns[16264] = 25'b00111111_10000110_11000101_0;
      patterns[16265] = 25'b00111111_10000111_11000110_0;
      patterns[16266] = 25'b00111111_10001000_11000111_0;
      patterns[16267] = 25'b00111111_10001001_11001000_0;
      patterns[16268] = 25'b00111111_10001010_11001001_0;
      patterns[16269] = 25'b00111111_10001011_11001010_0;
      patterns[16270] = 25'b00111111_10001100_11001011_0;
      patterns[16271] = 25'b00111111_10001101_11001100_0;
      patterns[16272] = 25'b00111111_10001110_11001101_0;
      patterns[16273] = 25'b00111111_10001111_11001110_0;
      patterns[16274] = 25'b00111111_10010000_11001111_0;
      patterns[16275] = 25'b00111111_10010001_11010000_0;
      patterns[16276] = 25'b00111111_10010010_11010001_0;
      patterns[16277] = 25'b00111111_10010011_11010010_0;
      patterns[16278] = 25'b00111111_10010100_11010011_0;
      patterns[16279] = 25'b00111111_10010101_11010100_0;
      patterns[16280] = 25'b00111111_10010110_11010101_0;
      patterns[16281] = 25'b00111111_10010111_11010110_0;
      patterns[16282] = 25'b00111111_10011000_11010111_0;
      patterns[16283] = 25'b00111111_10011001_11011000_0;
      patterns[16284] = 25'b00111111_10011010_11011001_0;
      patterns[16285] = 25'b00111111_10011011_11011010_0;
      patterns[16286] = 25'b00111111_10011100_11011011_0;
      patterns[16287] = 25'b00111111_10011101_11011100_0;
      patterns[16288] = 25'b00111111_10011110_11011101_0;
      patterns[16289] = 25'b00111111_10011111_11011110_0;
      patterns[16290] = 25'b00111111_10100000_11011111_0;
      patterns[16291] = 25'b00111111_10100001_11100000_0;
      patterns[16292] = 25'b00111111_10100010_11100001_0;
      patterns[16293] = 25'b00111111_10100011_11100010_0;
      patterns[16294] = 25'b00111111_10100100_11100011_0;
      patterns[16295] = 25'b00111111_10100101_11100100_0;
      patterns[16296] = 25'b00111111_10100110_11100101_0;
      patterns[16297] = 25'b00111111_10100111_11100110_0;
      patterns[16298] = 25'b00111111_10101000_11100111_0;
      patterns[16299] = 25'b00111111_10101001_11101000_0;
      patterns[16300] = 25'b00111111_10101010_11101001_0;
      patterns[16301] = 25'b00111111_10101011_11101010_0;
      patterns[16302] = 25'b00111111_10101100_11101011_0;
      patterns[16303] = 25'b00111111_10101101_11101100_0;
      patterns[16304] = 25'b00111111_10101110_11101101_0;
      patterns[16305] = 25'b00111111_10101111_11101110_0;
      patterns[16306] = 25'b00111111_10110000_11101111_0;
      patterns[16307] = 25'b00111111_10110001_11110000_0;
      patterns[16308] = 25'b00111111_10110010_11110001_0;
      patterns[16309] = 25'b00111111_10110011_11110010_0;
      patterns[16310] = 25'b00111111_10110100_11110011_0;
      patterns[16311] = 25'b00111111_10110101_11110100_0;
      patterns[16312] = 25'b00111111_10110110_11110101_0;
      patterns[16313] = 25'b00111111_10110111_11110110_0;
      patterns[16314] = 25'b00111111_10111000_11110111_0;
      patterns[16315] = 25'b00111111_10111001_11111000_0;
      patterns[16316] = 25'b00111111_10111010_11111001_0;
      patterns[16317] = 25'b00111111_10111011_11111010_0;
      patterns[16318] = 25'b00111111_10111100_11111011_0;
      patterns[16319] = 25'b00111111_10111101_11111100_0;
      patterns[16320] = 25'b00111111_10111110_11111101_0;
      patterns[16321] = 25'b00111111_10111111_11111110_0;
      patterns[16322] = 25'b00111111_11000000_11111111_0;
      patterns[16323] = 25'b00111111_11000001_00000000_1;
      patterns[16324] = 25'b00111111_11000010_00000001_1;
      patterns[16325] = 25'b00111111_11000011_00000010_1;
      patterns[16326] = 25'b00111111_11000100_00000011_1;
      patterns[16327] = 25'b00111111_11000101_00000100_1;
      patterns[16328] = 25'b00111111_11000110_00000101_1;
      patterns[16329] = 25'b00111111_11000111_00000110_1;
      patterns[16330] = 25'b00111111_11001000_00000111_1;
      patterns[16331] = 25'b00111111_11001001_00001000_1;
      patterns[16332] = 25'b00111111_11001010_00001001_1;
      patterns[16333] = 25'b00111111_11001011_00001010_1;
      patterns[16334] = 25'b00111111_11001100_00001011_1;
      patterns[16335] = 25'b00111111_11001101_00001100_1;
      patterns[16336] = 25'b00111111_11001110_00001101_1;
      patterns[16337] = 25'b00111111_11001111_00001110_1;
      patterns[16338] = 25'b00111111_11010000_00001111_1;
      patterns[16339] = 25'b00111111_11010001_00010000_1;
      patterns[16340] = 25'b00111111_11010010_00010001_1;
      patterns[16341] = 25'b00111111_11010011_00010010_1;
      patterns[16342] = 25'b00111111_11010100_00010011_1;
      patterns[16343] = 25'b00111111_11010101_00010100_1;
      patterns[16344] = 25'b00111111_11010110_00010101_1;
      patterns[16345] = 25'b00111111_11010111_00010110_1;
      patterns[16346] = 25'b00111111_11011000_00010111_1;
      patterns[16347] = 25'b00111111_11011001_00011000_1;
      patterns[16348] = 25'b00111111_11011010_00011001_1;
      patterns[16349] = 25'b00111111_11011011_00011010_1;
      patterns[16350] = 25'b00111111_11011100_00011011_1;
      patterns[16351] = 25'b00111111_11011101_00011100_1;
      patterns[16352] = 25'b00111111_11011110_00011101_1;
      patterns[16353] = 25'b00111111_11011111_00011110_1;
      patterns[16354] = 25'b00111111_11100000_00011111_1;
      patterns[16355] = 25'b00111111_11100001_00100000_1;
      patterns[16356] = 25'b00111111_11100010_00100001_1;
      patterns[16357] = 25'b00111111_11100011_00100010_1;
      patterns[16358] = 25'b00111111_11100100_00100011_1;
      patterns[16359] = 25'b00111111_11100101_00100100_1;
      patterns[16360] = 25'b00111111_11100110_00100101_1;
      patterns[16361] = 25'b00111111_11100111_00100110_1;
      patterns[16362] = 25'b00111111_11101000_00100111_1;
      patterns[16363] = 25'b00111111_11101001_00101000_1;
      patterns[16364] = 25'b00111111_11101010_00101001_1;
      patterns[16365] = 25'b00111111_11101011_00101010_1;
      patterns[16366] = 25'b00111111_11101100_00101011_1;
      patterns[16367] = 25'b00111111_11101101_00101100_1;
      patterns[16368] = 25'b00111111_11101110_00101101_1;
      patterns[16369] = 25'b00111111_11101111_00101110_1;
      patterns[16370] = 25'b00111111_11110000_00101111_1;
      patterns[16371] = 25'b00111111_11110001_00110000_1;
      patterns[16372] = 25'b00111111_11110010_00110001_1;
      patterns[16373] = 25'b00111111_11110011_00110010_1;
      patterns[16374] = 25'b00111111_11110100_00110011_1;
      patterns[16375] = 25'b00111111_11110101_00110100_1;
      patterns[16376] = 25'b00111111_11110110_00110101_1;
      patterns[16377] = 25'b00111111_11110111_00110110_1;
      patterns[16378] = 25'b00111111_11111000_00110111_1;
      patterns[16379] = 25'b00111111_11111001_00111000_1;
      patterns[16380] = 25'b00111111_11111010_00111001_1;
      patterns[16381] = 25'b00111111_11111011_00111010_1;
      patterns[16382] = 25'b00111111_11111100_00111011_1;
      patterns[16383] = 25'b00111111_11111101_00111100_1;
      patterns[16384] = 25'b00111111_11111110_00111101_1;
      patterns[16385] = 25'b00111111_11111111_00111110_1;
      patterns[16386] = 25'b01000000_00000000_01000000_0;
      patterns[16387] = 25'b01000000_00000001_01000001_0;
      patterns[16388] = 25'b01000000_00000010_01000010_0;
      patterns[16389] = 25'b01000000_00000011_01000011_0;
      patterns[16390] = 25'b01000000_00000100_01000100_0;
      patterns[16391] = 25'b01000000_00000101_01000101_0;
      patterns[16392] = 25'b01000000_00000110_01000110_0;
      patterns[16393] = 25'b01000000_00000111_01000111_0;
      patterns[16394] = 25'b01000000_00001000_01001000_0;
      patterns[16395] = 25'b01000000_00001001_01001001_0;
      patterns[16396] = 25'b01000000_00001010_01001010_0;
      patterns[16397] = 25'b01000000_00001011_01001011_0;
      patterns[16398] = 25'b01000000_00001100_01001100_0;
      patterns[16399] = 25'b01000000_00001101_01001101_0;
      patterns[16400] = 25'b01000000_00001110_01001110_0;
      patterns[16401] = 25'b01000000_00001111_01001111_0;
      patterns[16402] = 25'b01000000_00010000_01010000_0;
      patterns[16403] = 25'b01000000_00010001_01010001_0;
      patterns[16404] = 25'b01000000_00010010_01010010_0;
      patterns[16405] = 25'b01000000_00010011_01010011_0;
      patterns[16406] = 25'b01000000_00010100_01010100_0;
      patterns[16407] = 25'b01000000_00010101_01010101_0;
      patterns[16408] = 25'b01000000_00010110_01010110_0;
      patterns[16409] = 25'b01000000_00010111_01010111_0;
      patterns[16410] = 25'b01000000_00011000_01011000_0;
      patterns[16411] = 25'b01000000_00011001_01011001_0;
      patterns[16412] = 25'b01000000_00011010_01011010_0;
      patterns[16413] = 25'b01000000_00011011_01011011_0;
      patterns[16414] = 25'b01000000_00011100_01011100_0;
      patterns[16415] = 25'b01000000_00011101_01011101_0;
      patterns[16416] = 25'b01000000_00011110_01011110_0;
      patterns[16417] = 25'b01000000_00011111_01011111_0;
      patterns[16418] = 25'b01000000_00100000_01100000_0;
      patterns[16419] = 25'b01000000_00100001_01100001_0;
      patterns[16420] = 25'b01000000_00100010_01100010_0;
      patterns[16421] = 25'b01000000_00100011_01100011_0;
      patterns[16422] = 25'b01000000_00100100_01100100_0;
      patterns[16423] = 25'b01000000_00100101_01100101_0;
      patterns[16424] = 25'b01000000_00100110_01100110_0;
      patterns[16425] = 25'b01000000_00100111_01100111_0;
      patterns[16426] = 25'b01000000_00101000_01101000_0;
      patterns[16427] = 25'b01000000_00101001_01101001_0;
      patterns[16428] = 25'b01000000_00101010_01101010_0;
      patterns[16429] = 25'b01000000_00101011_01101011_0;
      patterns[16430] = 25'b01000000_00101100_01101100_0;
      patterns[16431] = 25'b01000000_00101101_01101101_0;
      patterns[16432] = 25'b01000000_00101110_01101110_0;
      patterns[16433] = 25'b01000000_00101111_01101111_0;
      patterns[16434] = 25'b01000000_00110000_01110000_0;
      patterns[16435] = 25'b01000000_00110001_01110001_0;
      patterns[16436] = 25'b01000000_00110010_01110010_0;
      patterns[16437] = 25'b01000000_00110011_01110011_0;
      patterns[16438] = 25'b01000000_00110100_01110100_0;
      patterns[16439] = 25'b01000000_00110101_01110101_0;
      patterns[16440] = 25'b01000000_00110110_01110110_0;
      patterns[16441] = 25'b01000000_00110111_01110111_0;
      patterns[16442] = 25'b01000000_00111000_01111000_0;
      patterns[16443] = 25'b01000000_00111001_01111001_0;
      patterns[16444] = 25'b01000000_00111010_01111010_0;
      patterns[16445] = 25'b01000000_00111011_01111011_0;
      patterns[16446] = 25'b01000000_00111100_01111100_0;
      patterns[16447] = 25'b01000000_00111101_01111101_0;
      patterns[16448] = 25'b01000000_00111110_01111110_0;
      patterns[16449] = 25'b01000000_00111111_01111111_0;
      patterns[16450] = 25'b01000000_01000000_10000000_0;
      patterns[16451] = 25'b01000000_01000001_10000001_0;
      patterns[16452] = 25'b01000000_01000010_10000010_0;
      patterns[16453] = 25'b01000000_01000011_10000011_0;
      patterns[16454] = 25'b01000000_01000100_10000100_0;
      patterns[16455] = 25'b01000000_01000101_10000101_0;
      patterns[16456] = 25'b01000000_01000110_10000110_0;
      patterns[16457] = 25'b01000000_01000111_10000111_0;
      patterns[16458] = 25'b01000000_01001000_10001000_0;
      patterns[16459] = 25'b01000000_01001001_10001001_0;
      patterns[16460] = 25'b01000000_01001010_10001010_0;
      patterns[16461] = 25'b01000000_01001011_10001011_0;
      patterns[16462] = 25'b01000000_01001100_10001100_0;
      patterns[16463] = 25'b01000000_01001101_10001101_0;
      patterns[16464] = 25'b01000000_01001110_10001110_0;
      patterns[16465] = 25'b01000000_01001111_10001111_0;
      patterns[16466] = 25'b01000000_01010000_10010000_0;
      patterns[16467] = 25'b01000000_01010001_10010001_0;
      patterns[16468] = 25'b01000000_01010010_10010010_0;
      patterns[16469] = 25'b01000000_01010011_10010011_0;
      patterns[16470] = 25'b01000000_01010100_10010100_0;
      patterns[16471] = 25'b01000000_01010101_10010101_0;
      patterns[16472] = 25'b01000000_01010110_10010110_0;
      patterns[16473] = 25'b01000000_01010111_10010111_0;
      patterns[16474] = 25'b01000000_01011000_10011000_0;
      patterns[16475] = 25'b01000000_01011001_10011001_0;
      patterns[16476] = 25'b01000000_01011010_10011010_0;
      patterns[16477] = 25'b01000000_01011011_10011011_0;
      patterns[16478] = 25'b01000000_01011100_10011100_0;
      patterns[16479] = 25'b01000000_01011101_10011101_0;
      patterns[16480] = 25'b01000000_01011110_10011110_0;
      patterns[16481] = 25'b01000000_01011111_10011111_0;
      patterns[16482] = 25'b01000000_01100000_10100000_0;
      patterns[16483] = 25'b01000000_01100001_10100001_0;
      patterns[16484] = 25'b01000000_01100010_10100010_0;
      patterns[16485] = 25'b01000000_01100011_10100011_0;
      patterns[16486] = 25'b01000000_01100100_10100100_0;
      patterns[16487] = 25'b01000000_01100101_10100101_0;
      patterns[16488] = 25'b01000000_01100110_10100110_0;
      patterns[16489] = 25'b01000000_01100111_10100111_0;
      patterns[16490] = 25'b01000000_01101000_10101000_0;
      patterns[16491] = 25'b01000000_01101001_10101001_0;
      patterns[16492] = 25'b01000000_01101010_10101010_0;
      patterns[16493] = 25'b01000000_01101011_10101011_0;
      patterns[16494] = 25'b01000000_01101100_10101100_0;
      patterns[16495] = 25'b01000000_01101101_10101101_0;
      patterns[16496] = 25'b01000000_01101110_10101110_0;
      patterns[16497] = 25'b01000000_01101111_10101111_0;
      patterns[16498] = 25'b01000000_01110000_10110000_0;
      patterns[16499] = 25'b01000000_01110001_10110001_0;
      patterns[16500] = 25'b01000000_01110010_10110010_0;
      patterns[16501] = 25'b01000000_01110011_10110011_0;
      patterns[16502] = 25'b01000000_01110100_10110100_0;
      patterns[16503] = 25'b01000000_01110101_10110101_0;
      patterns[16504] = 25'b01000000_01110110_10110110_0;
      patterns[16505] = 25'b01000000_01110111_10110111_0;
      patterns[16506] = 25'b01000000_01111000_10111000_0;
      patterns[16507] = 25'b01000000_01111001_10111001_0;
      patterns[16508] = 25'b01000000_01111010_10111010_0;
      patterns[16509] = 25'b01000000_01111011_10111011_0;
      patterns[16510] = 25'b01000000_01111100_10111100_0;
      patterns[16511] = 25'b01000000_01111101_10111101_0;
      patterns[16512] = 25'b01000000_01111110_10111110_0;
      patterns[16513] = 25'b01000000_01111111_10111111_0;
      patterns[16514] = 25'b01000000_10000000_11000000_0;
      patterns[16515] = 25'b01000000_10000001_11000001_0;
      patterns[16516] = 25'b01000000_10000010_11000010_0;
      patterns[16517] = 25'b01000000_10000011_11000011_0;
      patterns[16518] = 25'b01000000_10000100_11000100_0;
      patterns[16519] = 25'b01000000_10000101_11000101_0;
      patterns[16520] = 25'b01000000_10000110_11000110_0;
      patterns[16521] = 25'b01000000_10000111_11000111_0;
      patterns[16522] = 25'b01000000_10001000_11001000_0;
      patterns[16523] = 25'b01000000_10001001_11001001_0;
      patterns[16524] = 25'b01000000_10001010_11001010_0;
      patterns[16525] = 25'b01000000_10001011_11001011_0;
      patterns[16526] = 25'b01000000_10001100_11001100_0;
      patterns[16527] = 25'b01000000_10001101_11001101_0;
      patterns[16528] = 25'b01000000_10001110_11001110_0;
      patterns[16529] = 25'b01000000_10001111_11001111_0;
      patterns[16530] = 25'b01000000_10010000_11010000_0;
      patterns[16531] = 25'b01000000_10010001_11010001_0;
      patterns[16532] = 25'b01000000_10010010_11010010_0;
      patterns[16533] = 25'b01000000_10010011_11010011_0;
      patterns[16534] = 25'b01000000_10010100_11010100_0;
      patterns[16535] = 25'b01000000_10010101_11010101_0;
      patterns[16536] = 25'b01000000_10010110_11010110_0;
      patterns[16537] = 25'b01000000_10010111_11010111_0;
      patterns[16538] = 25'b01000000_10011000_11011000_0;
      patterns[16539] = 25'b01000000_10011001_11011001_0;
      patterns[16540] = 25'b01000000_10011010_11011010_0;
      patterns[16541] = 25'b01000000_10011011_11011011_0;
      patterns[16542] = 25'b01000000_10011100_11011100_0;
      patterns[16543] = 25'b01000000_10011101_11011101_0;
      patterns[16544] = 25'b01000000_10011110_11011110_0;
      patterns[16545] = 25'b01000000_10011111_11011111_0;
      patterns[16546] = 25'b01000000_10100000_11100000_0;
      patterns[16547] = 25'b01000000_10100001_11100001_0;
      patterns[16548] = 25'b01000000_10100010_11100010_0;
      patterns[16549] = 25'b01000000_10100011_11100011_0;
      patterns[16550] = 25'b01000000_10100100_11100100_0;
      patterns[16551] = 25'b01000000_10100101_11100101_0;
      patterns[16552] = 25'b01000000_10100110_11100110_0;
      patterns[16553] = 25'b01000000_10100111_11100111_0;
      patterns[16554] = 25'b01000000_10101000_11101000_0;
      patterns[16555] = 25'b01000000_10101001_11101001_0;
      patterns[16556] = 25'b01000000_10101010_11101010_0;
      patterns[16557] = 25'b01000000_10101011_11101011_0;
      patterns[16558] = 25'b01000000_10101100_11101100_0;
      patterns[16559] = 25'b01000000_10101101_11101101_0;
      patterns[16560] = 25'b01000000_10101110_11101110_0;
      patterns[16561] = 25'b01000000_10101111_11101111_0;
      patterns[16562] = 25'b01000000_10110000_11110000_0;
      patterns[16563] = 25'b01000000_10110001_11110001_0;
      patterns[16564] = 25'b01000000_10110010_11110010_0;
      patterns[16565] = 25'b01000000_10110011_11110011_0;
      patterns[16566] = 25'b01000000_10110100_11110100_0;
      patterns[16567] = 25'b01000000_10110101_11110101_0;
      patterns[16568] = 25'b01000000_10110110_11110110_0;
      patterns[16569] = 25'b01000000_10110111_11110111_0;
      patterns[16570] = 25'b01000000_10111000_11111000_0;
      patterns[16571] = 25'b01000000_10111001_11111001_0;
      patterns[16572] = 25'b01000000_10111010_11111010_0;
      patterns[16573] = 25'b01000000_10111011_11111011_0;
      patterns[16574] = 25'b01000000_10111100_11111100_0;
      patterns[16575] = 25'b01000000_10111101_11111101_0;
      patterns[16576] = 25'b01000000_10111110_11111110_0;
      patterns[16577] = 25'b01000000_10111111_11111111_0;
      patterns[16578] = 25'b01000000_11000000_00000000_1;
      patterns[16579] = 25'b01000000_11000001_00000001_1;
      patterns[16580] = 25'b01000000_11000010_00000010_1;
      patterns[16581] = 25'b01000000_11000011_00000011_1;
      patterns[16582] = 25'b01000000_11000100_00000100_1;
      patterns[16583] = 25'b01000000_11000101_00000101_1;
      patterns[16584] = 25'b01000000_11000110_00000110_1;
      patterns[16585] = 25'b01000000_11000111_00000111_1;
      patterns[16586] = 25'b01000000_11001000_00001000_1;
      patterns[16587] = 25'b01000000_11001001_00001001_1;
      patterns[16588] = 25'b01000000_11001010_00001010_1;
      patterns[16589] = 25'b01000000_11001011_00001011_1;
      patterns[16590] = 25'b01000000_11001100_00001100_1;
      patterns[16591] = 25'b01000000_11001101_00001101_1;
      patterns[16592] = 25'b01000000_11001110_00001110_1;
      patterns[16593] = 25'b01000000_11001111_00001111_1;
      patterns[16594] = 25'b01000000_11010000_00010000_1;
      patterns[16595] = 25'b01000000_11010001_00010001_1;
      patterns[16596] = 25'b01000000_11010010_00010010_1;
      patterns[16597] = 25'b01000000_11010011_00010011_1;
      patterns[16598] = 25'b01000000_11010100_00010100_1;
      patterns[16599] = 25'b01000000_11010101_00010101_1;
      patterns[16600] = 25'b01000000_11010110_00010110_1;
      patterns[16601] = 25'b01000000_11010111_00010111_1;
      patterns[16602] = 25'b01000000_11011000_00011000_1;
      patterns[16603] = 25'b01000000_11011001_00011001_1;
      patterns[16604] = 25'b01000000_11011010_00011010_1;
      patterns[16605] = 25'b01000000_11011011_00011011_1;
      patterns[16606] = 25'b01000000_11011100_00011100_1;
      patterns[16607] = 25'b01000000_11011101_00011101_1;
      patterns[16608] = 25'b01000000_11011110_00011110_1;
      patterns[16609] = 25'b01000000_11011111_00011111_1;
      patterns[16610] = 25'b01000000_11100000_00100000_1;
      patterns[16611] = 25'b01000000_11100001_00100001_1;
      patterns[16612] = 25'b01000000_11100010_00100010_1;
      patterns[16613] = 25'b01000000_11100011_00100011_1;
      patterns[16614] = 25'b01000000_11100100_00100100_1;
      patterns[16615] = 25'b01000000_11100101_00100101_1;
      patterns[16616] = 25'b01000000_11100110_00100110_1;
      patterns[16617] = 25'b01000000_11100111_00100111_1;
      patterns[16618] = 25'b01000000_11101000_00101000_1;
      patterns[16619] = 25'b01000000_11101001_00101001_1;
      patterns[16620] = 25'b01000000_11101010_00101010_1;
      patterns[16621] = 25'b01000000_11101011_00101011_1;
      patterns[16622] = 25'b01000000_11101100_00101100_1;
      patterns[16623] = 25'b01000000_11101101_00101101_1;
      patterns[16624] = 25'b01000000_11101110_00101110_1;
      patterns[16625] = 25'b01000000_11101111_00101111_1;
      patterns[16626] = 25'b01000000_11110000_00110000_1;
      patterns[16627] = 25'b01000000_11110001_00110001_1;
      patterns[16628] = 25'b01000000_11110010_00110010_1;
      patterns[16629] = 25'b01000000_11110011_00110011_1;
      patterns[16630] = 25'b01000000_11110100_00110100_1;
      patterns[16631] = 25'b01000000_11110101_00110101_1;
      patterns[16632] = 25'b01000000_11110110_00110110_1;
      patterns[16633] = 25'b01000000_11110111_00110111_1;
      patterns[16634] = 25'b01000000_11111000_00111000_1;
      patterns[16635] = 25'b01000000_11111001_00111001_1;
      patterns[16636] = 25'b01000000_11111010_00111010_1;
      patterns[16637] = 25'b01000000_11111011_00111011_1;
      patterns[16638] = 25'b01000000_11111100_00111100_1;
      patterns[16639] = 25'b01000000_11111101_00111101_1;
      patterns[16640] = 25'b01000000_11111110_00111110_1;
      patterns[16641] = 25'b01000000_11111111_00111111_1;
      patterns[16642] = 25'b01000001_00000000_01000001_0;
      patterns[16643] = 25'b01000001_00000001_01000010_0;
      patterns[16644] = 25'b01000001_00000010_01000011_0;
      patterns[16645] = 25'b01000001_00000011_01000100_0;
      patterns[16646] = 25'b01000001_00000100_01000101_0;
      patterns[16647] = 25'b01000001_00000101_01000110_0;
      patterns[16648] = 25'b01000001_00000110_01000111_0;
      patterns[16649] = 25'b01000001_00000111_01001000_0;
      patterns[16650] = 25'b01000001_00001000_01001001_0;
      patterns[16651] = 25'b01000001_00001001_01001010_0;
      patterns[16652] = 25'b01000001_00001010_01001011_0;
      patterns[16653] = 25'b01000001_00001011_01001100_0;
      patterns[16654] = 25'b01000001_00001100_01001101_0;
      patterns[16655] = 25'b01000001_00001101_01001110_0;
      patterns[16656] = 25'b01000001_00001110_01001111_0;
      patterns[16657] = 25'b01000001_00001111_01010000_0;
      patterns[16658] = 25'b01000001_00010000_01010001_0;
      patterns[16659] = 25'b01000001_00010001_01010010_0;
      patterns[16660] = 25'b01000001_00010010_01010011_0;
      patterns[16661] = 25'b01000001_00010011_01010100_0;
      patterns[16662] = 25'b01000001_00010100_01010101_0;
      patterns[16663] = 25'b01000001_00010101_01010110_0;
      patterns[16664] = 25'b01000001_00010110_01010111_0;
      patterns[16665] = 25'b01000001_00010111_01011000_0;
      patterns[16666] = 25'b01000001_00011000_01011001_0;
      patterns[16667] = 25'b01000001_00011001_01011010_0;
      patterns[16668] = 25'b01000001_00011010_01011011_0;
      patterns[16669] = 25'b01000001_00011011_01011100_0;
      patterns[16670] = 25'b01000001_00011100_01011101_0;
      patterns[16671] = 25'b01000001_00011101_01011110_0;
      patterns[16672] = 25'b01000001_00011110_01011111_0;
      patterns[16673] = 25'b01000001_00011111_01100000_0;
      patterns[16674] = 25'b01000001_00100000_01100001_0;
      patterns[16675] = 25'b01000001_00100001_01100010_0;
      patterns[16676] = 25'b01000001_00100010_01100011_0;
      patterns[16677] = 25'b01000001_00100011_01100100_0;
      patterns[16678] = 25'b01000001_00100100_01100101_0;
      patterns[16679] = 25'b01000001_00100101_01100110_0;
      patterns[16680] = 25'b01000001_00100110_01100111_0;
      patterns[16681] = 25'b01000001_00100111_01101000_0;
      patterns[16682] = 25'b01000001_00101000_01101001_0;
      patterns[16683] = 25'b01000001_00101001_01101010_0;
      patterns[16684] = 25'b01000001_00101010_01101011_0;
      patterns[16685] = 25'b01000001_00101011_01101100_0;
      patterns[16686] = 25'b01000001_00101100_01101101_0;
      patterns[16687] = 25'b01000001_00101101_01101110_0;
      patterns[16688] = 25'b01000001_00101110_01101111_0;
      patterns[16689] = 25'b01000001_00101111_01110000_0;
      patterns[16690] = 25'b01000001_00110000_01110001_0;
      patterns[16691] = 25'b01000001_00110001_01110010_0;
      patterns[16692] = 25'b01000001_00110010_01110011_0;
      patterns[16693] = 25'b01000001_00110011_01110100_0;
      patterns[16694] = 25'b01000001_00110100_01110101_0;
      patterns[16695] = 25'b01000001_00110101_01110110_0;
      patterns[16696] = 25'b01000001_00110110_01110111_0;
      patterns[16697] = 25'b01000001_00110111_01111000_0;
      patterns[16698] = 25'b01000001_00111000_01111001_0;
      patterns[16699] = 25'b01000001_00111001_01111010_0;
      patterns[16700] = 25'b01000001_00111010_01111011_0;
      patterns[16701] = 25'b01000001_00111011_01111100_0;
      patterns[16702] = 25'b01000001_00111100_01111101_0;
      patterns[16703] = 25'b01000001_00111101_01111110_0;
      patterns[16704] = 25'b01000001_00111110_01111111_0;
      patterns[16705] = 25'b01000001_00111111_10000000_0;
      patterns[16706] = 25'b01000001_01000000_10000001_0;
      patterns[16707] = 25'b01000001_01000001_10000010_0;
      patterns[16708] = 25'b01000001_01000010_10000011_0;
      patterns[16709] = 25'b01000001_01000011_10000100_0;
      patterns[16710] = 25'b01000001_01000100_10000101_0;
      patterns[16711] = 25'b01000001_01000101_10000110_0;
      patterns[16712] = 25'b01000001_01000110_10000111_0;
      patterns[16713] = 25'b01000001_01000111_10001000_0;
      patterns[16714] = 25'b01000001_01001000_10001001_0;
      patterns[16715] = 25'b01000001_01001001_10001010_0;
      patterns[16716] = 25'b01000001_01001010_10001011_0;
      patterns[16717] = 25'b01000001_01001011_10001100_0;
      patterns[16718] = 25'b01000001_01001100_10001101_0;
      patterns[16719] = 25'b01000001_01001101_10001110_0;
      patterns[16720] = 25'b01000001_01001110_10001111_0;
      patterns[16721] = 25'b01000001_01001111_10010000_0;
      patterns[16722] = 25'b01000001_01010000_10010001_0;
      patterns[16723] = 25'b01000001_01010001_10010010_0;
      patterns[16724] = 25'b01000001_01010010_10010011_0;
      patterns[16725] = 25'b01000001_01010011_10010100_0;
      patterns[16726] = 25'b01000001_01010100_10010101_0;
      patterns[16727] = 25'b01000001_01010101_10010110_0;
      patterns[16728] = 25'b01000001_01010110_10010111_0;
      patterns[16729] = 25'b01000001_01010111_10011000_0;
      patterns[16730] = 25'b01000001_01011000_10011001_0;
      patterns[16731] = 25'b01000001_01011001_10011010_0;
      patterns[16732] = 25'b01000001_01011010_10011011_0;
      patterns[16733] = 25'b01000001_01011011_10011100_0;
      patterns[16734] = 25'b01000001_01011100_10011101_0;
      patterns[16735] = 25'b01000001_01011101_10011110_0;
      patterns[16736] = 25'b01000001_01011110_10011111_0;
      patterns[16737] = 25'b01000001_01011111_10100000_0;
      patterns[16738] = 25'b01000001_01100000_10100001_0;
      patterns[16739] = 25'b01000001_01100001_10100010_0;
      patterns[16740] = 25'b01000001_01100010_10100011_0;
      patterns[16741] = 25'b01000001_01100011_10100100_0;
      patterns[16742] = 25'b01000001_01100100_10100101_0;
      patterns[16743] = 25'b01000001_01100101_10100110_0;
      patterns[16744] = 25'b01000001_01100110_10100111_0;
      patterns[16745] = 25'b01000001_01100111_10101000_0;
      patterns[16746] = 25'b01000001_01101000_10101001_0;
      patterns[16747] = 25'b01000001_01101001_10101010_0;
      patterns[16748] = 25'b01000001_01101010_10101011_0;
      patterns[16749] = 25'b01000001_01101011_10101100_0;
      patterns[16750] = 25'b01000001_01101100_10101101_0;
      patterns[16751] = 25'b01000001_01101101_10101110_0;
      patterns[16752] = 25'b01000001_01101110_10101111_0;
      patterns[16753] = 25'b01000001_01101111_10110000_0;
      patterns[16754] = 25'b01000001_01110000_10110001_0;
      patterns[16755] = 25'b01000001_01110001_10110010_0;
      patterns[16756] = 25'b01000001_01110010_10110011_0;
      patterns[16757] = 25'b01000001_01110011_10110100_0;
      patterns[16758] = 25'b01000001_01110100_10110101_0;
      patterns[16759] = 25'b01000001_01110101_10110110_0;
      patterns[16760] = 25'b01000001_01110110_10110111_0;
      patterns[16761] = 25'b01000001_01110111_10111000_0;
      patterns[16762] = 25'b01000001_01111000_10111001_0;
      patterns[16763] = 25'b01000001_01111001_10111010_0;
      patterns[16764] = 25'b01000001_01111010_10111011_0;
      patterns[16765] = 25'b01000001_01111011_10111100_0;
      patterns[16766] = 25'b01000001_01111100_10111101_0;
      patterns[16767] = 25'b01000001_01111101_10111110_0;
      patterns[16768] = 25'b01000001_01111110_10111111_0;
      patterns[16769] = 25'b01000001_01111111_11000000_0;
      patterns[16770] = 25'b01000001_10000000_11000001_0;
      patterns[16771] = 25'b01000001_10000001_11000010_0;
      patterns[16772] = 25'b01000001_10000010_11000011_0;
      patterns[16773] = 25'b01000001_10000011_11000100_0;
      patterns[16774] = 25'b01000001_10000100_11000101_0;
      patterns[16775] = 25'b01000001_10000101_11000110_0;
      patterns[16776] = 25'b01000001_10000110_11000111_0;
      patterns[16777] = 25'b01000001_10000111_11001000_0;
      patterns[16778] = 25'b01000001_10001000_11001001_0;
      patterns[16779] = 25'b01000001_10001001_11001010_0;
      patterns[16780] = 25'b01000001_10001010_11001011_0;
      patterns[16781] = 25'b01000001_10001011_11001100_0;
      patterns[16782] = 25'b01000001_10001100_11001101_0;
      patterns[16783] = 25'b01000001_10001101_11001110_0;
      patterns[16784] = 25'b01000001_10001110_11001111_0;
      patterns[16785] = 25'b01000001_10001111_11010000_0;
      patterns[16786] = 25'b01000001_10010000_11010001_0;
      patterns[16787] = 25'b01000001_10010001_11010010_0;
      patterns[16788] = 25'b01000001_10010010_11010011_0;
      patterns[16789] = 25'b01000001_10010011_11010100_0;
      patterns[16790] = 25'b01000001_10010100_11010101_0;
      patterns[16791] = 25'b01000001_10010101_11010110_0;
      patterns[16792] = 25'b01000001_10010110_11010111_0;
      patterns[16793] = 25'b01000001_10010111_11011000_0;
      patterns[16794] = 25'b01000001_10011000_11011001_0;
      patterns[16795] = 25'b01000001_10011001_11011010_0;
      patterns[16796] = 25'b01000001_10011010_11011011_0;
      patterns[16797] = 25'b01000001_10011011_11011100_0;
      patterns[16798] = 25'b01000001_10011100_11011101_0;
      patterns[16799] = 25'b01000001_10011101_11011110_0;
      patterns[16800] = 25'b01000001_10011110_11011111_0;
      patterns[16801] = 25'b01000001_10011111_11100000_0;
      patterns[16802] = 25'b01000001_10100000_11100001_0;
      patterns[16803] = 25'b01000001_10100001_11100010_0;
      patterns[16804] = 25'b01000001_10100010_11100011_0;
      patterns[16805] = 25'b01000001_10100011_11100100_0;
      patterns[16806] = 25'b01000001_10100100_11100101_0;
      patterns[16807] = 25'b01000001_10100101_11100110_0;
      patterns[16808] = 25'b01000001_10100110_11100111_0;
      patterns[16809] = 25'b01000001_10100111_11101000_0;
      patterns[16810] = 25'b01000001_10101000_11101001_0;
      patterns[16811] = 25'b01000001_10101001_11101010_0;
      patterns[16812] = 25'b01000001_10101010_11101011_0;
      patterns[16813] = 25'b01000001_10101011_11101100_0;
      patterns[16814] = 25'b01000001_10101100_11101101_0;
      patterns[16815] = 25'b01000001_10101101_11101110_0;
      patterns[16816] = 25'b01000001_10101110_11101111_0;
      patterns[16817] = 25'b01000001_10101111_11110000_0;
      patterns[16818] = 25'b01000001_10110000_11110001_0;
      patterns[16819] = 25'b01000001_10110001_11110010_0;
      patterns[16820] = 25'b01000001_10110010_11110011_0;
      patterns[16821] = 25'b01000001_10110011_11110100_0;
      patterns[16822] = 25'b01000001_10110100_11110101_0;
      patterns[16823] = 25'b01000001_10110101_11110110_0;
      patterns[16824] = 25'b01000001_10110110_11110111_0;
      patterns[16825] = 25'b01000001_10110111_11111000_0;
      patterns[16826] = 25'b01000001_10111000_11111001_0;
      patterns[16827] = 25'b01000001_10111001_11111010_0;
      patterns[16828] = 25'b01000001_10111010_11111011_0;
      patterns[16829] = 25'b01000001_10111011_11111100_0;
      patterns[16830] = 25'b01000001_10111100_11111101_0;
      patterns[16831] = 25'b01000001_10111101_11111110_0;
      patterns[16832] = 25'b01000001_10111110_11111111_0;
      patterns[16833] = 25'b01000001_10111111_00000000_1;
      patterns[16834] = 25'b01000001_11000000_00000001_1;
      patterns[16835] = 25'b01000001_11000001_00000010_1;
      patterns[16836] = 25'b01000001_11000010_00000011_1;
      patterns[16837] = 25'b01000001_11000011_00000100_1;
      patterns[16838] = 25'b01000001_11000100_00000101_1;
      patterns[16839] = 25'b01000001_11000101_00000110_1;
      patterns[16840] = 25'b01000001_11000110_00000111_1;
      patterns[16841] = 25'b01000001_11000111_00001000_1;
      patterns[16842] = 25'b01000001_11001000_00001001_1;
      patterns[16843] = 25'b01000001_11001001_00001010_1;
      patterns[16844] = 25'b01000001_11001010_00001011_1;
      patterns[16845] = 25'b01000001_11001011_00001100_1;
      patterns[16846] = 25'b01000001_11001100_00001101_1;
      patterns[16847] = 25'b01000001_11001101_00001110_1;
      patterns[16848] = 25'b01000001_11001110_00001111_1;
      patterns[16849] = 25'b01000001_11001111_00010000_1;
      patterns[16850] = 25'b01000001_11010000_00010001_1;
      patterns[16851] = 25'b01000001_11010001_00010010_1;
      patterns[16852] = 25'b01000001_11010010_00010011_1;
      patterns[16853] = 25'b01000001_11010011_00010100_1;
      patterns[16854] = 25'b01000001_11010100_00010101_1;
      patterns[16855] = 25'b01000001_11010101_00010110_1;
      patterns[16856] = 25'b01000001_11010110_00010111_1;
      patterns[16857] = 25'b01000001_11010111_00011000_1;
      patterns[16858] = 25'b01000001_11011000_00011001_1;
      patterns[16859] = 25'b01000001_11011001_00011010_1;
      patterns[16860] = 25'b01000001_11011010_00011011_1;
      patterns[16861] = 25'b01000001_11011011_00011100_1;
      patterns[16862] = 25'b01000001_11011100_00011101_1;
      patterns[16863] = 25'b01000001_11011101_00011110_1;
      patterns[16864] = 25'b01000001_11011110_00011111_1;
      patterns[16865] = 25'b01000001_11011111_00100000_1;
      patterns[16866] = 25'b01000001_11100000_00100001_1;
      patterns[16867] = 25'b01000001_11100001_00100010_1;
      patterns[16868] = 25'b01000001_11100010_00100011_1;
      patterns[16869] = 25'b01000001_11100011_00100100_1;
      patterns[16870] = 25'b01000001_11100100_00100101_1;
      patterns[16871] = 25'b01000001_11100101_00100110_1;
      patterns[16872] = 25'b01000001_11100110_00100111_1;
      patterns[16873] = 25'b01000001_11100111_00101000_1;
      patterns[16874] = 25'b01000001_11101000_00101001_1;
      patterns[16875] = 25'b01000001_11101001_00101010_1;
      patterns[16876] = 25'b01000001_11101010_00101011_1;
      patterns[16877] = 25'b01000001_11101011_00101100_1;
      patterns[16878] = 25'b01000001_11101100_00101101_1;
      patterns[16879] = 25'b01000001_11101101_00101110_1;
      patterns[16880] = 25'b01000001_11101110_00101111_1;
      patterns[16881] = 25'b01000001_11101111_00110000_1;
      patterns[16882] = 25'b01000001_11110000_00110001_1;
      patterns[16883] = 25'b01000001_11110001_00110010_1;
      patterns[16884] = 25'b01000001_11110010_00110011_1;
      patterns[16885] = 25'b01000001_11110011_00110100_1;
      patterns[16886] = 25'b01000001_11110100_00110101_1;
      patterns[16887] = 25'b01000001_11110101_00110110_1;
      patterns[16888] = 25'b01000001_11110110_00110111_1;
      patterns[16889] = 25'b01000001_11110111_00111000_1;
      patterns[16890] = 25'b01000001_11111000_00111001_1;
      patterns[16891] = 25'b01000001_11111001_00111010_1;
      patterns[16892] = 25'b01000001_11111010_00111011_1;
      patterns[16893] = 25'b01000001_11111011_00111100_1;
      patterns[16894] = 25'b01000001_11111100_00111101_1;
      patterns[16895] = 25'b01000001_11111101_00111110_1;
      patterns[16896] = 25'b01000001_11111110_00111111_1;
      patterns[16897] = 25'b01000001_11111111_01000000_1;
      patterns[16898] = 25'b01000010_00000000_01000010_0;
      patterns[16899] = 25'b01000010_00000001_01000011_0;
      patterns[16900] = 25'b01000010_00000010_01000100_0;
      patterns[16901] = 25'b01000010_00000011_01000101_0;
      patterns[16902] = 25'b01000010_00000100_01000110_0;
      patterns[16903] = 25'b01000010_00000101_01000111_0;
      patterns[16904] = 25'b01000010_00000110_01001000_0;
      patterns[16905] = 25'b01000010_00000111_01001001_0;
      patterns[16906] = 25'b01000010_00001000_01001010_0;
      patterns[16907] = 25'b01000010_00001001_01001011_0;
      patterns[16908] = 25'b01000010_00001010_01001100_0;
      patterns[16909] = 25'b01000010_00001011_01001101_0;
      patterns[16910] = 25'b01000010_00001100_01001110_0;
      patterns[16911] = 25'b01000010_00001101_01001111_0;
      patterns[16912] = 25'b01000010_00001110_01010000_0;
      patterns[16913] = 25'b01000010_00001111_01010001_0;
      patterns[16914] = 25'b01000010_00010000_01010010_0;
      patterns[16915] = 25'b01000010_00010001_01010011_0;
      patterns[16916] = 25'b01000010_00010010_01010100_0;
      patterns[16917] = 25'b01000010_00010011_01010101_0;
      patterns[16918] = 25'b01000010_00010100_01010110_0;
      patterns[16919] = 25'b01000010_00010101_01010111_0;
      patterns[16920] = 25'b01000010_00010110_01011000_0;
      patterns[16921] = 25'b01000010_00010111_01011001_0;
      patterns[16922] = 25'b01000010_00011000_01011010_0;
      patterns[16923] = 25'b01000010_00011001_01011011_0;
      patterns[16924] = 25'b01000010_00011010_01011100_0;
      patterns[16925] = 25'b01000010_00011011_01011101_0;
      patterns[16926] = 25'b01000010_00011100_01011110_0;
      patterns[16927] = 25'b01000010_00011101_01011111_0;
      patterns[16928] = 25'b01000010_00011110_01100000_0;
      patterns[16929] = 25'b01000010_00011111_01100001_0;
      patterns[16930] = 25'b01000010_00100000_01100010_0;
      patterns[16931] = 25'b01000010_00100001_01100011_0;
      patterns[16932] = 25'b01000010_00100010_01100100_0;
      patterns[16933] = 25'b01000010_00100011_01100101_0;
      patterns[16934] = 25'b01000010_00100100_01100110_0;
      patterns[16935] = 25'b01000010_00100101_01100111_0;
      patterns[16936] = 25'b01000010_00100110_01101000_0;
      patterns[16937] = 25'b01000010_00100111_01101001_0;
      patterns[16938] = 25'b01000010_00101000_01101010_0;
      patterns[16939] = 25'b01000010_00101001_01101011_0;
      patterns[16940] = 25'b01000010_00101010_01101100_0;
      patterns[16941] = 25'b01000010_00101011_01101101_0;
      patterns[16942] = 25'b01000010_00101100_01101110_0;
      patterns[16943] = 25'b01000010_00101101_01101111_0;
      patterns[16944] = 25'b01000010_00101110_01110000_0;
      patterns[16945] = 25'b01000010_00101111_01110001_0;
      patterns[16946] = 25'b01000010_00110000_01110010_0;
      patterns[16947] = 25'b01000010_00110001_01110011_0;
      patterns[16948] = 25'b01000010_00110010_01110100_0;
      patterns[16949] = 25'b01000010_00110011_01110101_0;
      patterns[16950] = 25'b01000010_00110100_01110110_0;
      patterns[16951] = 25'b01000010_00110101_01110111_0;
      patterns[16952] = 25'b01000010_00110110_01111000_0;
      patterns[16953] = 25'b01000010_00110111_01111001_0;
      patterns[16954] = 25'b01000010_00111000_01111010_0;
      patterns[16955] = 25'b01000010_00111001_01111011_0;
      patterns[16956] = 25'b01000010_00111010_01111100_0;
      patterns[16957] = 25'b01000010_00111011_01111101_0;
      patterns[16958] = 25'b01000010_00111100_01111110_0;
      patterns[16959] = 25'b01000010_00111101_01111111_0;
      patterns[16960] = 25'b01000010_00111110_10000000_0;
      patterns[16961] = 25'b01000010_00111111_10000001_0;
      patterns[16962] = 25'b01000010_01000000_10000010_0;
      patterns[16963] = 25'b01000010_01000001_10000011_0;
      patterns[16964] = 25'b01000010_01000010_10000100_0;
      patterns[16965] = 25'b01000010_01000011_10000101_0;
      patterns[16966] = 25'b01000010_01000100_10000110_0;
      patterns[16967] = 25'b01000010_01000101_10000111_0;
      patterns[16968] = 25'b01000010_01000110_10001000_0;
      patterns[16969] = 25'b01000010_01000111_10001001_0;
      patterns[16970] = 25'b01000010_01001000_10001010_0;
      patterns[16971] = 25'b01000010_01001001_10001011_0;
      patterns[16972] = 25'b01000010_01001010_10001100_0;
      patterns[16973] = 25'b01000010_01001011_10001101_0;
      patterns[16974] = 25'b01000010_01001100_10001110_0;
      patterns[16975] = 25'b01000010_01001101_10001111_0;
      patterns[16976] = 25'b01000010_01001110_10010000_0;
      patterns[16977] = 25'b01000010_01001111_10010001_0;
      patterns[16978] = 25'b01000010_01010000_10010010_0;
      patterns[16979] = 25'b01000010_01010001_10010011_0;
      patterns[16980] = 25'b01000010_01010010_10010100_0;
      patterns[16981] = 25'b01000010_01010011_10010101_0;
      patterns[16982] = 25'b01000010_01010100_10010110_0;
      patterns[16983] = 25'b01000010_01010101_10010111_0;
      patterns[16984] = 25'b01000010_01010110_10011000_0;
      patterns[16985] = 25'b01000010_01010111_10011001_0;
      patterns[16986] = 25'b01000010_01011000_10011010_0;
      patterns[16987] = 25'b01000010_01011001_10011011_0;
      patterns[16988] = 25'b01000010_01011010_10011100_0;
      patterns[16989] = 25'b01000010_01011011_10011101_0;
      patterns[16990] = 25'b01000010_01011100_10011110_0;
      patterns[16991] = 25'b01000010_01011101_10011111_0;
      patterns[16992] = 25'b01000010_01011110_10100000_0;
      patterns[16993] = 25'b01000010_01011111_10100001_0;
      patterns[16994] = 25'b01000010_01100000_10100010_0;
      patterns[16995] = 25'b01000010_01100001_10100011_0;
      patterns[16996] = 25'b01000010_01100010_10100100_0;
      patterns[16997] = 25'b01000010_01100011_10100101_0;
      patterns[16998] = 25'b01000010_01100100_10100110_0;
      patterns[16999] = 25'b01000010_01100101_10100111_0;
      patterns[17000] = 25'b01000010_01100110_10101000_0;
      patterns[17001] = 25'b01000010_01100111_10101001_0;
      patterns[17002] = 25'b01000010_01101000_10101010_0;
      patterns[17003] = 25'b01000010_01101001_10101011_0;
      patterns[17004] = 25'b01000010_01101010_10101100_0;
      patterns[17005] = 25'b01000010_01101011_10101101_0;
      patterns[17006] = 25'b01000010_01101100_10101110_0;
      patterns[17007] = 25'b01000010_01101101_10101111_0;
      patterns[17008] = 25'b01000010_01101110_10110000_0;
      patterns[17009] = 25'b01000010_01101111_10110001_0;
      patterns[17010] = 25'b01000010_01110000_10110010_0;
      patterns[17011] = 25'b01000010_01110001_10110011_0;
      patterns[17012] = 25'b01000010_01110010_10110100_0;
      patterns[17013] = 25'b01000010_01110011_10110101_0;
      patterns[17014] = 25'b01000010_01110100_10110110_0;
      patterns[17015] = 25'b01000010_01110101_10110111_0;
      patterns[17016] = 25'b01000010_01110110_10111000_0;
      patterns[17017] = 25'b01000010_01110111_10111001_0;
      patterns[17018] = 25'b01000010_01111000_10111010_0;
      patterns[17019] = 25'b01000010_01111001_10111011_0;
      patterns[17020] = 25'b01000010_01111010_10111100_0;
      patterns[17021] = 25'b01000010_01111011_10111101_0;
      patterns[17022] = 25'b01000010_01111100_10111110_0;
      patterns[17023] = 25'b01000010_01111101_10111111_0;
      patterns[17024] = 25'b01000010_01111110_11000000_0;
      patterns[17025] = 25'b01000010_01111111_11000001_0;
      patterns[17026] = 25'b01000010_10000000_11000010_0;
      patterns[17027] = 25'b01000010_10000001_11000011_0;
      patterns[17028] = 25'b01000010_10000010_11000100_0;
      patterns[17029] = 25'b01000010_10000011_11000101_0;
      patterns[17030] = 25'b01000010_10000100_11000110_0;
      patterns[17031] = 25'b01000010_10000101_11000111_0;
      patterns[17032] = 25'b01000010_10000110_11001000_0;
      patterns[17033] = 25'b01000010_10000111_11001001_0;
      patterns[17034] = 25'b01000010_10001000_11001010_0;
      patterns[17035] = 25'b01000010_10001001_11001011_0;
      patterns[17036] = 25'b01000010_10001010_11001100_0;
      patterns[17037] = 25'b01000010_10001011_11001101_0;
      patterns[17038] = 25'b01000010_10001100_11001110_0;
      patterns[17039] = 25'b01000010_10001101_11001111_0;
      patterns[17040] = 25'b01000010_10001110_11010000_0;
      patterns[17041] = 25'b01000010_10001111_11010001_0;
      patterns[17042] = 25'b01000010_10010000_11010010_0;
      patterns[17043] = 25'b01000010_10010001_11010011_0;
      patterns[17044] = 25'b01000010_10010010_11010100_0;
      patterns[17045] = 25'b01000010_10010011_11010101_0;
      patterns[17046] = 25'b01000010_10010100_11010110_0;
      patterns[17047] = 25'b01000010_10010101_11010111_0;
      patterns[17048] = 25'b01000010_10010110_11011000_0;
      patterns[17049] = 25'b01000010_10010111_11011001_0;
      patterns[17050] = 25'b01000010_10011000_11011010_0;
      patterns[17051] = 25'b01000010_10011001_11011011_0;
      patterns[17052] = 25'b01000010_10011010_11011100_0;
      patterns[17053] = 25'b01000010_10011011_11011101_0;
      patterns[17054] = 25'b01000010_10011100_11011110_0;
      patterns[17055] = 25'b01000010_10011101_11011111_0;
      patterns[17056] = 25'b01000010_10011110_11100000_0;
      patterns[17057] = 25'b01000010_10011111_11100001_0;
      patterns[17058] = 25'b01000010_10100000_11100010_0;
      patterns[17059] = 25'b01000010_10100001_11100011_0;
      patterns[17060] = 25'b01000010_10100010_11100100_0;
      patterns[17061] = 25'b01000010_10100011_11100101_0;
      patterns[17062] = 25'b01000010_10100100_11100110_0;
      patterns[17063] = 25'b01000010_10100101_11100111_0;
      patterns[17064] = 25'b01000010_10100110_11101000_0;
      patterns[17065] = 25'b01000010_10100111_11101001_0;
      patterns[17066] = 25'b01000010_10101000_11101010_0;
      patterns[17067] = 25'b01000010_10101001_11101011_0;
      patterns[17068] = 25'b01000010_10101010_11101100_0;
      patterns[17069] = 25'b01000010_10101011_11101101_0;
      patterns[17070] = 25'b01000010_10101100_11101110_0;
      patterns[17071] = 25'b01000010_10101101_11101111_0;
      patterns[17072] = 25'b01000010_10101110_11110000_0;
      patterns[17073] = 25'b01000010_10101111_11110001_0;
      patterns[17074] = 25'b01000010_10110000_11110010_0;
      patterns[17075] = 25'b01000010_10110001_11110011_0;
      patterns[17076] = 25'b01000010_10110010_11110100_0;
      patterns[17077] = 25'b01000010_10110011_11110101_0;
      patterns[17078] = 25'b01000010_10110100_11110110_0;
      patterns[17079] = 25'b01000010_10110101_11110111_0;
      patterns[17080] = 25'b01000010_10110110_11111000_0;
      patterns[17081] = 25'b01000010_10110111_11111001_0;
      patterns[17082] = 25'b01000010_10111000_11111010_0;
      patterns[17083] = 25'b01000010_10111001_11111011_0;
      patterns[17084] = 25'b01000010_10111010_11111100_0;
      patterns[17085] = 25'b01000010_10111011_11111101_0;
      patterns[17086] = 25'b01000010_10111100_11111110_0;
      patterns[17087] = 25'b01000010_10111101_11111111_0;
      patterns[17088] = 25'b01000010_10111110_00000000_1;
      patterns[17089] = 25'b01000010_10111111_00000001_1;
      patterns[17090] = 25'b01000010_11000000_00000010_1;
      patterns[17091] = 25'b01000010_11000001_00000011_1;
      patterns[17092] = 25'b01000010_11000010_00000100_1;
      patterns[17093] = 25'b01000010_11000011_00000101_1;
      patterns[17094] = 25'b01000010_11000100_00000110_1;
      patterns[17095] = 25'b01000010_11000101_00000111_1;
      patterns[17096] = 25'b01000010_11000110_00001000_1;
      patterns[17097] = 25'b01000010_11000111_00001001_1;
      patterns[17098] = 25'b01000010_11001000_00001010_1;
      patterns[17099] = 25'b01000010_11001001_00001011_1;
      patterns[17100] = 25'b01000010_11001010_00001100_1;
      patterns[17101] = 25'b01000010_11001011_00001101_1;
      patterns[17102] = 25'b01000010_11001100_00001110_1;
      patterns[17103] = 25'b01000010_11001101_00001111_1;
      patterns[17104] = 25'b01000010_11001110_00010000_1;
      patterns[17105] = 25'b01000010_11001111_00010001_1;
      patterns[17106] = 25'b01000010_11010000_00010010_1;
      patterns[17107] = 25'b01000010_11010001_00010011_1;
      patterns[17108] = 25'b01000010_11010010_00010100_1;
      patterns[17109] = 25'b01000010_11010011_00010101_1;
      patterns[17110] = 25'b01000010_11010100_00010110_1;
      patterns[17111] = 25'b01000010_11010101_00010111_1;
      patterns[17112] = 25'b01000010_11010110_00011000_1;
      patterns[17113] = 25'b01000010_11010111_00011001_1;
      patterns[17114] = 25'b01000010_11011000_00011010_1;
      patterns[17115] = 25'b01000010_11011001_00011011_1;
      patterns[17116] = 25'b01000010_11011010_00011100_1;
      patterns[17117] = 25'b01000010_11011011_00011101_1;
      patterns[17118] = 25'b01000010_11011100_00011110_1;
      patterns[17119] = 25'b01000010_11011101_00011111_1;
      patterns[17120] = 25'b01000010_11011110_00100000_1;
      patterns[17121] = 25'b01000010_11011111_00100001_1;
      patterns[17122] = 25'b01000010_11100000_00100010_1;
      patterns[17123] = 25'b01000010_11100001_00100011_1;
      patterns[17124] = 25'b01000010_11100010_00100100_1;
      patterns[17125] = 25'b01000010_11100011_00100101_1;
      patterns[17126] = 25'b01000010_11100100_00100110_1;
      patterns[17127] = 25'b01000010_11100101_00100111_1;
      patterns[17128] = 25'b01000010_11100110_00101000_1;
      patterns[17129] = 25'b01000010_11100111_00101001_1;
      patterns[17130] = 25'b01000010_11101000_00101010_1;
      patterns[17131] = 25'b01000010_11101001_00101011_1;
      patterns[17132] = 25'b01000010_11101010_00101100_1;
      patterns[17133] = 25'b01000010_11101011_00101101_1;
      patterns[17134] = 25'b01000010_11101100_00101110_1;
      patterns[17135] = 25'b01000010_11101101_00101111_1;
      patterns[17136] = 25'b01000010_11101110_00110000_1;
      patterns[17137] = 25'b01000010_11101111_00110001_1;
      patterns[17138] = 25'b01000010_11110000_00110010_1;
      patterns[17139] = 25'b01000010_11110001_00110011_1;
      patterns[17140] = 25'b01000010_11110010_00110100_1;
      patterns[17141] = 25'b01000010_11110011_00110101_1;
      patterns[17142] = 25'b01000010_11110100_00110110_1;
      patterns[17143] = 25'b01000010_11110101_00110111_1;
      patterns[17144] = 25'b01000010_11110110_00111000_1;
      patterns[17145] = 25'b01000010_11110111_00111001_1;
      patterns[17146] = 25'b01000010_11111000_00111010_1;
      patterns[17147] = 25'b01000010_11111001_00111011_1;
      patterns[17148] = 25'b01000010_11111010_00111100_1;
      patterns[17149] = 25'b01000010_11111011_00111101_1;
      patterns[17150] = 25'b01000010_11111100_00111110_1;
      patterns[17151] = 25'b01000010_11111101_00111111_1;
      patterns[17152] = 25'b01000010_11111110_01000000_1;
      patterns[17153] = 25'b01000010_11111111_01000001_1;
      patterns[17154] = 25'b01000011_00000000_01000011_0;
      patterns[17155] = 25'b01000011_00000001_01000100_0;
      patterns[17156] = 25'b01000011_00000010_01000101_0;
      patterns[17157] = 25'b01000011_00000011_01000110_0;
      patterns[17158] = 25'b01000011_00000100_01000111_0;
      patterns[17159] = 25'b01000011_00000101_01001000_0;
      patterns[17160] = 25'b01000011_00000110_01001001_0;
      patterns[17161] = 25'b01000011_00000111_01001010_0;
      patterns[17162] = 25'b01000011_00001000_01001011_0;
      patterns[17163] = 25'b01000011_00001001_01001100_0;
      patterns[17164] = 25'b01000011_00001010_01001101_0;
      patterns[17165] = 25'b01000011_00001011_01001110_0;
      patterns[17166] = 25'b01000011_00001100_01001111_0;
      patterns[17167] = 25'b01000011_00001101_01010000_0;
      patterns[17168] = 25'b01000011_00001110_01010001_0;
      patterns[17169] = 25'b01000011_00001111_01010010_0;
      patterns[17170] = 25'b01000011_00010000_01010011_0;
      patterns[17171] = 25'b01000011_00010001_01010100_0;
      patterns[17172] = 25'b01000011_00010010_01010101_0;
      patterns[17173] = 25'b01000011_00010011_01010110_0;
      patterns[17174] = 25'b01000011_00010100_01010111_0;
      patterns[17175] = 25'b01000011_00010101_01011000_0;
      patterns[17176] = 25'b01000011_00010110_01011001_0;
      patterns[17177] = 25'b01000011_00010111_01011010_0;
      patterns[17178] = 25'b01000011_00011000_01011011_0;
      patterns[17179] = 25'b01000011_00011001_01011100_0;
      patterns[17180] = 25'b01000011_00011010_01011101_0;
      patterns[17181] = 25'b01000011_00011011_01011110_0;
      patterns[17182] = 25'b01000011_00011100_01011111_0;
      patterns[17183] = 25'b01000011_00011101_01100000_0;
      patterns[17184] = 25'b01000011_00011110_01100001_0;
      patterns[17185] = 25'b01000011_00011111_01100010_0;
      patterns[17186] = 25'b01000011_00100000_01100011_0;
      patterns[17187] = 25'b01000011_00100001_01100100_0;
      patterns[17188] = 25'b01000011_00100010_01100101_0;
      patterns[17189] = 25'b01000011_00100011_01100110_0;
      patterns[17190] = 25'b01000011_00100100_01100111_0;
      patterns[17191] = 25'b01000011_00100101_01101000_0;
      patterns[17192] = 25'b01000011_00100110_01101001_0;
      patterns[17193] = 25'b01000011_00100111_01101010_0;
      patterns[17194] = 25'b01000011_00101000_01101011_0;
      patterns[17195] = 25'b01000011_00101001_01101100_0;
      patterns[17196] = 25'b01000011_00101010_01101101_0;
      patterns[17197] = 25'b01000011_00101011_01101110_0;
      patterns[17198] = 25'b01000011_00101100_01101111_0;
      patterns[17199] = 25'b01000011_00101101_01110000_0;
      patterns[17200] = 25'b01000011_00101110_01110001_0;
      patterns[17201] = 25'b01000011_00101111_01110010_0;
      patterns[17202] = 25'b01000011_00110000_01110011_0;
      patterns[17203] = 25'b01000011_00110001_01110100_0;
      patterns[17204] = 25'b01000011_00110010_01110101_0;
      patterns[17205] = 25'b01000011_00110011_01110110_0;
      patterns[17206] = 25'b01000011_00110100_01110111_0;
      patterns[17207] = 25'b01000011_00110101_01111000_0;
      patterns[17208] = 25'b01000011_00110110_01111001_0;
      patterns[17209] = 25'b01000011_00110111_01111010_0;
      patterns[17210] = 25'b01000011_00111000_01111011_0;
      patterns[17211] = 25'b01000011_00111001_01111100_0;
      patterns[17212] = 25'b01000011_00111010_01111101_0;
      patterns[17213] = 25'b01000011_00111011_01111110_0;
      patterns[17214] = 25'b01000011_00111100_01111111_0;
      patterns[17215] = 25'b01000011_00111101_10000000_0;
      patterns[17216] = 25'b01000011_00111110_10000001_0;
      patterns[17217] = 25'b01000011_00111111_10000010_0;
      patterns[17218] = 25'b01000011_01000000_10000011_0;
      patterns[17219] = 25'b01000011_01000001_10000100_0;
      patterns[17220] = 25'b01000011_01000010_10000101_0;
      patterns[17221] = 25'b01000011_01000011_10000110_0;
      patterns[17222] = 25'b01000011_01000100_10000111_0;
      patterns[17223] = 25'b01000011_01000101_10001000_0;
      patterns[17224] = 25'b01000011_01000110_10001001_0;
      patterns[17225] = 25'b01000011_01000111_10001010_0;
      patterns[17226] = 25'b01000011_01001000_10001011_0;
      patterns[17227] = 25'b01000011_01001001_10001100_0;
      patterns[17228] = 25'b01000011_01001010_10001101_0;
      patterns[17229] = 25'b01000011_01001011_10001110_0;
      patterns[17230] = 25'b01000011_01001100_10001111_0;
      patterns[17231] = 25'b01000011_01001101_10010000_0;
      patterns[17232] = 25'b01000011_01001110_10010001_0;
      patterns[17233] = 25'b01000011_01001111_10010010_0;
      patterns[17234] = 25'b01000011_01010000_10010011_0;
      patterns[17235] = 25'b01000011_01010001_10010100_0;
      patterns[17236] = 25'b01000011_01010010_10010101_0;
      patterns[17237] = 25'b01000011_01010011_10010110_0;
      patterns[17238] = 25'b01000011_01010100_10010111_0;
      patterns[17239] = 25'b01000011_01010101_10011000_0;
      patterns[17240] = 25'b01000011_01010110_10011001_0;
      patterns[17241] = 25'b01000011_01010111_10011010_0;
      patterns[17242] = 25'b01000011_01011000_10011011_0;
      patterns[17243] = 25'b01000011_01011001_10011100_0;
      patterns[17244] = 25'b01000011_01011010_10011101_0;
      patterns[17245] = 25'b01000011_01011011_10011110_0;
      patterns[17246] = 25'b01000011_01011100_10011111_0;
      patterns[17247] = 25'b01000011_01011101_10100000_0;
      patterns[17248] = 25'b01000011_01011110_10100001_0;
      patterns[17249] = 25'b01000011_01011111_10100010_0;
      patterns[17250] = 25'b01000011_01100000_10100011_0;
      patterns[17251] = 25'b01000011_01100001_10100100_0;
      patterns[17252] = 25'b01000011_01100010_10100101_0;
      patterns[17253] = 25'b01000011_01100011_10100110_0;
      patterns[17254] = 25'b01000011_01100100_10100111_0;
      patterns[17255] = 25'b01000011_01100101_10101000_0;
      patterns[17256] = 25'b01000011_01100110_10101001_0;
      patterns[17257] = 25'b01000011_01100111_10101010_0;
      patterns[17258] = 25'b01000011_01101000_10101011_0;
      patterns[17259] = 25'b01000011_01101001_10101100_0;
      patterns[17260] = 25'b01000011_01101010_10101101_0;
      patterns[17261] = 25'b01000011_01101011_10101110_0;
      patterns[17262] = 25'b01000011_01101100_10101111_0;
      patterns[17263] = 25'b01000011_01101101_10110000_0;
      patterns[17264] = 25'b01000011_01101110_10110001_0;
      patterns[17265] = 25'b01000011_01101111_10110010_0;
      patterns[17266] = 25'b01000011_01110000_10110011_0;
      patterns[17267] = 25'b01000011_01110001_10110100_0;
      patterns[17268] = 25'b01000011_01110010_10110101_0;
      patterns[17269] = 25'b01000011_01110011_10110110_0;
      patterns[17270] = 25'b01000011_01110100_10110111_0;
      patterns[17271] = 25'b01000011_01110101_10111000_0;
      patterns[17272] = 25'b01000011_01110110_10111001_0;
      patterns[17273] = 25'b01000011_01110111_10111010_0;
      patterns[17274] = 25'b01000011_01111000_10111011_0;
      patterns[17275] = 25'b01000011_01111001_10111100_0;
      patterns[17276] = 25'b01000011_01111010_10111101_0;
      patterns[17277] = 25'b01000011_01111011_10111110_0;
      patterns[17278] = 25'b01000011_01111100_10111111_0;
      patterns[17279] = 25'b01000011_01111101_11000000_0;
      patterns[17280] = 25'b01000011_01111110_11000001_0;
      patterns[17281] = 25'b01000011_01111111_11000010_0;
      patterns[17282] = 25'b01000011_10000000_11000011_0;
      patterns[17283] = 25'b01000011_10000001_11000100_0;
      patterns[17284] = 25'b01000011_10000010_11000101_0;
      patterns[17285] = 25'b01000011_10000011_11000110_0;
      patterns[17286] = 25'b01000011_10000100_11000111_0;
      patterns[17287] = 25'b01000011_10000101_11001000_0;
      patterns[17288] = 25'b01000011_10000110_11001001_0;
      patterns[17289] = 25'b01000011_10000111_11001010_0;
      patterns[17290] = 25'b01000011_10001000_11001011_0;
      patterns[17291] = 25'b01000011_10001001_11001100_0;
      patterns[17292] = 25'b01000011_10001010_11001101_0;
      patterns[17293] = 25'b01000011_10001011_11001110_0;
      patterns[17294] = 25'b01000011_10001100_11001111_0;
      patterns[17295] = 25'b01000011_10001101_11010000_0;
      patterns[17296] = 25'b01000011_10001110_11010001_0;
      patterns[17297] = 25'b01000011_10001111_11010010_0;
      patterns[17298] = 25'b01000011_10010000_11010011_0;
      patterns[17299] = 25'b01000011_10010001_11010100_0;
      patterns[17300] = 25'b01000011_10010010_11010101_0;
      patterns[17301] = 25'b01000011_10010011_11010110_0;
      patterns[17302] = 25'b01000011_10010100_11010111_0;
      patterns[17303] = 25'b01000011_10010101_11011000_0;
      patterns[17304] = 25'b01000011_10010110_11011001_0;
      patterns[17305] = 25'b01000011_10010111_11011010_0;
      patterns[17306] = 25'b01000011_10011000_11011011_0;
      patterns[17307] = 25'b01000011_10011001_11011100_0;
      patterns[17308] = 25'b01000011_10011010_11011101_0;
      patterns[17309] = 25'b01000011_10011011_11011110_0;
      patterns[17310] = 25'b01000011_10011100_11011111_0;
      patterns[17311] = 25'b01000011_10011101_11100000_0;
      patterns[17312] = 25'b01000011_10011110_11100001_0;
      patterns[17313] = 25'b01000011_10011111_11100010_0;
      patterns[17314] = 25'b01000011_10100000_11100011_0;
      patterns[17315] = 25'b01000011_10100001_11100100_0;
      patterns[17316] = 25'b01000011_10100010_11100101_0;
      patterns[17317] = 25'b01000011_10100011_11100110_0;
      patterns[17318] = 25'b01000011_10100100_11100111_0;
      patterns[17319] = 25'b01000011_10100101_11101000_0;
      patterns[17320] = 25'b01000011_10100110_11101001_0;
      patterns[17321] = 25'b01000011_10100111_11101010_0;
      patterns[17322] = 25'b01000011_10101000_11101011_0;
      patterns[17323] = 25'b01000011_10101001_11101100_0;
      patterns[17324] = 25'b01000011_10101010_11101101_0;
      patterns[17325] = 25'b01000011_10101011_11101110_0;
      patterns[17326] = 25'b01000011_10101100_11101111_0;
      patterns[17327] = 25'b01000011_10101101_11110000_0;
      patterns[17328] = 25'b01000011_10101110_11110001_0;
      patterns[17329] = 25'b01000011_10101111_11110010_0;
      patterns[17330] = 25'b01000011_10110000_11110011_0;
      patterns[17331] = 25'b01000011_10110001_11110100_0;
      patterns[17332] = 25'b01000011_10110010_11110101_0;
      patterns[17333] = 25'b01000011_10110011_11110110_0;
      patterns[17334] = 25'b01000011_10110100_11110111_0;
      patterns[17335] = 25'b01000011_10110101_11111000_0;
      patterns[17336] = 25'b01000011_10110110_11111001_0;
      patterns[17337] = 25'b01000011_10110111_11111010_0;
      patterns[17338] = 25'b01000011_10111000_11111011_0;
      patterns[17339] = 25'b01000011_10111001_11111100_0;
      patterns[17340] = 25'b01000011_10111010_11111101_0;
      patterns[17341] = 25'b01000011_10111011_11111110_0;
      patterns[17342] = 25'b01000011_10111100_11111111_0;
      patterns[17343] = 25'b01000011_10111101_00000000_1;
      patterns[17344] = 25'b01000011_10111110_00000001_1;
      patterns[17345] = 25'b01000011_10111111_00000010_1;
      patterns[17346] = 25'b01000011_11000000_00000011_1;
      patterns[17347] = 25'b01000011_11000001_00000100_1;
      patterns[17348] = 25'b01000011_11000010_00000101_1;
      patterns[17349] = 25'b01000011_11000011_00000110_1;
      patterns[17350] = 25'b01000011_11000100_00000111_1;
      patterns[17351] = 25'b01000011_11000101_00001000_1;
      patterns[17352] = 25'b01000011_11000110_00001001_1;
      patterns[17353] = 25'b01000011_11000111_00001010_1;
      patterns[17354] = 25'b01000011_11001000_00001011_1;
      patterns[17355] = 25'b01000011_11001001_00001100_1;
      patterns[17356] = 25'b01000011_11001010_00001101_1;
      patterns[17357] = 25'b01000011_11001011_00001110_1;
      patterns[17358] = 25'b01000011_11001100_00001111_1;
      patterns[17359] = 25'b01000011_11001101_00010000_1;
      patterns[17360] = 25'b01000011_11001110_00010001_1;
      patterns[17361] = 25'b01000011_11001111_00010010_1;
      patterns[17362] = 25'b01000011_11010000_00010011_1;
      patterns[17363] = 25'b01000011_11010001_00010100_1;
      patterns[17364] = 25'b01000011_11010010_00010101_1;
      patterns[17365] = 25'b01000011_11010011_00010110_1;
      patterns[17366] = 25'b01000011_11010100_00010111_1;
      patterns[17367] = 25'b01000011_11010101_00011000_1;
      patterns[17368] = 25'b01000011_11010110_00011001_1;
      patterns[17369] = 25'b01000011_11010111_00011010_1;
      patterns[17370] = 25'b01000011_11011000_00011011_1;
      patterns[17371] = 25'b01000011_11011001_00011100_1;
      patterns[17372] = 25'b01000011_11011010_00011101_1;
      patterns[17373] = 25'b01000011_11011011_00011110_1;
      patterns[17374] = 25'b01000011_11011100_00011111_1;
      patterns[17375] = 25'b01000011_11011101_00100000_1;
      patterns[17376] = 25'b01000011_11011110_00100001_1;
      patterns[17377] = 25'b01000011_11011111_00100010_1;
      patterns[17378] = 25'b01000011_11100000_00100011_1;
      patterns[17379] = 25'b01000011_11100001_00100100_1;
      patterns[17380] = 25'b01000011_11100010_00100101_1;
      patterns[17381] = 25'b01000011_11100011_00100110_1;
      patterns[17382] = 25'b01000011_11100100_00100111_1;
      patterns[17383] = 25'b01000011_11100101_00101000_1;
      patterns[17384] = 25'b01000011_11100110_00101001_1;
      patterns[17385] = 25'b01000011_11100111_00101010_1;
      patterns[17386] = 25'b01000011_11101000_00101011_1;
      patterns[17387] = 25'b01000011_11101001_00101100_1;
      patterns[17388] = 25'b01000011_11101010_00101101_1;
      patterns[17389] = 25'b01000011_11101011_00101110_1;
      patterns[17390] = 25'b01000011_11101100_00101111_1;
      patterns[17391] = 25'b01000011_11101101_00110000_1;
      patterns[17392] = 25'b01000011_11101110_00110001_1;
      patterns[17393] = 25'b01000011_11101111_00110010_1;
      patterns[17394] = 25'b01000011_11110000_00110011_1;
      patterns[17395] = 25'b01000011_11110001_00110100_1;
      patterns[17396] = 25'b01000011_11110010_00110101_1;
      patterns[17397] = 25'b01000011_11110011_00110110_1;
      patterns[17398] = 25'b01000011_11110100_00110111_1;
      patterns[17399] = 25'b01000011_11110101_00111000_1;
      patterns[17400] = 25'b01000011_11110110_00111001_1;
      patterns[17401] = 25'b01000011_11110111_00111010_1;
      patterns[17402] = 25'b01000011_11111000_00111011_1;
      patterns[17403] = 25'b01000011_11111001_00111100_1;
      patterns[17404] = 25'b01000011_11111010_00111101_1;
      patterns[17405] = 25'b01000011_11111011_00111110_1;
      patterns[17406] = 25'b01000011_11111100_00111111_1;
      patterns[17407] = 25'b01000011_11111101_01000000_1;
      patterns[17408] = 25'b01000011_11111110_01000001_1;
      patterns[17409] = 25'b01000011_11111111_01000010_1;
      patterns[17410] = 25'b01000100_00000000_01000100_0;
      patterns[17411] = 25'b01000100_00000001_01000101_0;
      patterns[17412] = 25'b01000100_00000010_01000110_0;
      patterns[17413] = 25'b01000100_00000011_01000111_0;
      patterns[17414] = 25'b01000100_00000100_01001000_0;
      patterns[17415] = 25'b01000100_00000101_01001001_0;
      patterns[17416] = 25'b01000100_00000110_01001010_0;
      patterns[17417] = 25'b01000100_00000111_01001011_0;
      patterns[17418] = 25'b01000100_00001000_01001100_0;
      patterns[17419] = 25'b01000100_00001001_01001101_0;
      patterns[17420] = 25'b01000100_00001010_01001110_0;
      patterns[17421] = 25'b01000100_00001011_01001111_0;
      patterns[17422] = 25'b01000100_00001100_01010000_0;
      patterns[17423] = 25'b01000100_00001101_01010001_0;
      patterns[17424] = 25'b01000100_00001110_01010010_0;
      patterns[17425] = 25'b01000100_00001111_01010011_0;
      patterns[17426] = 25'b01000100_00010000_01010100_0;
      patterns[17427] = 25'b01000100_00010001_01010101_0;
      patterns[17428] = 25'b01000100_00010010_01010110_0;
      patterns[17429] = 25'b01000100_00010011_01010111_0;
      patterns[17430] = 25'b01000100_00010100_01011000_0;
      patterns[17431] = 25'b01000100_00010101_01011001_0;
      patterns[17432] = 25'b01000100_00010110_01011010_0;
      patterns[17433] = 25'b01000100_00010111_01011011_0;
      patterns[17434] = 25'b01000100_00011000_01011100_0;
      patterns[17435] = 25'b01000100_00011001_01011101_0;
      patterns[17436] = 25'b01000100_00011010_01011110_0;
      patterns[17437] = 25'b01000100_00011011_01011111_0;
      patterns[17438] = 25'b01000100_00011100_01100000_0;
      patterns[17439] = 25'b01000100_00011101_01100001_0;
      patterns[17440] = 25'b01000100_00011110_01100010_0;
      patterns[17441] = 25'b01000100_00011111_01100011_0;
      patterns[17442] = 25'b01000100_00100000_01100100_0;
      patterns[17443] = 25'b01000100_00100001_01100101_0;
      patterns[17444] = 25'b01000100_00100010_01100110_0;
      patterns[17445] = 25'b01000100_00100011_01100111_0;
      patterns[17446] = 25'b01000100_00100100_01101000_0;
      patterns[17447] = 25'b01000100_00100101_01101001_0;
      patterns[17448] = 25'b01000100_00100110_01101010_0;
      patterns[17449] = 25'b01000100_00100111_01101011_0;
      patterns[17450] = 25'b01000100_00101000_01101100_0;
      patterns[17451] = 25'b01000100_00101001_01101101_0;
      patterns[17452] = 25'b01000100_00101010_01101110_0;
      patterns[17453] = 25'b01000100_00101011_01101111_0;
      patterns[17454] = 25'b01000100_00101100_01110000_0;
      patterns[17455] = 25'b01000100_00101101_01110001_0;
      patterns[17456] = 25'b01000100_00101110_01110010_0;
      patterns[17457] = 25'b01000100_00101111_01110011_0;
      patterns[17458] = 25'b01000100_00110000_01110100_0;
      patterns[17459] = 25'b01000100_00110001_01110101_0;
      patterns[17460] = 25'b01000100_00110010_01110110_0;
      patterns[17461] = 25'b01000100_00110011_01110111_0;
      patterns[17462] = 25'b01000100_00110100_01111000_0;
      patterns[17463] = 25'b01000100_00110101_01111001_0;
      patterns[17464] = 25'b01000100_00110110_01111010_0;
      patterns[17465] = 25'b01000100_00110111_01111011_0;
      patterns[17466] = 25'b01000100_00111000_01111100_0;
      patterns[17467] = 25'b01000100_00111001_01111101_0;
      patterns[17468] = 25'b01000100_00111010_01111110_0;
      patterns[17469] = 25'b01000100_00111011_01111111_0;
      patterns[17470] = 25'b01000100_00111100_10000000_0;
      patterns[17471] = 25'b01000100_00111101_10000001_0;
      patterns[17472] = 25'b01000100_00111110_10000010_0;
      patterns[17473] = 25'b01000100_00111111_10000011_0;
      patterns[17474] = 25'b01000100_01000000_10000100_0;
      patterns[17475] = 25'b01000100_01000001_10000101_0;
      patterns[17476] = 25'b01000100_01000010_10000110_0;
      patterns[17477] = 25'b01000100_01000011_10000111_0;
      patterns[17478] = 25'b01000100_01000100_10001000_0;
      patterns[17479] = 25'b01000100_01000101_10001001_0;
      patterns[17480] = 25'b01000100_01000110_10001010_0;
      patterns[17481] = 25'b01000100_01000111_10001011_0;
      patterns[17482] = 25'b01000100_01001000_10001100_0;
      patterns[17483] = 25'b01000100_01001001_10001101_0;
      patterns[17484] = 25'b01000100_01001010_10001110_0;
      patterns[17485] = 25'b01000100_01001011_10001111_0;
      patterns[17486] = 25'b01000100_01001100_10010000_0;
      patterns[17487] = 25'b01000100_01001101_10010001_0;
      patterns[17488] = 25'b01000100_01001110_10010010_0;
      patterns[17489] = 25'b01000100_01001111_10010011_0;
      patterns[17490] = 25'b01000100_01010000_10010100_0;
      patterns[17491] = 25'b01000100_01010001_10010101_0;
      patterns[17492] = 25'b01000100_01010010_10010110_0;
      patterns[17493] = 25'b01000100_01010011_10010111_0;
      patterns[17494] = 25'b01000100_01010100_10011000_0;
      patterns[17495] = 25'b01000100_01010101_10011001_0;
      patterns[17496] = 25'b01000100_01010110_10011010_0;
      patterns[17497] = 25'b01000100_01010111_10011011_0;
      patterns[17498] = 25'b01000100_01011000_10011100_0;
      patterns[17499] = 25'b01000100_01011001_10011101_0;
      patterns[17500] = 25'b01000100_01011010_10011110_0;
      patterns[17501] = 25'b01000100_01011011_10011111_0;
      patterns[17502] = 25'b01000100_01011100_10100000_0;
      patterns[17503] = 25'b01000100_01011101_10100001_0;
      patterns[17504] = 25'b01000100_01011110_10100010_0;
      patterns[17505] = 25'b01000100_01011111_10100011_0;
      patterns[17506] = 25'b01000100_01100000_10100100_0;
      patterns[17507] = 25'b01000100_01100001_10100101_0;
      patterns[17508] = 25'b01000100_01100010_10100110_0;
      patterns[17509] = 25'b01000100_01100011_10100111_0;
      patterns[17510] = 25'b01000100_01100100_10101000_0;
      patterns[17511] = 25'b01000100_01100101_10101001_0;
      patterns[17512] = 25'b01000100_01100110_10101010_0;
      patterns[17513] = 25'b01000100_01100111_10101011_0;
      patterns[17514] = 25'b01000100_01101000_10101100_0;
      patterns[17515] = 25'b01000100_01101001_10101101_0;
      patterns[17516] = 25'b01000100_01101010_10101110_0;
      patterns[17517] = 25'b01000100_01101011_10101111_0;
      patterns[17518] = 25'b01000100_01101100_10110000_0;
      patterns[17519] = 25'b01000100_01101101_10110001_0;
      patterns[17520] = 25'b01000100_01101110_10110010_0;
      patterns[17521] = 25'b01000100_01101111_10110011_0;
      patterns[17522] = 25'b01000100_01110000_10110100_0;
      patterns[17523] = 25'b01000100_01110001_10110101_0;
      patterns[17524] = 25'b01000100_01110010_10110110_0;
      patterns[17525] = 25'b01000100_01110011_10110111_0;
      patterns[17526] = 25'b01000100_01110100_10111000_0;
      patterns[17527] = 25'b01000100_01110101_10111001_0;
      patterns[17528] = 25'b01000100_01110110_10111010_0;
      patterns[17529] = 25'b01000100_01110111_10111011_0;
      patterns[17530] = 25'b01000100_01111000_10111100_0;
      patterns[17531] = 25'b01000100_01111001_10111101_0;
      patterns[17532] = 25'b01000100_01111010_10111110_0;
      patterns[17533] = 25'b01000100_01111011_10111111_0;
      patterns[17534] = 25'b01000100_01111100_11000000_0;
      patterns[17535] = 25'b01000100_01111101_11000001_0;
      patterns[17536] = 25'b01000100_01111110_11000010_0;
      patterns[17537] = 25'b01000100_01111111_11000011_0;
      patterns[17538] = 25'b01000100_10000000_11000100_0;
      patterns[17539] = 25'b01000100_10000001_11000101_0;
      patterns[17540] = 25'b01000100_10000010_11000110_0;
      patterns[17541] = 25'b01000100_10000011_11000111_0;
      patterns[17542] = 25'b01000100_10000100_11001000_0;
      patterns[17543] = 25'b01000100_10000101_11001001_0;
      patterns[17544] = 25'b01000100_10000110_11001010_0;
      patterns[17545] = 25'b01000100_10000111_11001011_0;
      patterns[17546] = 25'b01000100_10001000_11001100_0;
      patterns[17547] = 25'b01000100_10001001_11001101_0;
      patterns[17548] = 25'b01000100_10001010_11001110_0;
      patterns[17549] = 25'b01000100_10001011_11001111_0;
      patterns[17550] = 25'b01000100_10001100_11010000_0;
      patterns[17551] = 25'b01000100_10001101_11010001_0;
      patterns[17552] = 25'b01000100_10001110_11010010_0;
      patterns[17553] = 25'b01000100_10001111_11010011_0;
      patterns[17554] = 25'b01000100_10010000_11010100_0;
      patterns[17555] = 25'b01000100_10010001_11010101_0;
      patterns[17556] = 25'b01000100_10010010_11010110_0;
      patterns[17557] = 25'b01000100_10010011_11010111_0;
      patterns[17558] = 25'b01000100_10010100_11011000_0;
      patterns[17559] = 25'b01000100_10010101_11011001_0;
      patterns[17560] = 25'b01000100_10010110_11011010_0;
      patterns[17561] = 25'b01000100_10010111_11011011_0;
      patterns[17562] = 25'b01000100_10011000_11011100_0;
      patterns[17563] = 25'b01000100_10011001_11011101_0;
      patterns[17564] = 25'b01000100_10011010_11011110_0;
      patterns[17565] = 25'b01000100_10011011_11011111_0;
      patterns[17566] = 25'b01000100_10011100_11100000_0;
      patterns[17567] = 25'b01000100_10011101_11100001_0;
      patterns[17568] = 25'b01000100_10011110_11100010_0;
      patterns[17569] = 25'b01000100_10011111_11100011_0;
      patterns[17570] = 25'b01000100_10100000_11100100_0;
      patterns[17571] = 25'b01000100_10100001_11100101_0;
      patterns[17572] = 25'b01000100_10100010_11100110_0;
      patterns[17573] = 25'b01000100_10100011_11100111_0;
      patterns[17574] = 25'b01000100_10100100_11101000_0;
      patterns[17575] = 25'b01000100_10100101_11101001_0;
      patterns[17576] = 25'b01000100_10100110_11101010_0;
      patterns[17577] = 25'b01000100_10100111_11101011_0;
      patterns[17578] = 25'b01000100_10101000_11101100_0;
      patterns[17579] = 25'b01000100_10101001_11101101_0;
      patterns[17580] = 25'b01000100_10101010_11101110_0;
      patterns[17581] = 25'b01000100_10101011_11101111_0;
      patterns[17582] = 25'b01000100_10101100_11110000_0;
      patterns[17583] = 25'b01000100_10101101_11110001_0;
      patterns[17584] = 25'b01000100_10101110_11110010_0;
      patterns[17585] = 25'b01000100_10101111_11110011_0;
      patterns[17586] = 25'b01000100_10110000_11110100_0;
      patterns[17587] = 25'b01000100_10110001_11110101_0;
      patterns[17588] = 25'b01000100_10110010_11110110_0;
      patterns[17589] = 25'b01000100_10110011_11110111_0;
      patterns[17590] = 25'b01000100_10110100_11111000_0;
      patterns[17591] = 25'b01000100_10110101_11111001_0;
      patterns[17592] = 25'b01000100_10110110_11111010_0;
      patterns[17593] = 25'b01000100_10110111_11111011_0;
      patterns[17594] = 25'b01000100_10111000_11111100_0;
      patterns[17595] = 25'b01000100_10111001_11111101_0;
      patterns[17596] = 25'b01000100_10111010_11111110_0;
      patterns[17597] = 25'b01000100_10111011_11111111_0;
      patterns[17598] = 25'b01000100_10111100_00000000_1;
      patterns[17599] = 25'b01000100_10111101_00000001_1;
      patterns[17600] = 25'b01000100_10111110_00000010_1;
      patterns[17601] = 25'b01000100_10111111_00000011_1;
      patterns[17602] = 25'b01000100_11000000_00000100_1;
      patterns[17603] = 25'b01000100_11000001_00000101_1;
      patterns[17604] = 25'b01000100_11000010_00000110_1;
      patterns[17605] = 25'b01000100_11000011_00000111_1;
      patterns[17606] = 25'b01000100_11000100_00001000_1;
      patterns[17607] = 25'b01000100_11000101_00001001_1;
      patterns[17608] = 25'b01000100_11000110_00001010_1;
      patterns[17609] = 25'b01000100_11000111_00001011_1;
      patterns[17610] = 25'b01000100_11001000_00001100_1;
      patterns[17611] = 25'b01000100_11001001_00001101_1;
      patterns[17612] = 25'b01000100_11001010_00001110_1;
      patterns[17613] = 25'b01000100_11001011_00001111_1;
      patterns[17614] = 25'b01000100_11001100_00010000_1;
      patterns[17615] = 25'b01000100_11001101_00010001_1;
      patterns[17616] = 25'b01000100_11001110_00010010_1;
      patterns[17617] = 25'b01000100_11001111_00010011_1;
      patterns[17618] = 25'b01000100_11010000_00010100_1;
      patterns[17619] = 25'b01000100_11010001_00010101_1;
      patterns[17620] = 25'b01000100_11010010_00010110_1;
      patterns[17621] = 25'b01000100_11010011_00010111_1;
      patterns[17622] = 25'b01000100_11010100_00011000_1;
      patterns[17623] = 25'b01000100_11010101_00011001_1;
      patterns[17624] = 25'b01000100_11010110_00011010_1;
      patterns[17625] = 25'b01000100_11010111_00011011_1;
      patterns[17626] = 25'b01000100_11011000_00011100_1;
      patterns[17627] = 25'b01000100_11011001_00011101_1;
      patterns[17628] = 25'b01000100_11011010_00011110_1;
      patterns[17629] = 25'b01000100_11011011_00011111_1;
      patterns[17630] = 25'b01000100_11011100_00100000_1;
      patterns[17631] = 25'b01000100_11011101_00100001_1;
      patterns[17632] = 25'b01000100_11011110_00100010_1;
      patterns[17633] = 25'b01000100_11011111_00100011_1;
      patterns[17634] = 25'b01000100_11100000_00100100_1;
      patterns[17635] = 25'b01000100_11100001_00100101_1;
      patterns[17636] = 25'b01000100_11100010_00100110_1;
      patterns[17637] = 25'b01000100_11100011_00100111_1;
      patterns[17638] = 25'b01000100_11100100_00101000_1;
      patterns[17639] = 25'b01000100_11100101_00101001_1;
      patterns[17640] = 25'b01000100_11100110_00101010_1;
      patterns[17641] = 25'b01000100_11100111_00101011_1;
      patterns[17642] = 25'b01000100_11101000_00101100_1;
      patterns[17643] = 25'b01000100_11101001_00101101_1;
      patterns[17644] = 25'b01000100_11101010_00101110_1;
      patterns[17645] = 25'b01000100_11101011_00101111_1;
      patterns[17646] = 25'b01000100_11101100_00110000_1;
      patterns[17647] = 25'b01000100_11101101_00110001_1;
      patterns[17648] = 25'b01000100_11101110_00110010_1;
      patterns[17649] = 25'b01000100_11101111_00110011_1;
      patterns[17650] = 25'b01000100_11110000_00110100_1;
      patterns[17651] = 25'b01000100_11110001_00110101_1;
      patterns[17652] = 25'b01000100_11110010_00110110_1;
      patterns[17653] = 25'b01000100_11110011_00110111_1;
      patterns[17654] = 25'b01000100_11110100_00111000_1;
      patterns[17655] = 25'b01000100_11110101_00111001_1;
      patterns[17656] = 25'b01000100_11110110_00111010_1;
      patterns[17657] = 25'b01000100_11110111_00111011_1;
      patterns[17658] = 25'b01000100_11111000_00111100_1;
      patterns[17659] = 25'b01000100_11111001_00111101_1;
      patterns[17660] = 25'b01000100_11111010_00111110_1;
      patterns[17661] = 25'b01000100_11111011_00111111_1;
      patterns[17662] = 25'b01000100_11111100_01000000_1;
      patterns[17663] = 25'b01000100_11111101_01000001_1;
      patterns[17664] = 25'b01000100_11111110_01000010_1;
      patterns[17665] = 25'b01000100_11111111_01000011_1;
      patterns[17666] = 25'b01000101_00000000_01000101_0;
      patterns[17667] = 25'b01000101_00000001_01000110_0;
      patterns[17668] = 25'b01000101_00000010_01000111_0;
      patterns[17669] = 25'b01000101_00000011_01001000_0;
      patterns[17670] = 25'b01000101_00000100_01001001_0;
      patterns[17671] = 25'b01000101_00000101_01001010_0;
      patterns[17672] = 25'b01000101_00000110_01001011_0;
      patterns[17673] = 25'b01000101_00000111_01001100_0;
      patterns[17674] = 25'b01000101_00001000_01001101_0;
      patterns[17675] = 25'b01000101_00001001_01001110_0;
      patterns[17676] = 25'b01000101_00001010_01001111_0;
      patterns[17677] = 25'b01000101_00001011_01010000_0;
      patterns[17678] = 25'b01000101_00001100_01010001_0;
      patterns[17679] = 25'b01000101_00001101_01010010_0;
      patterns[17680] = 25'b01000101_00001110_01010011_0;
      patterns[17681] = 25'b01000101_00001111_01010100_0;
      patterns[17682] = 25'b01000101_00010000_01010101_0;
      patterns[17683] = 25'b01000101_00010001_01010110_0;
      patterns[17684] = 25'b01000101_00010010_01010111_0;
      patterns[17685] = 25'b01000101_00010011_01011000_0;
      patterns[17686] = 25'b01000101_00010100_01011001_0;
      patterns[17687] = 25'b01000101_00010101_01011010_0;
      patterns[17688] = 25'b01000101_00010110_01011011_0;
      patterns[17689] = 25'b01000101_00010111_01011100_0;
      patterns[17690] = 25'b01000101_00011000_01011101_0;
      patterns[17691] = 25'b01000101_00011001_01011110_0;
      patterns[17692] = 25'b01000101_00011010_01011111_0;
      patterns[17693] = 25'b01000101_00011011_01100000_0;
      patterns[17694] = 25'b01000101_00011100_01100001_0;
      patterns[17695] = 25'b01000101_00011101_01100010_0;
      patterns[17696] = 25'b01000101_00011110_01100011_0;
      patterns[17697] = 25'b01000101_00011111_01100100_0;
      patterns[17698] = 25'b01000101_00100000_01100101_0;
      patterns[17699] = 25'b01000101_00100001_01100110_0;
      patterns[17700] = 25'b01000101_00100010_01100111_0;
      patterns[17701] = 25'b01000101_00100011_01101000_0;
      patterns[17702] = 25'b01000101_00100100_01101001_0;
      patterns[17703] = 25'b01000101_00100101_01101010_0;
      patterns[17704] = 25'b01000101_00100110_01101011_0;
      patterns[17705] = 25'b01000101_00100111_01101100_0;
      patterns[17706] = 25'b01000101_00101000_01101101_0;
      patterns[17707] = 25'b01000101_00101001_01101110_0;
      patterns[17708] = 25'b01000101_00101010_01101111_0;
      patterns[17709] = 25'b01000101_00101011_01110000_0;
      patterns[17710] = 25'b01000101_00101100_01110001_0;
      patterns[17711] = 25'b01000101_00101101_01110010_0;
      patterns[17712] = 25'b01000101_00101110_01110011_0;
      patterns[17713] = 25'b01000101_00101111_01110100_0;
      patterns[17714] = 25'b01000101_00110000_01110101_0;
      patterns[17715] = 25'b01000101_00110001_01110110_0;
      patterns[17716] = 25'b01000101_00110010_01110111_0;
      patterns[17717] = 25'b01000101_00110011_01111000_0;
      patterns[17718] = 25'b01000101_00110100_01111001_0;
      patterns[17719] = 25'b01000101_00110101_01111010_0;
      patterns[17720] = 25'b01000101_00110110_01111011_0;
      patterns[17721] = 25'b01000101_00110111_01111100_0;
      patterns[17722] = 25'b01000101_00111000_01111101_0;
      patterns[17723] = 25'b01000101_00111001_01111110_0;
      patterns[17724] = 25'b01000101_00111010_01111111_0;
      patterns[17725] = 25'b01000101_00111011_10000000_0;
      patterns[17726] = 25'b01000101_00111100_10000001_0;
      patterns[17727] = 25'b01000101_00111101_10000010_0;
      patterns[17728] = 25'b01000101_00111110_10000011_0;
      patterns[17729] = 25'b01000101_00111111_10000100_0;
      patterns[17730] = 25'b01000101_01000000_10000101_0;
      patterns[17731] = 25'b01000101_01000001_10000110_0;
      patterns[17732] = 25'b01000101_01000010_10000111_0;
      patterns[17733] = 25'b01000101_01000011_10001000_0;
      patterns[17734] = 25'b01000101_01000100_10001001_0;
      patterns[17735] = 25'b01000101_01000101_10001010_0;
      patterns[17736] = 25'b01000101_01000110_10001011_0;
      patterns[17737] = 25'b01000101_01000111_10001100_0;
      patterns[17738] = 25'b01000101_01001000_10001101_0;
      patterns[17739] = 25'b01000101_01001001_10001110_0;
      patterns[17740] = 25'b01000101_01001010_10001111_0;
      patterns[17741] = 25'b01000101_01001011_10010000_0;
      patterns[17742] = 25'b01000101_01001100_10010001_0;
      patterns[17743] = 25'b01000101_01001101_10010010_0;
      patterns[17744] = 25'b01000101_01001110_10010011_0;
      patterns[17745] = 25'b01000101_01001111_10010100_0;
      patterns[17746] = 25'b01000101_01010000_10010101_0;
      patterns[17747] = 25'b01000101_01010001_10010110_0;
      patterns[17748] = 25'b01000101_01010010_10010111_0;
      patterns[17749] = 25'b01000101_01010011_10011000_0;
      patterns[17750] = 25'b01000101_01010100_10011001_0;
      patterns[17751] = 25'b01000101_01010101_10011010_0;
      patterns[17752] = 25'b01000101_01010110_10011011_0;
      patterns[17753] = 25'b01000101_01010111_10011100_0;
      patterns[17754] = 25'b01000101_01011000_10011101_0;
      patterns[17755] = 25'b01000101_01011001_10011110_0;
      patterns[17756] = 25'b01000101_01011010_10011111_0;
      patterns[17757] = 25'b01000101_01011011_10100000_0;
      patterns[17758] = 25'b01000101_01011100_10100001_0;
      patterns[17759] = 25'b01000101_01011101_10100010_0;
      patterns[17760] = 25'b01000101_01011110_10100011_0;
      patterns[17761] = 25'b01000101_01011111_10100100_0;
      patterns[17762] = 25'b01000101_01100000_10100101_0;
      patterns[17763] = 25'b01000101_01100001_10100110_0;
      patterns[17764] = 25'b01000101_01100010_10100111_0;
      patterns[17765] = 25'b01000101_01100011_10101000_0;
      patterns[17766] = 25'b01000101_01100100_10101001_0;
      patterns[17767] = 25'b01000101_01100101_10101010_0;
      patterns[17768] = 25'b01000101_01100110_10101011_0;
      patterns[17769] = 25'b01000101_01100111_10101100_0;
      patterns[17770] = 25'b01000101_01101000_10101101_0;
      patterns[17771] = 25'b01000101_01101001_10101110_0;
      patterns[17772] = 25'b01000101_01101010_10101111_0;
      patterns[17773] = 25'b01000101_01101011_10110000_0;
      patterns[17774] = 25'b01000101_01101100_10110001_0;
      patterns[17775] = 25'b01000101_01101101_10110010_0;
      patterns[17776] = 25'b01000101_01101110_10110011_0;
      patterns[17777] = 25'b01000101_01101111_10110100_0;
      patterns[17778] = 25'b01000101_01110000_10110101_0;
      patterns[17779] = 25'b01000101_01110001_10110110_0;
      patterns[17780] = 25'b01000101_01110010_10110111_0;
      patterns[17781] = 25'b01000101_01110011_10111000_0;
      patterns[17782] = 25'b01000101_01110100_10111001_0;
      patterns[17783] = 25'b01000101_01110101_10111010_0;
      patterns[17784] = 25'b01000101_01110110_10111011_0;
      patterns[17785] = 25'b01000101_01110111_10111100_0;
      patterns[17786] = 25'b01000101_01111000_10111101_0;
      patterns[17787] = 25'b01000101_01111001_10111110_0;
      patterns[17788] = 25'b01000101_01111010_10111111_0;
      patterns[17789] = 25'b01000101_01111011_11000000_0;
      patterns[17790] = 25'b01000101_01111100_11000001_0;
      patterns[17791] = 25'b01000101_01111101_11000010_0;
      patterns[17792] = 25'b01000101_01111110_11000011_0;
      patterns[17793] = 25'b01000101_01111111_11000100_0;
      patterns[17794] = 25'b01000101_10000000_11000101_0;
      patterns[17795] = 25'b01000101_10000001_11000110_0;
      patterns[17796] = 25'b01000101_10000010_11000111_0;
      patterns[17797] = 25'b01000101_10000011_11001000_0;
      patterns[17798] = 25'b01000101_10000100_11001001_0;
      patterns[17799] = 25'b01000101_10000101_11001010_0;
      patterns[17800] = 25'b01000101_10000110_11001011_0;
      patterns[17801] = 25'b01000101_10000111_11001100_0;
      patterns[17802] = 25'b01000101_10001000_11001101_0;
      patterns[17803] = 25'b01000101_10001001_11001110_0;
      patterns[17804] = 25'b01000101_10001010_11001111_0;
      patterns[17805] = 25'b01000101_10001011_11010000_0;
      patterns[17806] = 25'b01000101_10001100_11010001_0;
      patterns[17807] = 25'b01000101_10001101_11010010_0;
      patterns[17808] = 25'b01000101_10001110_11010011_0;
      patterns[17809] = 25'b01000101_10001111_11010100_0;
      patterns[17810] = 25'b01000101_10010000_11010101_0;
      patterns[17811] = 25'b01000101_10010001_11010110_0;
      patterns[17812] = 25'b01000101_10010010_11010111_0;
      patterns[17813] = 25'b01000101_10010011_11011000_0;
      patterns[17814] = 25'b01000101_10010100_11011001_0;
      patterns[17815] = 25'b01000101_10010101_11011010_0;
      patterns[17816] = 25'b01000101_10010110_11011011_0;
      patterns[17817] = 25'b01000101_10010111_11011100_0;
      patterns[17818] = 25'b01000101_10011000_11011101_0;
      patterns[17819] = 25'b01000101_10011001_11011110_0;
      patterns[17820] = 25'b01000101_10011010_11011111_0;
      patterns[17821] = 25'b01000101_10011011_11100000_0;
      patterns[17822] = 25'b01000101_10011100_11100001_0;
      patterns[17823] = 25'b01000101_10011101_11100010_0;
      patterns[17824] = 25'b01000101_10011110_11100011_0;
      patterns[17825] = 25'b01000101_10011111_11100100_0;
      patterns[17826] = 25'b01000101_10100000_11100101_0;
      patterns[17827] = 25'b01000101_10100001_11100110_0;
      patterns[17828] = 25'b01000101_10100010_11100111_0;
      patterns[17829] = 25'b01000101_10100011_11101000_0;
      patterns[17830] = 25'b01000101_10100100_11101001_0;
      patterns[17831] = 25'b01000101_10100101_11101010_0;
      patterns[17832] = 25'b01000101_10100110_11101011_0;
      patterns[17833] = 25'b01000101_10100111_11101100_0;
      patterns[17834] = 25'b01000101_10101000_11101101_0;
      patterns[17835] = 25'b01000101_10101001_11101110_0;
      patterns[17836] = 25'b01000101_10101010_11101111_0;
      patterns[17837] = 25'b01000101_10101011_11110000_0;
      patterns[17838] = 25'b01000101_10101100_11110001_0;
      patterns[17839] = 25'b01000101_10101101_11110010_0;
      patterns[17840] = 25'b01000101_10101110_11110011_0;
      patterns[17841] = 25'b01000101_10101111_11110100_0;
      patterns[17842] = 25'b01000101_10110000_11110101_0;
      patterns[17843] = 25'b01000101_10110001_11110110_0;
      patterns[17844] = 25'b01000101_10110010_11110111_0;
      patterns[17845] = 25'b01000101_10110011_11111000_0;
      patterns[17846] = 25'b01000101_10110100_11111001_0;
      patterns[17847] = 25'b01000101_10110101_11111010_0;
      patterns[17848] = 25'b01000101_10110110_11111011_0;
      patterns[17849] = 25'b01000101_10110111_11111100_0;
      patterns[17850] = 25'b01000101_10111000_11111101_0;
      patterns[17851] = 25'b01000101_10111001_11111110_0;
      patterns[17852] = 25'b01000101_10111010_11111111_0;
      patterns[17853] = 25'b01000101_10111011_00000000_1;
      patterns[17854] = 25'b01000101_10111100_00000001_1;
      patterns[17855] = 25'b01000101_10111101_00000010_1;
      patterns[17856] = 25'b01000101_10111110_00000011_1;
      patterns[17857] = 25'b01000101_10111111_00000100_1;
      patterns[17858] = 25'b01000101_11000000_00000101_1;
      patterns[17859] = 25'b01000101_11000001_00000110_1;
      patterns[17860] = 25'b01000101_11000010_00000111_1;
      patterns[17861] = 25'b01000101_11000011_00001000_1;
      patterns[17862] = 25'b01000101_11000100_00001001_1;
      patterns[17863] = 25'b01000101_11000101_00001010_1;
      patterns[17864] = 25'b01000101_11000110_00001011_1;
      patterns[17865] = 25'b01000101_11000111_00001100_1;
      patterns[17866] = 25'b01000101_11001000_00001101_1;
      patterns[17867] = 25'b01000101_11001001_00001110_1;
      patterns[17868] = 25'b01000101_11001010_00001111_1;
      patterns[17869] = 25'b01000101_11001011_00010000_1;
      patterns[17870] = 25'b01000101_11001100_00010001_1;
      patterns[17871] = 25'b01000101_11001101_00010010_1;
      patterns[17872] = 25'b01000101_11001110_00010011_1;
      patterns[17873] = 25'b01000101_11001111_00010100_1;
      patterns[17874] = 25'b01000101_11010000_00010101_1;
      patterns[17875] = 25'b01000101_11010001_00010110_1;
      patterns[17876] = 25'b01000101_11010010_00010111_1;
      patterns[17877] = 25'b01000101_11010011_00011000_1;
      patterns[17878] = 25'b01000101_11010100_00011001_1;
      patterns[17879] = 25'b01000101_11010101_00011010_1;
      patterns[17880] = 25'b01000101_11010110_00011011_1;
      patterns[17881] = 25'b01000101_11010111_00011100_1;
      patterns[17882] = 25'b01000101_11011000_00011101_1;
      patterns[17883] = 25'b01000101_11011001_00011110_1;
      patterns[17884] = 25'b01000101_11011010_00011111_1;
      patterns[17885] = 25'b01000101_11011011_00100000_1;
      patterns[17886] = 25'b01000101_11011100_00100001_1;
      patterns[17887] = 25'b01000101_11011101_00100010_1;
      patterns[17888] = 25'b01000101_11011110_00100011_1;
      patterns[17889] = 25'b01000101_11011111_00100100_1;
      patterns[17890] = 25'b01000101_11100000_00100101_1;
      patterns[17891] = 25'b01000101_11100001_00100110_1;
      patterns[17892] = 25'b01000101_11100010_00100111_1;
      patterns[17893] = 25'b01000101_11100011_00101000_1;
      patterns[17894] = 25'b01000101_11100100_00101001_1;
      patterns[17895] = 25'b01000101_11100101_00101010_1;
      patterns[17896] = 25'b01000101_11100110_00101011_1;
      patterns[17897] = 25'b01000101_11100111_00101100_1;
      patterns[17898] = 25'b01000101_11101000_00101101_1;
      patterns[17899] = 25'b01000101_11101001_00101110_1;
      patterns[17900] = 25'b01000101_11101010_00101111_1;
      patterns[17901] = 25'b01000101_11101011_00110000_1;
      patterns[17902] = 25'b01000101_11101100_00110001_1;
      patterns[17903] = 25'b01000101_11101101_00110010_1;
      patterns[17904] = 25'b01000101_11101110_00110011_1;
      patterns[17905] = 25'b01000101_11101111_00110100_1;
      patterns[17906] = 25'b01000101_11110000_00110101_1;
      patterns[17907] = 25'b01000101_11110001_00110110_1;
      patterns[17908] = 25'b01000101_11110010_00110111_1;
      patterns[17909] = 25'b01000101_11110011_00111000_1;
      patterns[17910] = 25'b01000101_11110100_00111001_1;
      patterns[17911] = 25'b01000101_11110101_00111010_1;
      patterns[17912] = 25'b01000101_11110110_00111011_1;
      patterns[17913] = 25'b01000101_11110111_00111100_1;
      patterns[17914] = 25'b01000101_11111000_00111101_1;
      patterns[17915] = 25'b01000101_11111001_00111110_1;
      patterns[17916] = 25'b01000101_11111010_00111111_1;
      patterns[17917] = 25'b01000101_11111011_01000000_1;
      patterns[17918] = 25'b01000101_11111100_01000001_1;
      patterns[17919] = 25'b01000101_11111101_01000010_1;
      patterns[17920] = 25'b01000101_11111110_01000011_1;
      patterns[17921] = 25'b01000101_11111111_01000100_1;
      patterns[17922] = 25'b01000110_00000000_01000110_0;
      patterns[17923] = 25'b01000110_00000001_01000111_0;
      patterns[17924] = 25'b01000110_00000010_01001000_0;
      patterns[17925] = 25'b01000110_00000011_01001001_0;
      patterns[17926] = 25'b01000110_00000100_01001010_0;
      patterns[17927] = 25'b01000110_00000101_01001011_0;
      patterns[17928] = 25'b01000110_00000110_01001100_0;
      patterns[17929] = 25'b01000110_00000111_01001101_0;
      patterns[17930] = 25'b01000110_00001000_01001110_0;
      patterns[17931] = 25'b01000110_00001001_01001111_0;
      patterns[17932] = 25'b01000110_00001010_01010000_0;
      patterns[17933] = 25'b01000110_00001011_01010001_0;
      patterns[17934] = 25'b01000110_00001100_01010010_0;
      patterns[17935] = 25'b01000110_00001101_01010011_0;
      patterns[17936] = 25'b01000110_00001110_01010100_0;
      patterns[17937] = 25'b01000110_00001111_01010101_0;
      patterns[17938] = 25'b01000110_00010000_01010110_0;
      patterns[17939] = 25'b01000110_00010001_01010111_0;
      patterns[17940] = 25'b01000110_00010010_01011000_0;
      patterns[17941] = 25'b01000110_00010011_01011001_0;
      patterns[17942] = 25'b01000110_00010100_01011010_0;
      patterns[17943] = 25'b01000110_00010101_01011011_0;
      patterns[17944] = 25'b01000110_00010110_01011100_0;
      patterns[17945] = 25'b01000110_00010111_01011101_0;
      patterns[17946] = 25'b01000110_00011000_01011110_0;
      patterns[17947] = 25'b01000110_00011001_01011111_0;
      patterns[17948] = 25'b01000110_00011010_01100000_0;
      patterns[17949] = 25'b01000110_00011011_01100001_0;
      patterns[17950] = 25'b01000110_00011100_01100010_0;
      patterns[17951] = 25'b01000110_00011101_01100011_0;
      patterns[17952] = 25'b01000110_00011110_01100100_0;
      patterns[17953] = 25'b01000110_00011111_01100101_0;
      patterns[17954] = 25'b01000110_00100000_01100110_0;
      patterns[17955] = 25'b01000110_00100001_01100111_0;
      patterns[17956] = 25'b01000110_00100010_01101000_0;
      patterns[17957] = 25'b01000110_00100011_01101001_0;
      patterns[17958] = 25'b01000110_00100100_01101010_0;
      patterns[17959] = 25'b01000110_00100101_01101011_0;
      patterns[17960] = 25'b01000110_00100110_01101100_0;
      patterns[17961] = 25'b01000110_00100111_01101101_0;
      patterns[17962] = 25'b01000110_00101000_01101110_0;
      patterns[17963] = 25'b01000110_00101001_01101111_0;
      patterns[17964] = 25'b01000110_00101010_01110000_0;
      patterns[17965] = 25'b01000110_00101011_01110001_0;
      patterns[17966] = 25'b01000110_00101100_01110010_0;
      patterns[17967] = 25'b01000110_00101101_01110011_0;
      patterns[17968] = 25'b01000110_00101110_01110100_0;
      patterns[17969] = 25'b01000110_00101111_01110101_0;
      patterns[17970] = 25'b01000110_00110000_01110110_0;
      patterns[17971] = 25'b01000110_00110001_01110111_0;
      patterns[17972] = 25'b01000110_00110010_01111000_0;
      patterns[17973] = 25'b01000110_00110011_01111001_0;
      patterns[17974] = 25'b01000110_00110100_01111010_0;
      patterns[17975] = 25'b01000110_00110101_01111011_0;
      patterns[17976] = 25'b01000110_00110110_01111100_0;
      patterns[17977] = 25'b01000110_00110111_01111101_0;
      patterns[17978] = 25'b01000110_00111000_01111110_0;
      patterns[17979] = 25'b01000110_00111001_01111111_0;
      patterns[17980] = 25'b01000110_00111010_10000000_0;
      patterns[17981] = 25'b01000110_00111011_10000001_0;
      patterns[17982] = 25'b01000110_00111100_10000010_0;
      patterns[17983] = 25'b01000110_00111101_10000011_0;
      patterns[17984] = 25'b01000110_00111110_10000100_0;
      patterns[17985] = 25'b01000110_00111111_10000101_0;
      patterns[17986] = 25'b01000110_01000000_10000110_0;
      patterns[17987] = 25'b01000110_01000001_10000111_0;
      patterns[17988] = 25'b01000110_01000010_10001000_0;
      patterns[17989] = 25'b01000110_01000011_10001001_0;
      patterns[17990] = 25'b01000110_01000100_10001010_0;
      patterns[17991] = 25'b01000110_01000101_10001011_0;
      patterns[17992] = 25'b01000110_01000110_10001100_0;
      patterns[17993] = 25'b01000110_01000111_10001101_0;
      patterns[17994] = 25'b01000110_01001000_10001110_0;
      patterns[17995] = 25'b01000110_01001001_10001111_0;
      patterns[17996] = 25'b01000110_01001010_10010000_0;
      patterns[17997] = 25'b01000110_01001011_10010001_0;
      patterns[17998] = 25'b01000110_01001100_10010010_0;
      patterns[17999] = 25'b01000110_01001101_10010011_0;
      patterns[18000] = 25'b01000110_01001110_10010100_0;
      patterns[18001] = 25'b01000110_01001111_10010101_0;
      patterns[18002] = 25'b01000110_01010000_10010110_0;
      patterns[18003] = 25'b01000110_01010001_10010111_0;
      patterns[18004] = 25'b01000110_01010010_10011000_0;
      patterns[18005] = 25'b01000110_01010011_10011001_0;
      patterns[18006] = 25'b01000110_01010100_10011010_0;
      patterns[18007] = 25'b01000110_01010101_10011011_0;
      patterns[18008] = 25'b01000110_01010110_10011100_0;
      patterns[18009] = 25'b01000110_01010111_10011101_0;
      patterns[18010] = 25'b01000110_01011000_10011110_0;
      patterns[18011] = 25'b01000110_01011001_10011111_0;
      patterns[18012] = 25'b01000110_01011010_10100000_0;
      patterns[18013] = 25'b01000110_01011011_10100001_0;
      patterns[18014] = 25'b01000110_01011100_10100010_0;
      patterns[18015] = 25'b01000110_01011101_10100011_0;
      patterns[18016] = 25'b01000110_01011110_10100100_0;
      patterns[18017] = 25'b01000110_01011111_10100101_0;
      patterns[18018] = 25'b01000110_01100000_10100110_0;
      patterns[18019] = 25'b01000110_01100001_10100111_0;
      patterns[18020] = 25'b01000110_01100010_10101000_0;
      patterns[18021] = 25'b01000110_01100011_10101001_0;
      patterns[18022] = 25'b01000110_01100100_10101010_0;
      patterns[18023] = 25'b01000110_01100101_10101011_0;
      patterns[18024] = 25'b01000110_01100110_10101100_0;
      patterns[18025] = 25'b01000110_01100111_10101101_0;
      patterns[18026] = 25'b01000110_01101000_10101110_0;
      patterns[18027] = 25'b01000110_01101001_10101111_0;
      patterns[18028] = 25'b01000110_01101010_10110000_0;
      patterns[18029] = 25'b01000110_01101011_10110001_0;
      patterns[18030] = 25'b01000110_01101100_10110010_0;
      patterns[18031] = 25'b01000110_01101101_10110011_0;
      patterns[18032] = 25'b01000110_01101110_10110100_0;
      patterns[18033] = 25'b01000110_01101111_10110101_0;
      patterns[18034] = 25'b01000110_01110000_10110110_0;
      patterns[18035] = 25'b01000110_01110001_10110111_0;
      patterns[18036] = 25'b01000110_01110010_10111000_0;
      patterns[18037] = 25'b01000110_01110011_10111001_0;
      patterns[18038] = 25'b01000110_01110100_10111010_0;
      patterns[18039] = 25'b01000110_01110101_10111011_0;
      patterns[18040] = 25'b01000110_01110110_10111100_0;
      patterns[18041] = 25'b01000110_01110111_10111101_0;
      patterns[18042] = 25'b01000110_01111000_10111110_0;
      patterns[18043] = 25'b01000110_01111001_10111111_0;
      patterns[18044] = 25'b01000110_01111010_11000000_0;
      patterns[18045] = 25'b01000110_01111011_11000001_0;
      patterns[18046] = 25'b01000110_01111100_11000010_0;
      patterns[18047] = 25'b01000110_01111101_11000011_0;
      patterns[18048] = 25'b01000110_01111110_11000100_0;
      patterns[18049] = 25'b01000110_01111111_11000101_0;
      patterns[18050] = 25'b01000110_10000000_11000110_0;
      patterns[18051] = 25'b01000110_10000001_11000111_0;
      patterns[18052] = 25'b01000110_10000010_11001000_0;
      patterns[18053] = 25'b01000110_10000011_11001001_0;
      patterns[18054] = 25'b01000110_10000100_11001010_0;
      patterns[18055] = 25'b01000110_10000101_11001011_0;
      patterns[18056] = 25'b01000110_10000110_11001100_0;
      patterns[18057] = 25'b01000110_10000111_11001101_0;
      patterns[18058] = 25'b01000110_10001000_11001110_0;
      patterns[18059] = 25'b01000110_10001001_11001111_0;
      patterns[18060] = 25'b01000110_10001010_11010000_0;
      patterns[18061] = 25'b01000110_10001011_11010001_0;
      patterns[18062] = 25'b01000110_10001100_11010010_0;
      patterns[18063] = 25'b01000110_10001101_11010011_0;
      patterns[18064] = 25'b01000110_10001110_11010100_0;
      patterns[18065] = 25'b01000110_10001111_11010101_0;
      patterns[18066] = 25'b01000110_10010000_11010110_0;
      patterns[18067] = 25'b01000110_10010001_11010111_0;
      patterns[18068] = 25'b01000110_10010010_11011000_0;
      patterns[18069] = 25'b01000110_10010011_11011001_0;
      patterns[18070] = 25'b01000110_10010100_11011010_0;
      patterns[18071] = 25'b01000110_10010101_11011011_0;
      patterns[18072] = 25'b01000110_10010110_11011100_0;
      patterns[18073] = 25'b01000110_10010111_11011101_0;
      patterns[18074] = 25'b01000110_10011000_11011110_0;
      patterns[18075] = 25'b01000110_10011001_11011111_0;
      patterns[18076] = 25'b01000110_10011010_11100000_0;
      patterns[18077] = 25'b01000110_10011011_11100001_0;
      patterns[18078] = 25'b01000110_10011100_11100010_0;
      patterns[18079] = 25'b01000110_10011101_11100011_0;
      patterns[18080] = 25'b01000110_10011110_11100100_0;
      patterns[18081] = 25'b01000110_10011111_11100101_0;
      patterns[18082] = 25'b01000110_10100000_11100110_0;
      patterns[18083] = 25'b01000110_10100001_11100111_0;
      patterns[18084] = 25'b01000110_10100010_11101000_0;
      patterns[18085] = 25'b01000110_10100011_11101001_0;
      patterns[18086] = 25'b01000110_10100100_11101010_0;
      patterns[18087] = 25'b01000110_10100101_11101011_0;
      patterns[18088] = 25'b01000110_10100110_11101100_0;
      patterns[18089] = 25'b01000110_10100111_11101101_0;
      patterns[18090] = 25'b01000110_10101000_11101110_0;
      patterns[18091] = 25'b01000110_10101001_11101111_0;
      patterns[18092] = 25'b01000110_10101010_11110000_0;
      patterns[18093] = 25'b01000110_10101011_11110001_0;
      patterns[18094] = 25'b01000110_10101100_11110010_0;
      patterns[18095] = 25'b01000110_10101101_11110011_0;
      patterns[18096] = 25'b01000110_10101110_11110100_0;
      patterns[18097] = 25'b01000110_10101111_11110101_0;
      patterns[18098] = 25'b01000110_10110000_11110110_0;
      patterns[18099] = 25'b01000110_10110001_11110111_0;
      patterns[18100] = 25'b01000110_10110010_11111000_0;
      patterns[18101] = 25'b01000110_10110011_11111001_0;
      patterns[18102] = 25'b01000110_10110100_11111010_0;
      patterns[18103] = 25'b01000110_10110101_11111011_0;
      patterns[18104] = 25'b01000110_10110110_11111100_0;
      patterns[18105] = 25'b01000110_10110111_11111101_0;
      patterns[18106] = 25'b01000110_10111000_11111110_0;
      patterns[18107] = 25'b01000110_10111001_11111111_0;
      patterns[18108] = 25'b01000110_10111010_00000000_1;
      patterns[18109] = 25'b01000110_10111011_00000001_1;
      patterns[18110] = 25'b01000110_10111100_00000010_1;
      patterns[18111] = 25'b01000110_10111101_00000011_1;
      patterns[18112] = 25'b01000110_10111110_00000100_1;
      patterns[18113] = 25'b01000110_10111111_00000101_1;
      patterns[18114] = 25'b01000110_11000000_00000110_1;
      patterns[18115] = 25'b01000110_11000001_00000111_1;
      patterns[18116] = 25'b01000110_11000010_00001000_1;
      patterns[18117] = 25'b01000110_11000011_00001001_1;
      patterns[18118] = 25'b01000110_11000100_00001010_1;
      patterns[18119] = 25'b01000110_11000101_00001011_1;
      patterns[18120] = 25'b01000110_11000110_00001100_1;
      patterns[18121] = 25'b01000110_11000111_00001101_1;
      patterns[18122] = 25'b01000110_11001000_00001110_1;
      patterns[18123] = 25'b01000110_11001001_00001111_1;
      patterns[18124] = 25'b01000110_11001010_00010000_1;
      patterns[18125] = 25'b01000110_11001011_00010001_1;
      patterns[18126] = 25'b01000110_11001100_00010010_1;
      patterns[18127] = 25'b01000110_11001101_00010011_1;
      patterns[18128] = 25'b01000110_11001110_00010100_1;
      patterns[18129] = 25'b01000110_11001111_00010101_1;
      patterns[18130] = 25'b01000110_11010000_00010110_1;
      patterns[18131] = 25'b01000110_11010001_00010111_1;
      patterns[18132] = 25'b01000110_11010010_00011000_1;
      patterns[18133] = 25'b01000110_11010011_00011001_1;
      patterns[18134] = 25'b01000110_11010100_00011010_1;
      patterns[18135] = 25'b01000110_11010101_00011011_1;
      patterns[18136] = 25'b01000110_11010110_00011100_1;
      patterns[18137] = 25'b01000110_11010111_00011101_1;
      patterns[18138] = 25'b01000110_11011000_00011110_1;
      patterns[18139] = 25'b01000110_11011001_00011111_1;
      patterns[18140] = 25'b01000110_11011010_00100000_1;
      patterns[18141] = 25'b01000110_11011011_00100001_1;
      patterns[18142] = 25'b01000110_11011100_00100010_1;
      patterns[18143] = 25'b01000110_11011101_00100011_1;
      patterns[18144] = 25'b01000110_11011110_00100100_1;
      patterns[18145] = 25'b01000110_11011111_00100101_1;
      patterns[18146] = 25'b01000110_11100000_00100110_1;
      patterns[18147] = 25'b01000110_11100001_00100111_1;
      patterns[18148] = 25'b01000110_11100010_00101000_1;
      patterns[18149] = 25'b01000110_11100011_00101001_1;
      patterns[18150] = 25'b01000110_11100100_00101010_1;
      patterns[18151] = 25'b01000110_11100101_00101011_1;
      patterns[18152] = 25'b01000110_11100110_00101100_1;
      patterns[18153] = 25'b01000110_11100111_00101101_1;
      patterns[18154] = 25'b01000110_11101000_00101110_1;
      patterns[18155] = 25'b01000110_11101001_00101111_1;
      patterns[18156] = 25'b01000110_11101010_00110000_1;
      patterns[18157] = 25'b01000110_11101011_00110001_1;
      patterns[18158] = 25'b01000110_11101100_00110010_1;
      patterns[18159] = 25'b01000110_11101101_00110011_1;
      patterns[18160] = 25'b01000110_11101110_00110100_1;
      patterns[18161] = 25'b01000110_11101111_00110101_1;
      patterns[18162] = 25'b01000110_11110000_00110110_1;
      patterns[18163] = 25'b01000110_11110001_00110111_1;
      patterns[18164] = 25'b01000110_11110010_00111000_1;
      patterns[18165] = 25'b01000110_11110011_00111001_1;
      patterns[18166] = 25'b01000110_11110100_00111010_1;
      patterns[18167] = 25'b01000110_11110101_00111011_1;
      patterns[18168] = 25'b01000110_11110110_00111100_1;
      patterns[18169] = 25'b01000110_11110111_00111101_1;
      patterns[18170] = 25'b01000110_11111000_00111110_1;
      patterns[18171] = 25'b01000110_11111001_00111111_1;
      patterns[18172] = 25'b01000110_11111010_01000000_1;
      patterns[18173] = 25'b01000110_11111011_01000001_1;
      patterns[18174] = 25'b01000110_11111100_01000010_1;
      patterns[18175] = 25'b01000110_11111101_01000011_1;
      patterns[18176] = 25'b01000110_11111110_01000100_1;
      patterns[18177] = 25'b01000110_11111111_01000101_1;
      patterns[18178] = 25'b01000111_00000000_01000111_0;
      patterns[18179] = 25'b01000111_00000001_01001000_0;
      patterns[18180] = 25'b01000111_00000010_01001001_0;
      patterns[18181] = 25'b01000111_00000011_01001010_0;
      patterns[18182] = 25'b01000111_00000100_01001011_0;
      patterns[18183] = 25'b01000111_00000101_01001100_0;
      patterns[18184] = 25'b01000111_00000110_01001101_0;
      patterns[18185] = 25'b01000111_00000111_01001110_0;
      patterns[18186] = 25'b01000111_00001000_01001111_0;
      patterns[18187] = 25'b01000111_00001001_01010000_0;
      patterns[18188] = 25'b01000111_00001010_01010001_0;
      patterns[18189] = 25'b01000111_00001011_01010010_0;
      patterns[18190] = 25'b01000111_00001100_01010011_0;
      patterns[18191] = 25'b01000111_00001101_01010100_0;
      patterns[18192] = 25'b01000111_00001110_01010101_0;
      patterns[18193] = 25'b01000111_00001111_01010110_0;
      patterns[18194] = 25'b01000111_00010000_01010111_0;
      patterns[18195] = 25'b01000111_00010001_01011000_0;
      patterns[18196] = 25'b01000111_00010010_01011001_0;
      patterns[18197] = 25'b01000111_00010011_01011010_0;
      patterns[18198] = 25'b01000111_00010100_01011011_0;
      patterns[18199] = 25'b01000111_00010101_01011100_0;
      patterns[18200] = 25'b01000111_00010110_01011101_0;
      patterns[18201] = 25'b01000111_00010111_01011110_0;
      patterns[18202] = 25'b01000111_00011000_01011111_0;
      patterns[18203] = 25'b01000111_00011001_01100000_0;
      patterns[18204] = 25'b01000111_00011010_01100001_0;
      patterns[18205] = 25'b01000111_00011011_01100010_0;
      patterns[18206] = 25'b01000111_00011100_01100011_0;
      patterns[18207] = 25'b01000111_00011101_01100100_0;
      patterns[18208] = 25'b01000111_00011110_01100101_0;
      patterns[18209] = 25'b01000111_00011111_01100110_0;
      patterns[18210] = 25'b01000111_00100000_01100111_0;
      patterns[18211] = 25'b01000111_00100001_01101000_0;
      patterns[18212] = 25'b01000111_00100010_01101001_0;
      patterns[18213] = 25'b01000111_00100011_01101010_0;
      patterns[18214] = 25'b01000111_00100100_01101011_0;
      patterns[18215] = 25'b01000111_00100101_01101100_0;
      patterns[18216] = 25'b01000111_00100110_01101101_0;
      patterns[18217] = 25'b01000111_00100111_01101110_0;
      patterns[18218] = 25'b01000111_00101000_01101111_0;
      patterns[18219] = 25'b01000111_00101001_01110000_0;
      patterns[18220] = 25'b01000111_00101010_01110001_0;
      patterns[18221] = 25'b01000111_00101011_01110010_0;
      patterns[18222] = 25'b01000111_00101100_01110011_0;
      patterns[18223] = 25'b01000111_00101101_01110100_0;
      patterns[18224] = 25'b01000111_00101110_01110101_0;
      patterns[18225] = 25'b01000111_00101111_01110110_0;
      patterns[18226] = 25'b01000111_00110000_01110111_0;
      patterns[18227] = 25'b01000111_00110001_01111000_0;
      patterns[18228] = 25'b01000111_00110010_01111001_0;
      patterns[18229] = 25'b01000111_00110011_01111010_0;
      patterns[18230] = 25'b01000111_00110100_01111011_0;
      patterns[18231] = 25'b01000111_00110101_01111100_0;
      patterns[18232] = 25'b01000111_00110110_01111101_0;
      patterns[18233] = 25'b01000111_00110111_01111110_0;
      patterns[18234] = 25'b01000111_00111000_01111111_0;
      patterns[18235] = 25'b01000111_00111001_10000000_0;
      patterns[18236] = 25'b01000111_00111010_10000001_0;
      patterns[18237] = 25'b01000111_00111011_10000010_0;
      patterns[18238] = 25'b01000111_00111100_10000011_0;
      patterns[18239] = 25'b01000111_00111101_10000100_0;
      patterns[18240] = 25'b01000111_00111110_10000101_0;
      patterns[18241] = 25'b01000111_00111111_10000110_0;
      patterns[18242] = 25'b01000111_01000000_10000111_0;
      patterns[18243] = 25'b01000111_01000001_10001000_0;
      patterns[18244] = 25'b01000111_01000010_10001001_0;
      patterns[18245] = 25'b01000111_01000011_10001010_0;
      patterns[18246] = 25'b01000111_01000100_10001011_0;
      patterns[18247] = 25'b01000111_01000101_10001100_0;
      patterns[18248] = 25'b01000111_01000110_10001101_0;
      patterns[18249] = 25'b01000111_01000111_10001110_0;
      patterns[18250] = 25'b01000111_01001000_10001111_0;
      patterns[18251] = 25'b01000111_01001001_10010000_0;
      patterns[18252] = 25'b01000111_01001010_10010001_0;
      patterns[18253] = 25'b01000111_01001011_10010010_0;
      patterns[18254] = 25'b01000111_01001100_10010011_0;
      patterns[18255] = 25'b01000111_01001101_10010100_0;
      patterns[18256] = 25'b01000111_01001110_10010101_0;
      patterns[18257] = 25'b01000111_01001111_10010110_0;
      patterns[18258] = 25'b01000111_01010000_10010111_0;
      patterns[18259] = 25'b01000111_01010001_10011000_0;
      patterns[18260] = 25'b01000111_01010010_10011001_0;
      patterns[18261] = 25'b01000111_01010011_10011010_0;
      patterns[18262] = 25'b01000111_01010100_10011011_0;
      patterns[18263] = 25'b01000111_01010101_10011100_0;
      patterns[18264] = 25'b01000111_01010110_10011101_0;
      patterns[18265] = 25'b01000111_01010111_10011110_0;
      patterns[18266] = 25'b01000111_01011000_10011111_0;
      patterns[18267] = 25'b01000111_01011001_10100000_0;
      patterns[18268] = 25'b01000111_01011010_10100001_0;
      patterns[18269] = 25'b01000111_01011011_10100010_0;
      patterns[18270] = 25'b01000111_01011100_10100011_0;
      patterns[18271] = 25'b01000111_01011101_10100100_0;
      patterns[18272] = 25'b01000111_01011110_10100101_0;
      patterns[18273] = 25'b01000111_01011111_10100110_0;
      patterns[18274] = 25'b01000111_01100000_10100111_0;
      patterns[18275] = 25'b01000111_01100001_10101000_0;
      patterns[18276] = 25'b01000111_01100010_10101001_0;
      patterns[18277] = 25'b01000111_01100011_10101010_0;
      patterns[18278] = 25'b01000111_01100100_10101011_0;
      patterns[18279] = 25'b01000111_01100101_10101100_0;
      patterns[18280] = 25'b01000111_01100110_10101101_0;
      patterns[18281] = 25'b01000111_01100111_10101110_0;
      patterns[18282] = 25'b01000111_01101000_10101111_0;
      patterns[18283] = 25'b01000111_01101001_10110000_0;
      patterns[18284] = 25'b01000111_01101010_10110001_0;
      patterns[18285] = 25'b01000111_01101011_10110010_0;
      patterns[18286] = 25'b01000111_01101100_10110011_0;
      patterns[18287] = 25'b01000111_01101101_10110100_0;
      patterns[18288] = 25'b01000111_01101110_10110101_0;
      patterns[18289] = 25'b01000111_01101111_10110110_0;
      patterns[18290] = 25'b01000111_01110000_10110111_0;
      patterns[18291] = 25'b01000111_01110001_10111000_0;
      patterns[18292] = 25'b01000111_01110010_10111001_0;
      patterns[18293] = 25'b01000111_01110011_10111010_0;
      patterns[18294] = 25'b01000111_01110100_10111011_0;
      patterns[18295] = 25'b01000111_01110101_10111100_0;
      patterns[18296] = 25'b01000111_01110110_10111101_0;
      patterns[18297] = 25'b01000111_01110111_10111110_0;
      patterns[18298] = 25'b01000111_01111000_10111111_0;
      patterns[18299] = 25'b01000111_01111001_11000000_0;
      patterns[18300] = 25'b01000111_01111010_11000001_0;
      patterns[18301] = 25'b01000111_01111011_11000010_0;
      patterns[18302] = 25'b01000111_01111100_11000011_0;
      patterns[18303] = 25'b01000111_01111101_11000100_0;
      patterns[18304] = 25'b01000111_01111110_11000101_0;
      patterns[18305] = 25'b01000111_01111111_11000110_0;
      patterns[18306] = 25'b01000111_10000000_11000111_0;
      patterns[18307] = 25'b01000111_10000001_11001000_0;
      patterns[18308] = 25'b01000111_10000010_11001001_0;
      patterns[18309] = 25'b01000111_10000011_11001010_0;
      patterns[18310] = 25'b01000111_10000100_11001011_0;
      patterns[18311] = 25'b01000111_10000101_11001100_0;
      patterns[18312] = 25'b01000111_10000110_11001101_0;
      patterns[18313] = 25'b01000111_10000111_11001110_0;
      patterns[18314] = 25'b01000111_10001000_11001111_0;
      patterns[18315] = 25'b01000111_10001001_11010000_0;
      patterns[18316] = 25'b01000111_10001010_11010001_0;
      patterns[18317] = 25'b01000111_10001011_11010010_0;
      patterns[18318] = 25'b01000111_10001100_11010011_0;
      patterns[18319] = 25'b01000111_10001101_11010100_0;
      patterns[18320] = 25'b01000111_10001110_11010101_0;
      patterns[18321] = 25'b01000111_10001111_11010110_0;
      patterns[18322] = 25'b01000111_10010000_11010111_0;
      patterns[18323] = 25'b01000111_10010001_11011000_0;
      patterns[18324] = 25'b01000111_10010010_11011001_0;
      patterns[18325] = 25'b01000111_10010011_11011010_0;
      patterns[18326] = 25'b01000111_10010100_11011011_0;
      patterns[18327] = 25'b01000111_10010101_11011100_0;
      patterns[18328] = 25'b01000111_10010110_11011101_0;
      patterns[18329] = 25'b01000111_10010111_11011110_0;
      patterns[18330] = 25'b01000111_10011000_11011111_0;
      patterns[18331] = 25'b01000111_10011001_11100000_0;
      patterns[18332] = 25'b01000111_10011010_11100001_0;
      patterns[18333] = 25'b01000111_10011011_11100010_0;
      patterns[18334] = 25'b01000111_10011100_11100011_0;
      patterns[18335] = 25'b01000111_10011101_11100100_0;
      patterns[18336] = 25'b01000111_10011110_11100101_0;
      patterns[18337] = 25'b01000111_10011111_11100110_0;
      patterns[18338] = 25'b01000111_10100000_11100111_0;
      patterns[18339] = 25'b01000111_10100001_11101000_0;
      patterns[18340] = 25'b01000111_10100010_11101001_0;
      patterns[18341] = 25'b01000111_10100011_11101010_0;
      patterns[18342] = 25'b01000111_10100100_11101011_0;
      patterns[18343] = 25'b01000111_10100101_11101100_0;
      patterns[18344] = 25'b01000111_10100110_11101101_0;
      patterns[18345] = 25'b01000111_10100111_11101110_0;
      patterns[18346] = 25'b01000111_10101000_11101111_0;
      patterns[18347] = 25'b01000111_10101001_11110000_0;
      patterns[18348] = 25'b01000111_10101010_11110001_0;
      patterns[18349] = 25'b01000111_10101011_11110010_0;
      patterns[18350] = 25'b01000111_10101100_11110011_0;
      patterns[18351] = 25'b01000111_10101101_11110100_0;
      patterns[18352] = 25'b01000111_10101110_11110101_0;
      patterns[18353] = 25'b01000111_10101111_11110110_0;
      patterns[18354] = 25'b01000111_10110000_11110111_0;
      patterns[18355] = 25'b01000111_10110001_11111000_0;
      patterns[18356] = 25'b01000111_10110010_11111001_0;
      patterns[18357] = 25'b01000111_10110011_11111010_0;
      patterns[18358] = 25'b01000111_10110100_11111011_0;
      patterns[18359] = 25'b01000111_10110101_11111100_0;
      patterns[18360] = 25'b01000111_10110110_11111101_0;
      patterns[18361] = 25'b01000111_10110111_11111110_0;
      patterns[18362] = 25'b01000111_10111000_11111111_0;
      patterns[18363] = 25'b01000111_10111001_00000000_1;
      patterns[18364] = 25'b01000111_10111010_00000001_1;
      patterns[18365] = 25'b01000111_10111011_00000010_1;
      patterns[18366] = 25'b01000111_10111100_00000011_1;
      patterns[18367] = 25'b01000111_10111101_00000100_1;
      patterns[18368] = 25'b01000111_10111110_00000101_1;
      patterns[18369] = 25'b01000111_10111111_00000110_1;
      patterns[18370] = 25'b01000111_11000000_00000111_1;
      patterns[18371] = 25'b01000111_11000001_00001000_1;
      patterns[18372] = 25'b01000111_11000010_00001001_1;
      patterns[18373] = 25'b01000111_11000011_00001010_1;
      patterns[18374] = 25'b01000111_11000100_00001011_1;
      patterns[18375] = 25'b01000111_11000101_00001100_1;
      patterns[18376] = 25'b01000111_11000110_00001101_1;
      patterns[18377] = 25'b01000111_11000111_00001110_1;
      patterns[18378] = 25'b01000111_11001000_00001111_1;
      patterns[18379] = 25'b01000111_11001001_00010000_1;
      patterns[18380] = 25'b01000111_11001010_00010001_1;
      patterns[18381] = 25'b01000111_11001011_00010010_1;
      patterns[18382] = 25'b01000111_11001100_00010011_1;
      patterns[18383] = 25'b01000111_11001101_00010100_1;
      patterns[18384] = 25'b01000111_11001110_00010101_1;
      patterns[18385] = 25'b01000111_11001111_00010110_1;
      patterns[18386] = 25'b01000111_11010000_00010111_1;
      patterns[18387] = 25'b01000111_11010001_00011000_1;
      patterns[18388] = 25'b01000111_11010010_00011001_1;
      patterns[18389] = 25'b01000111_11010011_00011010_1;
      patterns[18390] = 25'b01000111_11010100_00011011_1;
      patterns[18391] = 25'b01000111_11010101_00011100_1;
      patterns[18392] = 25'b01000111_11010110_00011101_1;
      patterns[18393] = 25'b01000111_11010111_00011110_1;
      patterns[18394] = 25'b01000111_11011000_00011111_1;
      patterns[18395] = 25'b01000111_11011001_00100000_1;
      patterns[18396] = 25'b01000111_11011010_00100001_1;
      patterns[18397] = 25'b01000111_11011011_00100010_1;
      patterns[18398] = 25'b01000111_11011100_00100011_1;
      patterns[18399] = 25'b01000111_11011101_00100100_1;
      patterns[18400] = 25'b01000111_11011110_00100101_1;
      patterns[18401] = 25'b01000111_11011111_00100110_1;
      patterns[18402] = 25'b01000111_11100000_00100111_1;
      patterns[18403] = 25'b01000111_11100001_00101000_1;
      patterns[18404] = 25'b01000111_11100010_00101001_1;
      patterns[18405] = 25'b01000111_11100011_00101010_1;
      patterns[18406] = 25'b01000111_11100100_00101011_1;
      patterns[18407] = 25'b01000111_11100101_00101100_1;
      patterns[18408] = 25'b01000111_11100110_00101101_1;
      patterns[18409] = 25'b01000111_11100111_00101110_1;
      patterns[18410] = 25'b01000111_11101000_00101111_1;
      patterns[18411] = 25'b01000111_11101001_00110000_1;
      patterns[18412] = 25'b01000111_11101010_00110001_1;
      patterns[18413] = 25'b01000111_11101011_00110010_1;
      patterns[18414] = 25'b01000111_11101100_00110011_1;
      patterns[18415] = 25'b01000111_11101101_00110100_1;
      patterns[18416] = 25'b01000111_11101110_00110101_1;
      patterns[18417] = 25'b01000111_11101111_00110110_1;
      patterns[18418] = 25'b01000111_11110000_00110111_1;
      patterns[18419] = 25'b01000111_11110001_00111000_1;
      patterns[18420] = 25'b01000111_11110010_00111001_1;
      patterns[18421] = 25'b01000111_11110011_00111010_1;
      patterns[18422] = 25'b01000111_11110100_00111011_1;
      patterns[18423] = 25'b01000111_11110101_00111100_1;
      patterns[18424] = 25'b01000111_11110110_00111101_1;
      patterns[18425] = 25'b01000111_11110111_00111110_1;
      patterns[18426] = 25'b01000111_11111000_00111111_1;
      patterns[18427] = 25'b01000111_11111001_01000000_1;
      patterns[18428] = 25'b01000111_11111010_01000001_1;
      patterns[18429] = 25'b01000111_11111011_01000010_1;
      patterns[18430] = 25'b01000111_11111100_01000011_1;
      patterns[18431] = 25'b01000111_11111101_01000100_1;
      patterns[18432] = 25'b01000111_11111110_01000101_1;
      patterns[18433] = 25'b01000111_11111111_01000110_1;
      patterns[18434] = 25'b01001000_00000000_01001000_0;
      patterns[18435] = 25'b01001000_00000001_01001001_0;
      patterns[18436] = 25'b01001000_00000010_01001010_0;
      patterns[18437] = 25'b01001000_00000011_01001011_0;
      patterns[18438] = 25'b01001000_00000100_01001100_0;
      patterns[18439] = 25'b01001000_00000101_01001101_0;
      patterns[18440] = 25'b01001000_00000110_01001110_0;
      patterns[18441] = 25'b01001000_00000111_01001111_0;
      patterns[18442] = 25'b01001000_00001000_01010000_0;
      patterns[18443] = 25'b01001000_00001001_01010001_0;
      patterns[18444] = 25'b01001000_00001010_01010010_0;
      patterns[18445] = 25'b01001000_00001011_01010011_0;
      patterns[18446] = 25'b01001000_00001100_01010100_0;
      patterns[18447] = 25'b01001000_00001101_01010101_0;
      patterns[18448] = 25'b01001000_00001110_01010110_0;
      patterns[18449] = 25'b01001000_00001111_01010111_0;
      patterns[18450] = 25'b01001000_00010000_01011000_0;
      patterns[18451] = 25'b01001000_00010001_01011001_0;
      patterns[18452] = 25'b01001000_00010010_01011010_0;
      patterns[18453] = 25'b01001000_00010011_01011011_0;
      patterns[18454] = 25'b01001000_00010100_01011100_0;
      patterns[18455] = 25'b01001000_00010101_01011101_0;
      patterns[18456] = 25'b01001000_00010110_01011110_0;
      patterns[18457] = 25'b01001000_00010111_01011111_0;
      patterns[18458] = 25'b01001000_00011000_01100000_0;
      patterns[18459] = 25'b01001000_00011001_01100001_0;
      patterns[18460] = 25'b01001000_00011010_01100010_0;
      patterns[18461] = 25'b01001000_00011011_01100011_0;
      patterns[18462] = 25'b01001000_00011100_01100100_0;
      patterns[18463] = 25'b01001000_00011101_01100101_0;
      patterns[18464] = 25'b01001000_00011110_01100110_0;
      patterns[18465] = 25'b01001000_00011111_01100111_0;
      patterns[18466] = 25'b01001000_00100000_01101000_0;
      patterns[18467] = 25'b01001000_00100001_01101001_0;
      patterns[18468] = 25'b01001000_00100010_01101010_0;
      patterns[18469] = 25'b01001000_00100011_01101011_0;
      patterns[18470] = 25'b01001000_00100100_01101100_0;
      patterns[18471] = 25'b01001000_00100101_01101101_0;
      patterns[18472] = 25'b01001000_00100110_01101110_0;
      patterns[18473] = 25'b01001000_00100111_01101111_0;
      patterns[18474] = 25'b01001000_00101000_01110000_0;
      patterns[18475] = 25'b01001000_00101001_01110001_0;
      patterns[18476] = 25'b01001000_00101010_01110010_0;
      patterns[18477] = 25'b01001000_00101011_01110011_0;
      patterns[18478] = 25'b01001000_00101100_01110100_0;
      patterns[18479] = 25'b01001000_00101101_01110101_0;
      patterns[18480] = 25'b01001000_00101110_01110110_0;
      patterns[18481] = 25'b01001000_00101111_01110111_0;
      patterns[18482] = 25'b01001000_00110000_01111000_0;
      patterns[18483] = 25'b01001000_00110001_01111001_0;
      patterns[18484] = 25'b01001000_00110010_01111010_0;
      patterns[18485] = 25'b01001000_00110011_01111011_0;
      patterns[18486] = 25'b01001000_00110100_01111100_0;
      patterns[18487] = 25'b01001000_00110101_01111101_0;
      patterns[18488] = 25'b01001000_00110110_01111110_0;
      patterns[18489] = 25'b01001000_00110111_01111111_0;
      patterns[18490] = 25'b01001000_00111000_10000000_0;
      patterns[18491] = 25'b01001000_00111001_10000001_0;
      patterns[18492] = 25'b01001000_00111010_10000010_0;
      patterns[18493] = 25'b01001000_00111011_10000011_0;
      patterns[18494] = 25'b01001000_00111100_10000100_0;
      patterns[18495] = 25'b01001000_00111101_10000101_0;
      patterns[18496] = 25'b01001000_00111110_10000110_0;
      patterns[18497] = 25'b01001000_00111111_10000111_0;
      patterns[18498] = 25'b01001000_01000000_10001000_0;
      patterns[18499] = 25'b01001000_01000001_10001001_0;
      patterns[18500] = 25'b01001000_01000010_10001010_0;
      patterns[18501] = 25'b01001000_01000011_10001011_0;
      patterns[18502] = 25'b01001000_01000100_10001100_0;
      patterns[18503] = 25'b01001000_01000101_10001101_0;
      patterns[18504] = 25'b01001000_01000110_10001110_0;
      patterns[18505] = 25'b01001000_01000111_10001111_0;
      patterns[18506] = 25'b01001000_01001000_10010000_0;
      patterns[18507] = 25'b01001000_01001001_10010001_0;
      patterns[18508] = 25'b01001000_01001010_10010010_0;
      patterns[18509] = 25'b01001000_01001011_10010011_0;
      patterns[18510] = 25'b01001000_01001100_10010100_0;
      patterns[18511] = 25'b01001000_01001101_10010101_0;
      patterns[18512] = 25'b01001000_01001110_10010110_0;
      patterns[18513] = 25'b01001000_01001111_10010111_0;
      patterns[18514] = 25'b01001000_01010000_10011000_0;
      patterns[18515] = 25'b01001000_01010001_10011001_0;
      patterns[18516] = 25'b01001000_01010010_10011010_0;
      patterns[18517] = 25'b01001000_01010011_10011011_0;
      patterns[18518] = 25'b01001000_01010100_10011100_0;
      patterns[18519] = 25'b01001000_01010101_10011101_0;
      patterns[18520] = 25'b01001000_01010110_10011110_0;
      patterns[18521] = 25'b01001000_01010111_10011111_0;
      patterns[18522] = 25'b01001000_01011000_10100000_0;
      patterns[18523] = 25'b01001000_01011001_10100001_0;
      patterns[18524] = 25'b01001000_01011010_10100010_0;
      patterns[18525] = 25'b01001000_01011011_10100011_0;
      patterns[18526] = 25'b01001000_01011100_10100100_0;
      patterns[18527] = 25'b01001000_01011101_10100101_0;
      patterns[18528] = 25'b01001000_01011110_10100110_0;
      patterns[18529] = 25'b01001000_01011111_10100111_0;
      patterns[18530] = 25'b01001000_01100000_10101000_0;
      patterns[18531] = 25'b01001000_01100001_10101001_0;
      patterns[18532] = 25'b01001000_01100010_10101010_0;
      patterns[18533] = 25'b01001000_01100011_10101011_0;
      patterns[18534] = 25'b01001000_01100100_10101100_0;
      patterns[18535] = 25'b01001000_01100101_10101101_0;
      patterns[18536] = 25'b01001000_01100110_10101110_0;
      patterns[18537] = 25'b01001000_01100111_10101111_0;
      patterns[18538] = 25'b01001000_01101000_10110000_0;
      patterns[18539] = 25'b01001000_01101001_10110001_0;
      patterns[18540] = 25'b01001000_01101010_10110010_0;
      patterns[18541] = 25'b01001000_01101011_10110011_0;
      patterns[18542] = 25'b01001000_01101100_10110100_0;
      patterns[18543] = 25'b01001000_01101101_10110101_0;
      patterns[18544] = 25'b01001000_01101110_10110110_0;
      patterns[18545] = 25'b01001000_01101111_10110111_0;
      patterns[18546] = 25'b01001000_01110000_10111000_0;
      patterns[18547] = 25'b01001000_01110001_10111001_0;
      patterns[18548] = 25'b01001000_01110010_10111010_0;
      patterns[18549] = 25'b01001000_01110011_10111011_0;
      patterns[18550] = 25'b01001000_01110100_10111100_0;
      patterns[18551] = 25'b01001000_01110101_10111101_0;
      patterns[18552] = 25'b01001000_01110110_10111110_0;
      patterns[18553] = 25'b01001000_01110111_10111111_0;
      patterns[18554] = 25'b01001000_01111000_11000000_0;
      patterns[18555] = 25'b01001000_01111001_11000001_0;
      patterns[18556] = 25'b01001000_01111010_11000010_0;
      patterns[18557] = 25'b01001000_01111011_11000011_0;
      patterns[18558] = 25'b01001000_01111100_11000100_0;
      patterns[18559] = 25'b01001000_01111101_11000101_0;
      patterns[18560] = 25'b01001000_01111110_11000110_0;
      patterns[18561] = 25'b01001000_01111111_11000111_0;
      patterns[18562] = 25'b01001000_10000000_11001000_0;
      patterns[18563] = 25'b01001000_10000001_11001001_0;
      patterns[18564] = 25'b01001000_10000010_11001010_0;
      patterns[18565] = 25'b01001000_10000011_11001011_0;
      patterns[18566] = 25'b01001000_10000100_11001100_0;
      patterns[18567] = 25'b01001000_10000101_11001101_0;
      patterns[18568] = 25'b01001000_10000110_11001110_0;
      patterns[18569] = 25'b01001000_10000111_11001111_0;
      patterns[18570] = 25'b01001000_10001000_11010000_0;
      patterns[18571] = 25'b01001000_10001001_11010001_0;
      patterns[18572] = 25'b01001000_10001010_11010010_0;
      patterns[18573] = 25'b01001000_10001011_11010011_0;
      patterns[18574] = 25'b01001000_10001100_11010100_0;
      patterns[18575] = 25'b01001000_10001101_11010101_0;
      patterns[18576] = 25'b01001000_10001110_11010110_0;
      patterns[18577] = 25'b01001000_10001111_11010111_0;
      patterns[18578] = 25'b01001000_10010000_11011000_0;
      patterns[18579] = 25'b01001000_10010001_11011001_0;
      patterns[18580] = 25'b01001000_10010010_11011010_0;
      patterns[18581] = 25'b01001000_10010011_11011011_0;
      patterns[18582] = 25'b01001000_10010100_11011100_0;
      patterns[18583] = 25'b01001000_10010101_11011101_0;
      patterns[18584] = 25'b01001000_10010110_11011110_0;
      patterns[18585] = 25'b01001000_10010111_11011111_0;
      patterns[18586] = 25'b01001000_10011000_11100000_0;
      patterns[18587] = 25'b01001000_10011001_11100001_0;
      patterns[18588] = 25'b01001000_10011010_11100010_0;
      patterns[18589] = 25'b01001000_10011011_11100011_0;
      patterns[18590] = 25'b01001000_10011100_11100100_0;
      patterns[18591] = 25'b01001000_10011101_11100101_0;
      patterns[18592] = 25'b01001000_10011110_11100110_0;
      patterns[18593] = 25'b01001000_10011111_11100111_0;
      patterns[18594] = 25'b01001000_10100000_11101000_0;
      patterns[18595] = 25'b01001000_10100001_11101001_0;
      patterns[18596] = 25'b01001000_10100010_11101010_0;
      patterns[18597] = 25'b01001000_10100011_11101011_0;
      patterns[18598] = 25'b01001000_10100100_11101100_0;
      patterns[18599] = 25'b01001000_10100101_11101101_0;
      patterns[18600] = 25'b01001000_10100110_11101110_0;
      patterns[18601] = 25'b01001000_10100111_11101111_0;
      patterns[18602] = 25'b01001000_10101000_11110000_0;
      patterns[18603] = 25'b01001000_10101001_11110001_0;
      patterns[18604] = 25'b01001000_10101010_11110010_0;
      patterns[18605] = 25'b01001000_10101011_11110011_0;
      patterns[18606] = 25'b01001000_10101100_11110100_0;
      patterns[18607] = 25'b01001000_10101101_11110101_0;
      patterns[18608] = 25'b01001000_10101110_11110110_0;
      patterns[18609] = 25'b01001000_10101111_11110111_0;
      patterns[18610] = 25'b01001000_10110000_11111000_0;
      patterns[18611] = 25'b01001000_10110001_11111001_0;
      patterns[18612] = 25'b01001000_10110010_11111010_0;
      patterns[18613] = 25'b01001000_10110011_11111011_0;
      patterns[18614] = 25'b01001000_10110100_11111100_0;
      patterns[18615] = 25'b01001000_10110101_11111101_0;
      patterns[18616] = 25'b01001000_10110110_11111110_0;
      patterns[18617] = 25'b01001000_10110111_11111111_0;
      patterns[18618] = 25'b01001000_10111000_00000000_1;
      patterns[18619] = 25'b01001000_10111001_00000001_1;
      patterns[18620] = 25'b01001000_10111010_00000010_1;
      patterns[18621] = 25'b01001000_10111011_00000011_1;
      patterns[18622] = 25'b01001000_10111100_00000100_1;
      patterns[18623] = 25'b01001000_10111101_00000101_1;
      patterns[18624] = 25'b01001000_10111110_00000110_1;
      patterns[18625] = 25'b01001000_10111111_00000111_1;
      patterns[18626] = 25'b01001000_11000000_00001000_1;
      patterns[18627] = 25'b01001000_11000001_00001001_1;
      patterns[18628] = 25'b01001000_11000010_00001010_1;
      patterns[18629] = 25'b01001000_11000011_00001011_1;
      patterns[18630] = 25'b01001000_11000100_00001100_1;
      patterns[18631] = 25'b01001000_11000101_00001101_1;
      patterns[18632] = 25'b01001000_11000110_00001110_1;
      patterns[18633] = 25'b01001000_11000111_00001111_1;
      patterns[18634] = 25'b01001000_11001000_00010000_1;
      patterns[18635] = 25'b01001000_11001001_00010001_1;
      patterns[18636] = 25'b01001000_11001010_00010010_1;
      patterns[18637] = 25'b01001000_11001011_00010011_1;
      patterns[18638] = 25'b01001000_11001100_00010100_1;
      patterns[18639] = 25'b01001000_11001101_00010101_1;
      patterns[18640] = 25'b01001000_11001110_00010110_1;
      patterns[18641] = 25'b01001000_11001111_00010111_1;
      patterns[18642] = 25'b01001000_11010000_00011000_1;
      patterns[18643] = 25'b01001000_11010001_00011001_1;
      patterns[18644] = 25'b01001000_11010010_00011010_1;
      patterns[18645] = 25'b01001000_11010011_00011011_1;
      patterns[18646] = 25'b01001000_11010100_00011100_1;
      patterns[18647] = 25'b01001000_11010101_00011101_1;
      patterns[18648] = 25'b01001000_11010110_00011110_1;
      patterns[18649] = 25'b01001000_11010111_00011111_1;
      patterns[18650] = 25'b01001000_11011000_00100000_1;
      patterns[18651] = 25'b01001000_11011001_00100001_1;
      patterns[18652] = 25'b01001000_11011010_00100010_1;
      patterns[18653] = 25'b01001000_11011011_00100011_1;
      patterns[18654] = 25'b01001000_11011100_00100100_1;
      patterns[18655] = 25'b01001000_11011101_00100101_1;
      patterns[18656] = 25'b01001000_11011110_00100110_1;
      patterns[18657] = 25'b01001000_11011111_00100111_1;
      patterns[18658] = 25'b01001000_11100000_00101000_1;
      patterns[18659] = 25'b01001000_11100001_00101001_1;
      patterns[18660] = 25'b01001000_11100010_00101010_1;
      patterns[18661] = 25'b01001000_11100011_00101011_1;
      patterns[18662] = 25'b01001000_11100100_00101100_1;
      patterns[18663] = 25'b01001000_11100101_00101101_1;
      patterns[18664] = 25'b01001000_11100110_00101110_1;
      patterns[18665] = 25'b01001000_11100111_00101111_1;
      patterns[18666] = 25'b01001000_11101000_00110000_1;
      patterns[18667] = 25'b01001000_11101001_00110001_1;
      patterns[18668] = 25'b01001000_11101010_00110010_1;
      patterns[18669] = 25'b01001000_11101011_00110011_1;
      patterns[18670] = 25'b01001000_11101100_00110100_1;
      patterns[18671] = 25'b01001000_11101101_00110101_1;
      patterns[18672] = 25'b01001000_11101110_00110110_1;
      patterns[18673] = 25'b01001000_11101111_00110111_1;
      patterns[18674] = 25'b01001000_11110000_00111000_1;
      patterns[18675] = 25'b01001000_11110001_00111001_1;
      patterns[18676] = 25'b01001000_11110010_00111010_1;
      patterns[18677] = 25'b01001000_11110011_00111011_1;
      patterns[18678] = 25'b01001000_11110100_00111100_1;
      patterns[18679] = 25'b01001000_11110101_00111101_1;
      patterns[18680] = 25'b01001000_11110110_00111110_1;
      patterns[18681] = 25'b01001000_11110111_00111111_1;
      patterns[18682] = 25'b01001000_11111000_01000000_1;
      patterns[18683] = 25'b01001000_11111001_01000001_1;
      patterns[18684] = 25'b01001000_11111010_01000010_1;
      patterns[18685] = 25'b01001000_11111011_01000011_1;
      patterns[18686] = 25'b01001000_11111100_01000100_1;
      patterns[18687] = 25'b01001000_11111101_01000101_1;
      patterns[18688] = 25'b01001000_11111110_01000110_1;
      patterns[18689] = 25'b01001000_11111111_01000111_1;
      patterns[18690] = 25'b01001001_00000000_01001001_0;
      patterns[18691] = 25'b01001001_00000001_01001010_0;
      patterns[18692] = 25'b01001001_00000010_01001011_0;
      patterns[18693] = 25'b01001001_00000011_01001100_0;
      patterns[18694] = 25'b01001001_00000100_01001101_0;
      patterns[18695] = 25'b01001001_00000101_01001110_0;
      patterns[18696] = 25'b01001001_00000110_01001111_0;
      patterns[18697] = 25'b01001001_00000111_01010000_0;
      patterns[18698] = 25'b01001001_00001000_01010001_0;
      patterns[18699] = 25'b01001001_00001001_01010010_0;
      patterns[18700] = 25'b01001001_00001010_01010011_0;
      patterns[18701] = 25'b01001001_00001011_01010100_0;
      patterns[18702] = 25'b01001001_00001100_01010101_0;
      patterns[18703] = 25'b01001001_00001101_01010110_0;
      patterns[18704] = 25'b01001001_00001110_01010111_0;
      patterns[18705] = 25'b01001001_00001111_01011000_0;
      patterns[18706] = 25'b01001001_00010000_01011001_0;
      patterns[18707] = 25'b01001001_00010001_01011010_0;
      patterns[18708] = 25'b01001001_00010010_01011011_0;
      patterns[18709] = 25'b01001001_00010011_01011100_0;
      patterns[18710] = 25'b01001001_00010100_01011101_0;
      patterns[18711] = 25'b01001001_00010101_01011110_0;
      patterns[18712] = 25'b01001001_00010110_01011111_0;
      patterns[18713] = 25'b01001001_00010111_01100000_0;
      patterns[18714] = 25'b01001001_00011000_01100001_0;
      patterns[18715] = 25'b01001001_00011001_01100010_0;
      patterns[18716] = 25'b01001001_00011010_01100011_0;
      patterns[18717] = 25'b01001001_00011011_01100100_0;
      patterns[18718] = 25'b01001001_00011100_01100101_0;
      patterns[18719] = 25'b01001001_00011101_01100110_0;
      patterns[18720] = 25'b01001001_00011110_01100111_0;
      patterns[18721] = 25'b01001001_00011111_01101000_0;
      patterns[18722] = 25'b01001001_00100000_01101001_0;
      patterns[18723] = 25'b01001001_00100001_01101010_0;
      patterns[18724] = 25'b01001001_00100010_01101011_0;
      patterns[18725] = 25'b01001001_00100011_01101100_0;
      patterns[18726] = 25'b01001001_00100100_01101101_0;
      patterns[18727] = 25'b01001001_00100101_01101110_0;
      patterns[18728] = 25'b01001001_00100110_01101111_0;
      patterns[18729] = 25'b01001001_00100111_01110000_0;
      patterns[18730] = 25'b01001001_00101000_01110001_0;
      patterns[18731] = 25'b01001001_00101001_01110010_0;
      patterns[18732] = 25'b01001001_00101010_01110011_0;
      patterns[18733] = 25'b01001001_00101011_01110100_0;
      patterns[18734] = 25'b01001001_00101100_01110101_0;
      patterns[18735] = 25'b01001001_00101101_01110110_0;
      patterns[18736] = 25'b01001001_00101110_01110111_0;
      patterns[18737] = 25'b01001001_00101111_01111000_0;
      patterns[18738] = 25'b01001001_00110000_01111001_0;
      patterns[18739] = 25'b01001001_00110001_01111010_0;
      patterns[18740] = 25'b01001001_00110010_01111011_0;
      patterns[18741] = 25'b01001001_00110011_01111100_0;
      patterns[18742] = 25'b01001001_00110100_01111101_0;
      patterns[18743] = 25'b01001001_00110101_01111110_0;
      patterns[18744] = 25'b01001001_00110110_01111111_0;
      patterns[18745] = 25'b01001001_00110111_10000000_0;
      patterns[18746] = 25'b01001001_00111000_10000001_0;
      patterns[18747] = 25'b01001001_00111001_10000010_0;
      patterns[18748] = 25'b01001001_00111010_10000011_0;
      patterns[18749] = 25'b01001001_00111011_10000100_0;
      patterns[18750] = 25'b01001001_00111100_10000101_0;
      patterns[18751] = 25'b01001001_00111101_10000110_0;
      patterns[18752] = 25'b01001001_00111110_10000111_0;
      patterns[18753] = 25'b01001001_00111111_10001000_0;
      patterns[18754] = 25'b01001001_01000000_10001001_0;
      patterns[18755] = 25'b01001001_01000001_10001010_0;
      patterns[18756] = 25'b01001001_01000010_10001011_0;
      patterns[18757] = 25'b01001001_01000011_10001100_0;
      patterns[18758] = 25'b01001001_01000100_10001101_0;
      patterns[18759] = 25'b01001001_01000101_10001110_0;
      patterns[18760] = 25'b01001001_01000110_10001111_0;
      patterns[18761] = 25'b01001001_01000111_10010000_0;
      patterns[18762] = 25'b01001001_01001000_10010001_0;
      patterns[18763] = 25'b01001001_01001001_10010010_0;
      patterns[18764] = 25'b01001001_01001010_10010011_0;
      patterns[18765] = 25'b01001001_01001011_10010100_0;
      patterns[18766] = 25'b01001001_01001100_10010101_0;
      patterns[18767] = 25'b01001001_01001101_10010110_0;
      patterns[18768] = 25'b01001001_01001110_10010111_0;
      patterns[18769] = 25'b01001001_01001111_10011000_0;
      patterns[18770] = 25'b01001001_01010000_10011001_0;
      patterns[18771] = 25'b01001001_01010001_10011010_0;
      patterns[18772] = 25'b01001001_01010010_10011011_0;
      patterns[18773] = 25'b01001001_01010011_10011100_0;
      patterns[18774] = 25'b01001001_01010100_10011101_0;
      patterns[18775] = 25'b01001001_01010101_10011110_0;
      patterns[18776] = 25'b01001001_01010110_10011111_0;
      patterns[18777] = 25'b01001001_01010111_10100000_0;
      patterns[18778] = 25'b01001001_01011000_10100001_0;
      patterns[18779] = 25'b01001001_01011001_10100010_0;
      patterns[18780] = 25'b01001001_01011010_10100011_0;
      patterns[18781] = 25'b01001001_01011011_10100100_0;
      patterns[18782] = 25'b01001001_01011100_10100101_0;
      patterns[18783] = 25'b01001001_01011101_10100110_0;
      patterns[18784] = 25'b01001001_01011110_10100111_0;
      patterns[18785] = 25'b01001001_01011111_10101000_0;
      patterns[18786] = 25'b01001001_01100000_10101001_0;
      patterns[18787] = 25'b01001001_01100001_10101010_0;
      patterns[18788] = 25'b01001001_01100010_10101011_0;
      patterns[18789] = 25'b01001001_01100011_10101100_0;
      patterns[18790] = 25'b01001001_01100100_10101101_0;
      patterns[18791] = 25'b01001001_01100101_10101110_0;
      patterns[18792] = 25'b01001001_01100110_10101111_0;
      patterns[18793] = 25'b01001001_01100111_10110000_0;
      patterns[18794] = 25'b01001001_01101000_10110001_0;
      patterns[18795] = 25'b01001001_01101001_10110010_0;
      patterns[18796] = 25'b01001001_01101010_10110011_0;
      patterns[18797] = 25'b01001001_01101011_10110100_0;
      patterns[18798] = 25'b01001001_01101100_10110101_0;
      patterns[18799] = 25'b01001001_01101101_10110110_0;
      patterns[18800] = 25'b01001001_01101110_10110111_0;
      patterns[18801] = 25'b01001001_01101111_10111000_0;
      patterns[18802] = 25'b01001001_01110000_10111001_0;
      patterns[18803] = 25'b01001001_01110001_10111010_0;
      patterns[18804] = 25'b01001001_01110010_10111011_0;
      patterns[18805] = 25'b01001001_01110011_10111100_0;
      patterns[18806] = 25'b01001001_01110100_10111101_0;
      patterns[18807] = 25'b01001001_01110101_10111110_0;
      patterns[18808] = 25'b01001001_01110110_10111111_0;
      patterns[18809] = 25'b01001001_01110111_11000000_0;
      patterns[18810] = 25'b01001001_01111000_11000001_0;
      patterns[18811] = 25'b01001001_01111001_11000010_0;
      patterns[18812] = 25'b01001001_01111010_11000011_0;
      patterns[18813] = 25'b01001001_01111011_11000100_0;
      patterns[18814] = 25'b01001001_01111100_11000101_0;
      patterns[18815] = 25'b01001001_01111101_11000110_0;
      patterns[18816] = 25'b01001001_01111110_11000111_0;
      patterns[18817] = 25'b01001001_01111111_11001000_0;
      patterns[18818] = 25'b01001001_10000000_11001001_0;
      patterns[18819] = 25'b01001001_10000001_11001010_0;
      patterns[18820] = 25'b01001001_10000010_11001011_0;
      patterns[18821] = 25'b01001001_10000011_11001100_0;
      patterns[18822] = 25'b01001001_10000100_11001101_0;
      patterns[18823] = 25'b01001001_10000101_11001110_0;
      patterns[18824] = 25'b01001001_10000110_11001111_0;
      patterns[18825] = 25'b01001001_10000111_11010000_0;
      patterns[18826] = 25'b01001001_10001000_11010001_0;
      patterns[18827] = 25'b01001001_10001001_11010010_0;
      patterns[18828] = 25'b01001001_10001010_11010011_0;
      patterns[18829] = 25'b01001001_10001011_11010100_0;
      patterns[18830] = 25'b01001001_10001100_11010101_0;
      patterns[18831] = 25'b01001001_10001101_11010110_0;
      patterns[18832] = 25'b01001001_10001110_11010111_0;
      patterns[18833] = 25'b01001001_10001111_11011000_0;
      patterns[18834] = 25'b01001001_10010000_11011001_0;
      patterns[18835] = 25'b01001001_10010001_11011010_0;
      patterns[18836] = 25'b01001001_10010010_11011011_0;
      patterns[18837] = 25'b01001001_10010011_11011100_0;
      patterns[18838] = 25'b01001001_10010100_11011101_0;
      patterns[18839] = 25'b01001001_10010101_11011110_0;
      patterns[18840] = 25'b01001001_10010110_11011111_0;
      patterns[18841] = 25'b01001001_10010111_11100000_0;
      patterns[18842] = 25'b01001001_10011000_11100001_0;
      patterns[18843] = 25'b01001001_10011001_11100010_0;
      patterns[18844] = 25'b01001001_10011010_11100011_0;
      patterns[18845] = 25'b01001001_10011011_11100100_0;
      patterns[18846] = 25'b01001001_10011100_11100101_0;
      patterns[18847] = 25'b01001001_10011101_11100110_0;
      patterns[18848] = 25'b01001001_10011110_11100111_0;
      patterns[18849] = 25'b01001001_10011111_11101000_0;
      patterns[18850] = 25'b01001001_10100000_11101001_0;
      patterns[18851] = 25'b01001001_10100001_11101010_0;
      patterns[18852] = 25'b01001001_10100010_11101011_0;
      patterns[18853] = 25'b01001001_10100011_11101100_0;
      patterns[18854] = 25'b01001001_10100100_11101101_0;
      patterns[18855] = 25'b01001001_10100101_11101110_0;
      patterns[18856] = 25'b01001001_10100110_11101111_0;
      patterns[18857] = 25'b01001001_10100111_11110000_0;
      patterns[18858] = 25'b01001001_10101000_11110001_0;
      patterns[18859] = 25'b01001001_10101001_11110010_0;
      patterns[18860] = 25'b01001001_10101010_11110011_0;
      patterns[18861] = 25'b01001001_10101011_11110100_0;
      patterns[18862] = 25'b01001001_10101100_11110101_0;
      patterns[18863] = 25'b01001001_10101101_11110110_0;
      patterns[18864] = 25'b01001001_10101110_11110111_0;
      patterns[18865] = 25'b01001001_10101111_11111000_0;
      patterns[18866] = 25'b01001001_10110000_11111001_0;
      patterns[18867] = 25'b01001001_10110001_11111010_0;
      patterns[18868] = 25'b01001001_10110010_11111011_0;
      patterns[18869] = 25'b01001001_10110011_11111100_0;
      patterns[18870] = 25'b01001001_10110100_11111101_0;
      patterns[18871] = 25'b01001001_10110101_11111110_0;
      patterns[18872] = 25'b01001001_10110110_11111111_0;
      patterns[18873] = 25'b01001001_10110111_00000000_1;
      patterns[18874] = 25'b01001001_10111000_00000001_1;
      patterns[18875] = 25'b01001001_10111001_00000010_1;
      patterns[18876] = 25'b01001001_10111010_00000011_1;
      patterns[18877] = 25'b01001001_10111011_00000100_1;
      patterns[18878] = 25'b01001001_10111100_00000101_1;
      patterns[18879] = 25'b01001001_10111101_00000110_1;
      patterns[18880] = 25'b01001001_10111110_00000111_1;
      patterns[18881] = 25'b01001001_10111111_00001000_1;
      patterns[18882] = 25'b01001001_11000000_00001001_1;
      patterns[18883] = 25'b01001001_11000001_00001010_1;
      patterns[18884] = 25'b01001001_11000010_00001011_1;
      patterns[18885] = 25'b01001001_11000011_00001100_1;
      patterns[18886] = 25'b01001001_11000100_00001101_1;
      patterns[18887] = 25'b01001001_11000101_00001110_1;
      patterns[18888] = 25'b01001001_11000110_00001111_1;
      patterns[18889] = 25'b01001001_11000111_00010000_1;
      patterns[18890] = 25'b01001001_11001000_00010001_1;
      patterns[18891] = 25'b01001001_11001001_00010010_1;
      patterns[18892] = 25'b01001001_11001010_00010011_1;
      patterns[18893] = 25'b01001001_11001011_00010100_1;
      patterns[18894] = 25'b01001001_11001100_00010101_1;
      patterns[18895] = 25'b01001001_11001101_00010110_1;
      patterns[18896] = 25'b01001001_11001110_00010111_1;
      patterns[18897] = 25'b01001001_11001111_00011000_1;
      patterns[18898] = 25'b01001001_11010000_00011001_1;
      patterns[18899] = 25'b01001001_11010001_00011010_1;
      patterns[18900] = 25'b01001001_11010010_00011011_1;
      patterns[18901] = 25'b01001001_11010011_00011100_1;
      patterns[18902] = 25'b01001001_11010100_00011101_1;
      patterns[18903] = 25'b01001001_11010101_00011110_1;
      patterns[18904] = 25'b01001001_11010110_00011111_1;
      patterns[18905] = 25'b01001001_11010111_00100000_1;
      patterns[18906] = 25'b01001001_11011000_00100001_1;
      patterns[18907] = 25'b01001001_11011001_00100010_1;
      patterns[18908] = 25'b01001001_11011010_00100011_1;
      patterns[18909] = 25'b01001001_11011011_00100100_1;
      patterns[18910] = 25'b01001001_11011100_00100101_1;
      patterns[18911] = 25'b01001001_11011101_00100110_1;
      patterns[18912] = 25'b01001001_11011110_00100111_1;
      patterns[18913] = 25'b01001001_11011111_00101000_1;
      patterns[18914] = 25'b01001001_11100000_00101001_1;
      patterns[18915] = 25'b01001001_11100001_00101010_1;
      patterns[18916] = 25'b01001001_11100010_00101011_1;
      patterns[18917] = 25'b01001001_11100011_00101100_1;
      patterns[18918] = 25'b01001001_11100100_00101101_1;
      patterns[18919] = 25'b01001001_11100101_00101110_1;
      patterns[18920] = 25'b01001001_11100110_00101111_1;
      patterns[18921] = 25'b01001001_11100111_00110000_1;
      patterns[18922] = 25'b01001001_11101000_00110001_1;
      patterns[18923] = 25'b01001001_11101001_00110010_1;
      patterns[18924] = 25'b01001001_11101010_00110011_1;
      patterns[18925] = 25'b01001001_11101011_00110100_1;
      patterns[18926] = 25'b01001001_11101100_00110101_1;
      patterns[18927] = 25'b01001001_11101101_00110110_1;
      patterns[18928] = 25'b01001001_11101110_00110111_1;
      patterns[18929] = 25'b01001001_11101111_00111000_1;
      patterns[18930] = 25'b01001001_11110000_00111001_1;
      patterns[18931] = 25'b01001001_11110001_00111010_1;
      patterns[18932] = 25'b01001001_11110010_00111011_1;
      patterns[18933] = 25'b01001001_11110011_00111100_1;
      patterns[18934] = 25'b01001001_11110100_00111101_1;
      patterns[18935] = 25'b01001001_11110101_00111110_1;
      patterns[18936] = 25'b01001001_11110110_00111111_1;
      patterns[18937] = 25'b01001001_11110111_01000000_1;
      patterns[18938] = 25'b01001001_11111000_01000001_1;
      patterns[18939] = 25'b01001001_11111001_01000010_1;
      patterns[18940] = 25'b01001001_11111010_01000011_1;
      patterns[18941] = 25'b01001001_11111011_01000100_1;
      patterns[18942] = 25'b01001001_11111100_01000101_1;
      patterns[18943] = 25'b01001001_11111101_01000110_1;
      patterns[18944] = 25'b01001001_11111110_01000111_1;
      patterns[18945] = 25'b01001001_11111111_01001000_1;
      patterns[18946] = 25'b01001010_00000000_01001010_0;
      patterns[18947] = 25'b01001010_00000001_01001011_0;
      patterns[18948] = 25'b01001010_00000010_01001100_0;
      patterns[18949] = 25'b01001010_00000011_01001101_0;
      patterns[18950] = 25'b01001010_00000100_01001110_0;
      patterns[18951] = 25'b01001010_00000101_01001111_0;
      patterns[18952] = 25'b01001010_00000110_01010000_0;
      patterns[18953] = 25'b01001010_00000111_01010001_0;
      patterns[18954] = 25'b01001010_00001000_01010010_0;
      patterns[18955] = 25'b01001010_00001001_01010011_0;
      patterns[18956] = 25'b01001010_00001010_01010100_0;
      patterns[18957] = 25'b01001010_00001011_01010101_0;
      patterns[18958] = 25'b01001010_00001100_01010110_0;
      patterns[18959] = 25'b01001010_00001101_01010111_0;
      patterns[18960] = 25'b01001010_00001110_01011000_0;
      patterns[18961] = 25'b01001010_00001111_01011001_0;
      patterns[18962] = 25'b01001010_00010000_01011010_0;
      patterns[18963] = 25'b01001010_00010001_01011011_0;
      patterns[18964] = 25'b01001010_00010010_01011100_0;
      patterns[18965] = 25'b01001010_00010011_01011101_0;
      patterns[18966] = 25'b01001010_00010100_01011110_0;
      patterns[18967] = 25'b01001010_00010101_01011111_0;
      patterns[18968] = 25'b01001010_00010110_01100000_0;
      patterns[18969] = 25'b01001010_00010111_01100001_0;
      patterns[18970] = 25'b01001010_00011000_01100010_0;
      patterns[18971] = 25'b01001010_00011001_01100011_0;
      patterns[18972] = 25'b01001010_00011010_01100100_0;
      patterns[18973] = 25'b01001010_00011011_01100101_0;
      patterns[18974] = 25'b01001010_00011100_01100110_0;
      patterns[18975] = 25'b01001010_00011101_01100111_0;
      patterns[18976] = 25'b01001010_00011110_01101000_0;
      patterns[18977] = 25'b01001010_00011111_01101001_0;
      patterns[18978] = 25'b01001010_00100000_01101010_0;
      patterns[18979] = 25'b01001010_00100001_01101011_0;
      patterns[18980] = 25'b01001010_00100010_01101100_0;
      patterns[18981] = 25'b01001010_00100011_01101101_0;
      patterns[18982] = 25'b01001010_00100100_01101110_0;
      patterns[18983] = 25'b01001010_00100101_01101111_0;
      patterns[18984] = 25'b01001010_00100110_01110000_0;
      patterns[18985] = 25'b01001010_00100111_01110001_0;
      patterns[18986] = 25'b01001010_00101000_01110010_0;
      patterns[18987] = 25'b01001010_00101001_01110011_0;
      patterns[18988] = 25'b01001010_00101010_01110100_0;
      patterns[18989] = 25'b01001010_00101011_01110101_0;
      patterns[18990] = 25'b01001010_00101100_01110110_0;
      patterns[18991] = 25'b01001010_00101101_01110111_0;
      patterns[18992] = 25'b01001010_00101110_01111000_0;
      patterns[18993] = 25'b01001010_00101111_01111001_0;
      patterns[18994] = 25'b01001010_00110000_01111010_0;
      patterns[18995] = 25'b01001010_00110001_01111011_0;
      patterns[18996] = 25'b01001010_00110010_01111100_0;
      patterns[18997] = 25'b01001010_00110011_01111101_0;
      patterns[18998] = 25'b01001010_00110100_01111110_0;
      patterns[18999] = 25'b01001010_00110101_01111111_0;
      patterns[19000] = 25'b01001010_00110110_10000000_0;
      patterns[19001] = 25'b01001010_00110111_10000001_0;
      patterns[19002] = 25'b01001010_00111000_10000010_0;
      patterns[19003] = 25'b01001010_00111001_10000011_0;
      patterns[19004] = 25'b01001010_00111010_10000100_0;
      patterns[19005] = 25'b01001010_00111011_10000101_0;
      patterns[19006] = 25'b01001010_00111100_10000110_0;
      patterns[19007] = 25'b01001010_00111101_10000111_0;
      patterns[19008] = 25'b01001010_00111110_10001000_0;
      patterns[19009] = 25'b01001010_00111111_10001001_0;
      patterns[19010] = 25'b01001010_01000000_10001010_0;
      patterns[19011] = 25'b01001010_01000001_10001011_0;
      patterns[19012] = 25'b01001010_01000010_10001100_0;
      patterns[19013] = 25'b01001010_01000011_10001101_0;
      patterns[19014] = 25'b01001010_01000100_10001110_0;
      patterns[19015] = 25'b01001010_01000101_10001111_0;
      patterns[19016] = 25'b01001010_01000110_10010000_0;
      patterns[19017] = 25'b01001010_01000111_10010001_0;
      patterns[19018] = 25'b01001010_01001000_10010010_0;
      patterns[19019] = 25'b01001010_01001001_10010011_0;
      patterns[19020] = 25'b01001010_01001010_10010100_0;
      patterns[19021] = 25'b01001010_01001011_10010101_0;
      patterns[19022] = 25'b01001010_01001100_10010110_0;
      patterns[19023] = 25'b01001010_01001101_10010111_0;
      patterns[19024] = 25'b01001010_01001110_10011000_0;
      patterns[19025] = 25'b01001010_01001111_10011001_0;
      patterns[19026] = 25'b01001010_01010000_10011010_0;
      patterns[19027] = 25'b01001010_01010001_10011011_0;
      patterns[19028] = 25'b01001010_01010010_10011100_0;
      patterns[19029] = 25'b01001010_01010011_10011101_0;
      patterns[19030] = 25'b01001010_01010100_10011110_0;
      patterns[19031] = 25'b01001010_01010101_10011111_0;
      patterns[19032] = 25'b01001010_01010110_10100000_0;
      patterns[19033] = 25'b01001010_01010111_10100001_0;
      patterns[19034] = 25'b01001010_01011000_10100010_0;
      patterns[19035] = 25'b01001010_01011001_10100011_0;
      patterns[19036] = 25'b01001010_01011010_10100100_0;
      patterns[19037] = 25'b01001010_01011011_10100101_0;
      patterns[19038] = 25'b01001010_01011100_10100110_0;
      patterns[19039] = 25'b01001010_01011101_10100111_0;
      patterns[19040] = 25'b01001010_01011110_10101000_0;
      patterns[19041] = 25'b01001010_01011111_10101001_0;
      patterns[19042] = 25'b01001010_01100000_10101010_0;
      patterns[19043] = 25'b01001010_01100001_10101011_0;
      patterns[19044] = 25'b01001010_01100010_10101100_0;
      patterns[19045] = 25'b01001010_01100011_10101101_0;
      patterns[19046] = 25'b01001010_01100100_10101110_0;
      patterns[19047] = 25'b01001010_01100101_10101111_0;
      patterns[19048] = 25'b01001010_01100110_10110000_0;
      patterns[19049] = 25'b01001010_01100111_10110001_0;
      patterns[19050] = 25'b01001010_01101000_10110010_0;
      patterns[19051] = 25'b01001010_01101001_10110011_0;
      patterns[19052] = 25'b01001010_01101010_10110100_0;
      patterns[19053] = 25'b01001010_01101011_10110101_0;
      patterns[19054] = 25'b01001010_01101100_10110110_0;
      patterns[19055] = 25'b01001010_01101101_10110111_0;
      patterns[19056] = 25'b01001010_01101110_10111000_0;
      patterns[19057] = 25'b01001010_01101111_10111001_0;
      patterns[19058] = 25'b01001010_01110000_10111010_0;
      patterns[19059] = 25'b01001010_01110001_10111011_0;
      patterns[19060] = 25'b01001010_01110010_10111100_0;
      patterns[19061] = 25'b01001010_01110011_10111101_0;
      patterns[19062] = 25'b01001010_01110100_10111110_0;
      patterns[19063] = 25'b01001010_01110101_10111111_0;
      patterns[19064] = 25'b01001010_01110110_11000000_0;
      patterns[19065] = 25'b01001010_01110111_11000001_0;
      patterns[19066] = 25'b01001010_01111000_11000010_0;
      patterns[19067] = 25'b01001010_01111001_11000011_0;
      patterns[19068] = 25'b01001010_01111010_11000100_0;
      patterns[19069] = 25'b01001010_01111011_11000101_0;
      patterns[19070] = 25'b01001010_01111100_11000110_0;
      patterns[19071] = 25'b01001010_01111101_11000111_0;
      patterns[19072] = 25'b01001010_01111110_11001000_0;
      patterns[19073] = 25'b01001010_01111111_11001001_0;
      patterns[19074] = 25'b01001010_10000000_11001010_0;
      patterns[19075] = 25'b01001010_10000001_11001011_0;
      patterns[19076] = 25'b01001010_10000010_11001100_0;
      patterns[19077] = 25'b01001010_10000011_11001101_0;
      patterns[19078] = 25'b01001010_10000100_11001110_0;
      patterns[19079] = 25'b01001010_10000101_11001111_0;
      patterns[19080] = 25'b01001010_10000110_11010000_0;
      patterns[19081] = 25'b01001010_10000111_11010001_0;
      patterns[19082] = 25'b01001010_10001000_11010010_0;
      patterns[19083] = 25'b01001010_10001001_11010011_0;
      patterns[19084] = 25'b01001010_10001010_11010100_0;
      patterns[19085] = 25'b01001010_10001011_11010101_0;
      patterns[19086] = 25'b01001010_10001100_11010110_0;
      patterns[19087] = 25'b01001010_10001101_11010111_0;
      patterns[19088] = 25'b01001010_10001110_11011000_0;
      patterns[19089] = 25'b01001010_10001111_11011001_0;
      patterns[19090] = 25'b01001010_10010000_11011010_0;
      patterns[19091] = 25'b01001010_10010001_11011011_0;
      patterns[19092] = 25'b01001010_10010010_11011100_0;
      patterns[19093] = 25'b01001010_10010011_11011101_0;
      patterns[19094] = 25'b01001010_10010100_11011110_0;
      patterns[19095] = 25'b01001010_10010101_11011111_0;
      patterns[19096] = 25'b01001010_10010110_11100000_0;
      patterns[19097] = 25'b01001010_10010111_11100001_0;
      patterns[19098] = 25'b01001010_10011000_11100010_0;
      patterns[19099] = 25'b01001010_10011001_11100011_0;
      patterns[19100] = 25'b01001010_10011010_11100100_0;
      patterns[19101] = 25'b01001010_10011011_11100101_0;
      patterns[19102] = 25'b01001010_10011100_11100110_0;
      patterns[19103] = 25'b01001010_10011101_11100111_0;
      patterns[19104] = 25'b01001010_10011110_11101000_0;
      patterns[19105] = 25'b01001010_10011111_11101001_0;
      patterns[19106] = 25'b01001010_10100000_11101010_0;
      patterns[19107] = 25'b01001010_10100001_11101011_0;
      patterns[19108] = 25'b01001010_10100010_11101100_0;
      patterns[19109] = 25'b01001010_10100011_11101101_0;
      patterns[19110] = 25'b01001010_10100100_11101110_0;
      patterns[19111] = 25'b01001010_10100101_11101111_0;
      patterns[19112] = 25'b01001010_10100110_11110000_0;
      patterns[19113] = 25'b01001010_10100111_11110001_0;
      patterns[19114] = 25'b01001010_10101000_11110010_0;
      patterns[19115] = 25'b01001010_10101001_11110011_0;
      patterns[19116] = 25'b01001010_10101010_11110100_0;
      patterns[19117] = 25'b01001010_10101011_11110101_0;
      patterns[19118] = 25'b01001010_10101100_11110110_0;
      patterns[19119] = 25'b01001010_10101101_11110111_0;
      patterns[19120] = 25'b01001010_10101110_11111000_0;
      patterns[19121] = 25'b01001010_10101111_11111001_0;
      patterns[19122] = 25'b01001010_10110000_11111010_0;
      patterns[19123] = 25'b01001010_10110001_11111011_0;
      patterns[19124] = 25'b01001010_10110010_11111100_0;
      patterns[19125] = 25'b01001010_10110011_11111101_0;
      patterns[19126] = 25'b01001010_10110100_11111110_0;
      patterns[19127] = 25'b01001010_10110101_11111111_0;
      patterns[19128] = 25'b01001010_10110110_00000000_1;
      patterns[19129] = 25'b01001010_10110111_00000001_1;
      patterns[19130] = 25'b01001010_10111000_00000010_1;
      patterns[19131] = 25'b01001010_10111001_00000011_1;
      patterns[19132] = 25'b01001010_10111010_00000100_1;
      patterns[19133] = 25'b01001010_10111011_00000101_1;
      patterns[19134] = 25'b01001010_10111100_00000110_1;
      patterns[19135] = 25'b01001010_10111101_00000111_1;
      patterns[19136] = 25'b01001010_10111110_00001000_1;
      patterns[19137] = 25'b01001010_10111111_00001001_1;
      patterns[19138] = 25'b01001010_11000000_00001010_1;
      patterns[19139] = 25'b01001010_11000001_00001011_1;
      patterns[19140] = 25'b01001010_11000010_00001100_1;
      patterns[19141] = 25'b01001010_11000011_00001101_1;
      patterns[19142] = 25'b01001010_11000100_00001110_1;
      patterns[19143] = 25'b01001010_11000101_00001111_1;
      patterns[19144] = 25'b01001010_11000110_00010000_1;
      patterns[19145] = 25'b01001010_11000111_00010001_1;
      patterns[19146] = 25'b01001010_11001000_00010010_1;
      patterns[19147] = 25'b01001010_11001001_00010011_1;
      patterns[19148] = 25'b01001010_11001010_00010100_1;
      patterns[19149] = 25'b01001010_11001011_00010101_1;
      patterns[19150] = 25'b01001010_11001100_00010110_1;
      patterns[19151] = 25'b01001010_11001101_00010111_1;
      patterns[19152] = 25'b01001010_11001110_00011000_1;
      patterns[19153] = 25'b01001010_11001111_00011001_1;
      patterns[19154] = 25'b01001010_11010000_00011010_1;
      patterns[19155] = 25'b01001010_11010001_00011011_1;
      patterns[19156] = 25'b01001010_11010010_00011100_1;
      patterns[19157] = 25'b01001010_11010011_00011101_1;
      patterns[19158] = 25'b01001010_11010100_00011110_1;
      patterns[19159] = 25'b01001010_11010101_00011111_1;
      patterns[19160] = 25'b01001010_11010110_00100000_1;
      patterns[19161] = 25'b01001010_11010111_00100001_1;
      patterns[19162] = 25'b01001010_11011000_00100010_1;
      patterns[19163] = 25'b01001010_11011001_00100011_1;
      patterns[19164] = 25'b01001010_11011010_00100100_1;
      patterns[19165] = 25'b01001010_11011011_00100101_1;
      patterns[19166] = 25'b01001010_11011100_00100110_1;
      patterns[19167] = 25'b01001010_11011101_00100111_1;
      patterns[19168] = 25'b01001010_11011110_00101000_1;
      patterns[19169] = 25'b01001010_11011111_00101001_1;
      patterns[19170] = 25'b01001010_11100000_00101010_1;
      patterns[19171] = 25'b01001010_11100001_00101011_1;
      patterns[19172] = 25'b01001010_11100010_00101100_1;
      patterns[19173] = 25'b01001010_11100011_00101101_1;
      patterns[19174] = 25'b01001010_11100100_00101110_1;
      patterns[19175] = 25'b01001010_11100101_00101111_1;
      patterns[19176] = 25'b01001010_11100110_00110000_1;
      patterns[19177] = 25'b01001010_11100111_00110001_1;
      patterns[19178] = 25'b01001010_11101000_00110010_1;
      patterns[19179] = 25'b01001010_11101001_00110011_1;
      patterns[19180] = 25'b01001010_11101010_00110100_1;
      patterns[19181] = 25'b01001010_11101011_00110101_1;
      patterns[19182] = 25'b01001010_11101100_00110110_1;
      patterns[19183] = 25'b01001010_11101101_00110111_1;
      patterns[19184] = 25'b01001010_11101110_00111000_1;
      patterns[19185] = 25'b01001010_11101111_00111001_1;
      patterns[19186] = 25'b01001010_11110000_00111010_1;
      patterns[19187] = 25'b01001010_11110001_00111011_1;
      patterns[19188] = 25'b01001010_11110010_00111100_1;
      patterns[19189] = 25'b01001010_11110011_00111101_1;
      patterns[19190] = 25'b01001010_11110100_00111110_1;
      patterns[19191] = 25'b01001010_11110101_00111111_1;
      patterns[19192] = 25'b01001010_11110110_01000000_1;
      patterns[19193] = 25'b01001010_11110111_01000001_1;
      patterns[19194] = 25'b01001010_11111000_01000010_1;
      patterns[19195] = 25'b01001010_11111001_01000011_1;
      patterns[19196] = 25'b01001010_11111010_01000100_1;
      patterns[19197] = 25'b01001010_11111011_01000101_1;
      patterns[19198] = 25'b01001010_11111100_01000110_1;
      patterns[19199] = 25'b01001010_11111101_01000111_1;
      patterns[19200] = 25'b01001010_11111110_01001000_1;
      patterns[19201] = 25'b01001010_11111111_01001001_1;
      patterns[19202] = 25'b01001011_00000000_01001011_0;
      patterns[19203] = 25'b01001011_00000001_01001100_0;
      patterns[19204] = 25'b01001011_00000010_01001101_0;
      patterns[19205] = 25'b01001011_00000011_01001110_0;
      patterns[19206] = 25'b01001011_00000100_01001111_0;
      patterns[19207] = 25'b01001011_00000101_01010000_0;
      patterns[19208] = 25'b01001011_00000110_01010001_0;
      patterns[19209] = 25'b01001011_00000111_01010010_0;
      patterns[19210] = 25'b01001011_00001000_01010011_0;
      patterns[19211] = 25'b01001011_00001001_01010100_0;
      patterns[19212] = 25'b01001011_00001010_01010101_0;
      patterns[19213] = 25'b01001011_00001011_01010110_0;
      patterns[19214] = 25'b01001011_00001100_01010111_0;
      patterns[19215] = 25'b01001011_00001101_01011000_0;
      patterns[19216] = 25'b01001011_00001110_01011001_0;
      patterns[19217] = 25'b01001011_00001111_01011010_0;
      patterns[19218] = 25'b01001011_00010000_01011011_0;
      patterns[19219] = 25'b01001011_00010001_01011100_0;
      patterns[19220] = 25'b01001011_00010010_01011101_0;
      patterns[19221] = 25'b01001011_00010011_01011110_0;
      patterns[19222] = 25'b01001011_00010100_01011111_0;
      patterns[19223] = 25'b01001011_00010101_01100000_0;
      patterns[19224] = 25'b01001011_00010110_01100001_0;
      patterns[19225] = 25'b01001011_00010111_01100010_0;
      patterns[19226] = 25'b01001011_00011000_01100011_0;
      patterns[19227] = 25'b01001011_00011001_01100100_0;
      patterns[19228] = 25'b01001011_00011010_01100101_0;
      patterns[19229] = 25'b01001011_00011011_01100110_0;
      patterns[19230] = 25'b01001011_00011100_01100111_0;
      patterns[19231] = 25'b01001011_00011101_01101000_0;
      patterns[19232] = 25'b01001011_00011110_01101001_0;
      patterns[19233] = 25'b01001011_00011111_01101010_0;
      patterns[19234] = 25'b01001011_00100000_01101011_0;
      patterns[19235] = 25'b01001011_00100001_01101100_0;
      patterns[19236] = 25'b01001011_00100010_01101101_0;
      patterns[19237] = 25'b01001011_00100011_01101110_0;
      patterns[19238] = 25'b01001011_00100100_01101111_0;
      patterns[19239] = 25'b01001011_00100101_01110000_0;
      patterns[19240] = 25'b01001011_00100110_01110001_0;
      patterns[19241] = 25'b01001011_00100111_01110010_0;
      patterns[19242] = 25'b01001011_00101000_01110011_0;
      patterns[19243] = 25'b01001011_00101001_01110100_0;
      patterns[19244] = 25'b01001011_00101010_01110101_0;
      patterns[19245] = 25'b01001011_00101011_01110110_0;
      patterns[19246] = 25'b01001011_00101100_01110111_0;
      patterns[19247] = 25'b01001011_00101101_01111000_0;
      patterns[19248] = 25'b01001011_00101110_01111001_0;
      patterns[19249] = 25'b01001011_00101111_01111010_0;
      patterns[19250] = 25'b01001011_00110000_01111011_0;
      patterns[19251] = 25'b01001011_00110001_01111100_0;
      patterns[19252] = 25'b01001011_00110010_01111101_0;
      patterns[19253] = 25'b01001011_00110011_01111110_0;
      patterns[19254] = 25'b01001011_00110100_01111111_0;
      patterns[19255] = 25'b01001011_00110101_10000000_0;
      patterns[19256] = 25'b01001011_00110110_10000001_0;
      patterns[19257] = 25'b01001011_00110111_10000010_0;
      patterns[19258] = 25'b01001011_00111000_10000011_0;
      patterns[19259] = 25'b01001011_00111001_10000100_0;
      patterns[19260] = 25'b01001011_00111010_10000101_0;
      patterns[19261] = 25'b01001011_00111011_10000110_0;
      patterns[19262] = 25'b01001011_00111100_10000111_0;
      patterns[19263] = 25'b01001011_00111101_10001000_0;
      patterns[19264] = 25'b01001011_00111110_10001001_0;
      patterns[19265] = 25'b01001011_00111111_10001010_0;
      patterns[19266] = 25'b01001011_01000000_10001011_0;
      patterns[19267] = 25'b01001011_01000001_10001100_0;
      patterns[19268] = 25'b01001011_01000010_10001101_0;
      patterns[19269] = 25'b01001011_01000011_10001110_0;
      patterns[19270] = 25'b01001011_01000100_10001111_0;
      patterns[19271] = 25'b01001011_01000101_10010000_0;
      patterns[19272] = 25'b01001011_01000110_10010001_0;
      patterns[19273] = 25'b01001011_01000111_10010010_0;
      patterns[19274] = 25'b01001011_01001000_10010011_0;
      patterns[19275] = 25'b01001011_01001001_10010100_0;
      patterns[19276] = 25'b01001011_01001010_10010101_0;
      patterns[19277] = 25'b01001011_01001011_10010110_0;
      patterns[19278] = 25'b01001011_01001100_10010111_0;
      patterns[19279] = 25'b01001011_01001101_10011000_0;
      patterns[19280] = 25'b01001011_01001110_10011001_0;
      patterns[19281] = 25'b01001011_01001111_10011010_0;
      patterns[19282] = 25'b01001011_01010000_10011011_0;
      patterns[19283] = 25'b01001011_01010001_10011100_0;
      patterns[19284] = 25'b01001011_01010010_10011101_0;
      patterns[19285] = 25'b01001011_01010011_10011110_0;
      patterns[19286] = 25'b01001011_01010100_10011111_0;
      patterns[19287] = 25'b01001011_01010101_10100000_0;
      patterns[19288] = 25'b01001011_01010110_10100001_0;
      patterns[19289] = 25'b01001011_01010111_10100010_0;
      patterns[19290] = 25'b01001011_01011000_10100011_0;
      patterns[19291] = 25'b01001011_01011001_10100100_0;
      patterns[19292] = 25'b01001011_01011010_10100101_0;
      patterns[19293] = 25'b01001011_01011011_10100110_0;
      patterns[19294] = 25'b01001011_01011100_10100111_0;
      patterns[19295] = 25'b01001011_01011101_10101000_0;
      patterns[19296] = 25'b01001011_01011110_10101001_0;
      patterns[19297] = 25'b01001011_01011111_10101010_0;
      patterns[19298] = 25'b01001011_01100000_10101011_0;
      patterns[19299] = 25'b01001011_01100001_10101100_0;
      patterns[19300] = 25'b01001011_01100010_10101101_0;
      patterns[19301] = 25'b01001011_01100011_10101110_0;
      patterns[19302] = 25'b01001011_01100100_10101111_0;
      patterns[19303] = 25'b01001011_01100101_10110000_0;
      patterns[19304] = 25'b01001011_01100110_10110001_0;
      patterns[19305] = 25'b01001011_01100111_10110010_0;
      patterns[19306] = 25'b01001011_01101000_10110011_0;
      patterns[19307] = 25'b01001011_01101001_10110100_0;
      patterns[19308] = 25'b01001011_01101010_10110101_0;
      patterns[19309] = 25'b01001011_01101011_10110110_0;
      patterns[19310] = 25'b01001011_01101100_10110111_0;
      patterns[19311] = 25'b01001011_01101101_10111000_0;
      patterns[19312] = 25'b01001011_01101110_10111001_0;
      patterns[19313] = 25'b01001011_01101111_10111010_0;
      patterns[19314] = 25'b01001011_01110000_10111011_0;
      patterns[19315] = 25'b01001011_01110001_10111100_0;
      patterns[19316] = 25'b01001011_01110010_10111101_0;
      patterns[19317] = 25'b01001011_01110011_10111110_0;
      patterns[19318] = 25'b01001011_01110100_10111111_0;
      patterns[19319] = 25'b01001011_01110101_11000000_0;
      patterns[19320] = 25'b01001011_01110110_11000001_0;
      patterns[19321] = 25'b01001011_01110111_11000010_0;
      patterns[19322] = 25'b01001011_01111000_11000011_0;
      patterns[19323] = 25'b01001011_01111001_11000100_0;
      patterns[19324] = 25'b01001011_01111010_11000101_0;
      patterns[19325] = 25'b01001011_01111011_11000110_0;
      patterns[19326] = 25'b01001011_01111100_11000111_0;
      patterns[19327] = 25'b01001011_01111101_11001000_0;
      patterns[19328] = 25'b01001011_01111110_11001001_0;
      patterns[19329] = 25'b01001011_01111111_11001010_0;
      patterns[19330] = 25'b01001011_10000000_11001011_0;
      patterns[19331] = 25'b01001011_10000001_11001100_0;
      patterns[19332] = 25'b01001011_10000010_11001101_0;
      patterns[19333] = 25'b01001011_10000011_11001110_0;
      patterns[19334] = 25'b01001011_10000100_11001111_0;
      patterns[19335] = 25'b01001011_10000101_11010000_0;
      patterns[19336] = 25'b01001011_10000110_11010001_0;
      patterns[19337] = 25'b01001011_10000111_11010010_0;
      patterns[19338] = 25'b01001011_10001000_11010011_0;
      patterns[19339] = 25'b01001011_10001001_11010100_0;
      patterns[19340] = 25'b01001011_10001010_11010101_0;
      patterns[19341] = 25'b01001011_10001011_11010110_0;
      patterns[19342] = 25'b01001011_10001100_11010111_0;
      patterns[19343] = 25'b01001011_10001101_11011000_0;
      patterns[19344] = 25'b01001011_10001110_11011001_0;
      patterns[19345] = 25'b01001011_10001111_11011010_0;
      patterns[19346] = 25'b01001011_10010000_11011011_0;
      patterns[19347] = 25'b01001011_10010001_11011100_0;
      patterns[19348] = 25'b01001011_10010010_11011101_0;
      patterns[19349] = 25'b01001011_10010011_11011110_0;
      patterns[19350] = 25'b01001011_10010100_11011111_0;
      patterns[19351] = 25'b01001011_10010101_11100000_0;
      patterns[19352] = 25'b01001011_10010110_11100001_0;
      patterns[19353] = 25'b01001011_10010111_11100010_0;
      patterns[19354] = 25'b01001011_10011000_11100011_0;
      patterns[19355] = 25'b01001011_10011001_11100100_0;
      patterns[19356] = 25'b01001011_10011010_11100101_0;
      patterns[19357] = 25'b01001011_10011011_11100110_0;
      patterns[19358] = 25'b01001011_10011100_11100111_0;
      patterns[19359] = 25'b01001011_10011101_11101000_0;
      patterns[19360] = 25'b01001011_10011110_11101001_0;
      patterns[19361] = 25'b01001011_10011111_11101010_0;
      patterns[19362] = 25'b01001011_10100000_11101011_0;
      patterns[19363] = 25'b01001011_10100001_11101100_0;
      patterns[19364] = 25'b01001011_10100010_11101101_0;
      patterns[19365] = 25'b01001011_10100011_11101110_0;
      patterns[19366] = 25'b01001011_10100100_11101111_0;
      patterns[19367] = 25'b01001011_10100101_11110000_0;
      patterns[19368] = 25'b01001011_10100110_11110001_0;
      patterns[19369] = 25'b01001011_10100111_11110010_0;
      patterns[19370] = 25'b01001011_10101000_11110011_0;
      patterns[19371] = 25'b01001011_10101001_11110100_0;
      patterns[19372] = 25'b01001011_10101010_11110101_0;
      patterns[19373] = 25'b01001011_10101011_11110110_0;
      patterns[19374] = 25'b01001011_10101100_11110111_0;
      patterns[19375] = 25'b01001011_10101101_11111000_0;
      patterns[19376] = 25'b01001011_10101110_11111001_0;
      patterns[19377] = 25'b01001011_10101111_11111010_0;
      patterns[19378] = 25'b01001011_10110000_11111011_0;
      patterns[19379] = 25'b01001011_10110001_11111100_0;
      patterns[19380] = 25'b01001011_10110010_11111101_0;
      patterns[19381] = 25'b01001011_10110011_11111110_0;
      patterns[19382] = 25'b01001011_10110100_11111111_0;
      patterns[19383] = 25'b01001011_10110101_00000000_1;
      patterns[19384] = 25'b01001011_10110110_00000001_1;
      patterns[19385] = 25'b01001011_10110111_00000010_1;
      patterns[19386] = 25'b01001011_10111000_00000011_1;
      patterns[19387] = 25'b01001011_10111001_00000100_1;
      patterns[19388] = 25'b01001011_10111010_00000101_1;
      patterns[19389] = 25'b01001011_10111011_00000110_1;
      patterns[19390] = 25'b01001011_10111100_00000111_1;
      patterns[19391] = 25'b01001011_10111101_00001000_1;
      patterns[19392] = 25'b01001011_10111110_00001001_1;
      patterns[19393] = 25'b01001011_10111111_00001010_1;
      patterns[19394] = 25'b01001011_11000000_00001011_1;
      patterns[19395] = 25'b01001011_11000001_00001100_1;
      patterns[19396] = 25'b01001011_11000010_00001101_1;
      patterns[19397] = 25'b01001011_11000011_00001110_1;
      patterns[19398] = 25'b01001011_11000100_00001111_1;
      patterns[19399] = 25'b01001011_11000101_00010000_1;
      patterns[19400] = 25'b01001011_11000110_00010001_1;
      patterns[19401] = 25'b01001011_11000111_00010010_1;
      patterns[19402] = 25'b01001011_11001000_00010011_1;
      patterns[19403] = 25'b01001011_11001001_00010100_1;
      patterns[19404] = 25'b01001011_11001010_00010101_1;
      patterns[19405] = 25'b01001011_11001011_00010110_1;
      patterns[19406] = 25'b01001011_11001100_00010111_1;
      patterns[19407] = 25'b01001011_11001101_00011000_1;
      patterns[19408] = 25'b01001011_11001110_00011001_1;
      patterns[19409] = 25'b01001011_11001111_00011010_1;
      patterns[19410] = 25'b01001011_11010000_00011011_1;
      patterns[19411] = 25'b01001011_11010001_00011100_1;
      patterns[19412] = 25'b01001011_11010010_00011101_1;
      patterns[19413] = 25'b01001011_11010011_00011110_1;
      patterns[19414] = 25'b01001011_11010100_00011111_1;
      patterns[19415] = 25'b01001011_11010101_00100000_1;
      patterns[19416] = 25'b01001011_11010110_00100001_1;
      patterns[19417] = 25'b01001011_11010111_00100010_1;
      patterns[19418] = 25'b01001011_11011000_00100011_1;
      patterns[19419] = 25'b01001011_11011001_00100100_1;
      patterns[19420] = 25'b01001011_11011010_00100101_1;
      patterns[19421] = 25'b01001011_11011011_00100110_1;
      patterns[19422] = 25'b01001011_11011100_00100111_1;
      patterns[19423] = 25'b01001011_11011101_00101000_1;
      patterns[19424] = 25'b01001011_11011110_00101001_1;
      patterns[19425] = 25'b01001011_11011111_00101010_1;
      patterns[19426] = 25'b01001011_11100000_00101011_1;
      patterns[19427] = 25'b01001011_11100001_00101100_1;
      patterns[19428] = 25'b01001011_11100010_00101101_1;
      patterns[19429] = 25'b01001011_11100011_00101110_1;
      patterns[19430] = 25'b01001011_11100100_00101111_1;
      patterns[19431] = 25'b01001011_11100101_00110000_1;
      patterns[19432] = 25'b01001011_11100110_00110001_1;
      patterns[19433] = 25'b01001011_11100111_00110010_1;
      patterns[19434] = 25'b01001011_11101000_00110011_1;
      patterns[19435] = 25'b01001011_11101001_00110100_1;
      patterns[19436] = 25'b01001011_11101010_00110101_1;
      patterns[19437] = 25'b01001011_11101011_00110110_1;
      patterns[19438] = 25'b01001011_11101100_00110111_1;
      patterns[19439] = 25'b01001011_11101101_00111000_1;
      patterns[19440] = 25'b01001011_11101110_00111001_1;
      patterns[19441] = 25'b01001011_11101111_00111010_1;
      patterns[19442] = 25'b01001011_11110000_00111011_1;
      patterns[19443] = 25'b01001011_11110001_00111100_1;
      patterns[19444] = 25'b01001011_11110010_00111101_1;
      patterns[19445] = 25'b01001011_11110011_00111110_1;
      patterns[19446] = 25'b01001011_11110100_00111111_1;
      patterns[19447] = 25'b01001011_11110101_01000000_1;
      patterns[19448] = 25'b01001011_11110110_01000001_1;
      patterns[19449] = 25'b01001011_11110111_01000010_1;
      patterns[19450] = 25'b01001011_11111000_01000011_1;
      patterns[19451] = 25'b01001011_11111001_01000100_1;
      patterns[19452] = 25'b01001011_11111010_01000101_1;
      patterns[19453] = 25'b01001011_11111011_01000110_1;
      patterns[19454] = 25'b01001011_11111100_01000111_1;
      patterns[19455] = 25'b01001011_11111101_01001000_1;
      patterns[19456] = 25'b01001011_11111110_01001001_1;
      patterns[19457] = 25'b01001011_11111111_01001010_1;
      patterns[19458] = 25'b01001100_00000000_01001100_0;
      patterns[19459] = 25'b01001100_00000001_01001101_0;
      patterns[19460] = 25'b01001100_00000010_01001110_0;
      patterns[19461] = 25'b01001100_00000011_01001111_0;
      patterns[19462] = 25'b01001100_00000100_01010000_0;
      patterns[19463] = 25'b01001100_00000101_01010001_0;
      patterns[19464] = 25'b01001100_00000110_01010010_0;
      patterns[19465] = 25'b01001100_00000111_01010011_0;
      patterns[19466] = 25'b01001100_00001000_01010100_0;
      patterns[19467] = 25'b01001100_00001001_01010101_0;
      patterns[19468] = 25'b01001100_00001010_01010110_0;
      patterns[19469] = 25'b01001100_00001011_01010111_0;
      patterns[19470] = 25'b01001100_00001100_01011000_0;
      patterns[19471] = 25'b01001100_00001101_01011001_0;
      patterns[19472] = 25'b01001100_00001110_01011010_0;
      patterns[19473] = 25'b01001100_00001111_01011011_0;
      patterns[19474] = 25'b01001100_00010000_01011100_0;
      patterns[19475] = 25'b01001100_00010001_01011101_0;
      patterns[19476] = 25'b01001100_00010010_01011110_0;
      patterns[19477] = 25'b01001100_00010011_01011111_0;
      patterns[19478] = 25'b01001100_00010100_01100000_0;
      patterns[19479] = 25'b01001100_00010101_01100001_0;
      patterns[19480] = 25'b01001100_00010110_01100010_0;
      patterns[19481] = 25'b01001100_00010111_01100011_0;
      patterns[19482] = 25'b01001100_00011000_01100100_0;
      patterns[19483] = 25'b01001100_00011001_01100101_0;
      patterns[19484] = 25'b01001100_00011010_01100110_0;
      patterns[19485] = 25'b01001100_00011011_01100111_0;
      patterns[19486] = 25'b01001100_00011100_01101000_0;
      patterns[19487] = 25'b01001100_00011101_01101001_0;
      patterns[19488] = 25'b01001100_00011110_01101010_0;
      patterns[19489] = 25'b01001100_00011111_01101011_0;
      patterns[19490] = 25'b01001100_00100000_01101100_0;
      patterns[19491] = 25'b01001100_00100001_01101101_0;
      patterns[19492] = 25'b01001100_00100010_01101110_0;
      patterns[19493] = 25'b01001100_00100011_01101111_0;
      patterns[19494] = 25'b01001100_00100100_01110000_0;
      patterns[19495] = 25'b01001100_00100101_01110001_0;
      patterns[19496] = 25'b01001100_00100110_01110010_0;
      patterns[19497] = 25'b01001100_00100111_01110011_0;
      patterns[19498] = 25'b01001100_00101000_01110100_0;
      patterns[19499] = 25'b01001100_00101001_01110101_0;
      patterns[19500] = 25'b01001100_00101010_01110110_0;
      patterns[19501] = 25'b01001100_00101011_01110111_0;
      patterns[19502] = 25'b01001100_00101100_01111000_0;
      patterns[19503] = 25'b01001100_00101101_01111001_0;
      patterns[19504] = 25'b01001100_00101110_01111010_0;
      patterns[19505] = 25'b01001100_00101111_01111011_0;
      patterns[19506] = 25'b01001100_00110000_01111100_0;
      patterns[19507] = 25'b01001100_00110001_01111101_0;
      patterns[19508] = 25'b01001100_00110010_01111110_0;
      patterns[19509] = 25'b01001100_00110011_01111111_0;
      patterns[19510] = 25'b01001100_00110100_10000000_0;
      patterns[19511] = 25'b01001100_00110101_10000001_0;
      patterns[19512] = 25'b01001100_00110110_10000010_0;
      patterns[19513] = 25'b01001100_00110111_10000011_0;
      patterns[19514] = 25'b01001100_00111000_10000100_0;
      patterns[19515] = 25'b01001100_00111001_10000101_0;
      patterns[19516] = 25'b01001100_00111010_10000110_0;
      patterns[19517] = 25'b01001100_00111011_10000111_0;
      patterns[19518] = 25'b01001100_00111100_10001000_0;
      patterns[19519] = 25'b01001100_00111101_10001001_0;
      patterns[19520] = 25'b01001100_00111110_10001010_0;
      patterns[19521] = 25'b01001100_00111111_10001011_0;
      patterns[19522] = 25'b01001100_01000000_10001100_0;
      patterns[19523] = 25'b01001100_01000001_10001101_0;
      patterns[19524] = 25'b01001100_01000010_10001110_0;
      patterns[19525] = 25'b01001100_01000011_10001111_0;
      patterns[19526] = 25'b01001100_01000100_10010000_0;
      patterns[19527] = 25'b01001100_01000101_10010001_0;
      patterns[19528] = 25'b01001100_01000110_10010010_0;
      patterns[19529] = 25'b01001100_01000111_10010011_0;
      patterns[19530] = 25'b01001100_01001000_10010100_0;
      patterns[19531] = 25'b01001100_01001001_10010101_0;
      patterns[19532] = 25'b01001100_01001010_10010110_0;
      patterns[19533] = 25'b01001100_01001011_10010111_0;
      patterns[19534] = 25'b01001100_01001100_10011000_0;
      patterns[19535] = 25'b01001100_01001101_10011001_0;
      patterns[19536] = 25'b01001100_01001110_10011010_0;
      patterns[19537] = 25'b01001100_01001111_10011011_0;
      patterns[19538] = 25'b01001100_01010000_10011100_0;
      patterns[19539] = 25'b01001100_01010001_10011101_0;
      patterns[19540] = 25'b01001100_01010010_10011110_0;
      patterns[19541] = 25'b01001100_01010011_10011111_0;
      patterns[19542] = 25'b01001100_01010100_10100000_0;
      patterns[19543] = 25'b01001100_01010101_10100001_0;
      patterns[19544] = 25'b01001100_01010110_10100010_0;
      patterns[19545] = 25'b01001100_01010111_10100011_0;
      patterns[19546] = 25'b01001100_01011000_10100100_0;
      patterns[19547] = 25'b01001100_01011001_10100101_0;
      patterns[19548] = 25'b01001100_01011010_10100110_0;
      patterns[19549] = 25'b01001100_01011011_10100111_0;
      patterns[19550] = 25'b01001100_01011100_10101000_0;
      patterns[19551] = 25'b01001100_01011101_10101001_0;
      patterns[19552] = 25'b01001100_01011110_10101010_0;
      patterns[19553] = 25'b01001100_01011111_10101011_0;
      patterns[19554] = 25'b01001100_01100000_10101100_0;
      patterns[19555] = 25'b01001100_01100001_10101101_0;
      patterns[19556] = 25'b01001100_01100010_10101110_0;
      patterns[19557] = 25'b01001100_01100011_10101111_0;
      patterns[19558] = 25'b01001100_01100100_10110000_0;
      patterns[19559] = 25'b01001100_01100101_10110001_0;
      patterns[19560] = 25'b01001100_01100110_10110010_0;
      patterns[19561] = 25'b01001100_01100111_10110011_0;
      patterns[19562] = 25'b01001100_01101000_10110100_0;
      patterns[19563] = 25'b01001100_01101001_10110101_0;
      patterns[19564] = 25'b01001100_01101010_10110110_0;
      patterns[19565] = 25'b01001100_01101011_10110111_0;
      patterns[19566] = 25'b01001100_01101100_10111000_0;
      patterns[19567] = 25'b01001100_01101101_10111001_0;
      patterns[19568] = 25'b01001100_01101110_10111010_0;
      patterns[19569] = 25'b01001100_01101111_10111011_0;
      patterns[19570] = 25'b01001100_01110000_10111100_0;
      patterns[19571] = 25'b01001100_01110001_10111101_0;
      patterns[19572] = 25'b01001100_01110010_10111110_0;
      patterns[19573] = 25'b01001100_01110011_10111111_0;
      patterns[19574] = 25'b01001100_01110100_11000000_0;
      patterns[19575] = 25'b01001100_01110101_11000001_0;
      patterns[19576] = 25'b01001100_01110110_11000010_0;
      patterns[19577] = 25'b01001100_01110111_11000011_0;
      patterns[19578] = 25'b01001100_01111000_11000100_0;
      patterns[19579] = 25'b01001100_01111001_11000101_0;
      patterns[19580] = 25'b01001100_01111010_11000110_0;
      patterns[19581] = 25'b01001100_01111011_11000111_0;
      patterns[19582] = 25'b01001100_01111100_11001000_0;
      patterns[19583] = 25'b01001100_01111101_11001001_0;
      patterns[19584] = 25'b01001100_01111110_11001010_0;
      patterns[19585] = 25'b01001100_01111111_11001011_0;
      patterns[19586] = 25'b01001100_10000000_11001100_0;
      patterns[19587] = 25'b01001100_10000001_11001101_0;
      patterns[19588] = 25'b01001100_10000010_11001110_0;
      patterns[19589] = 25'b01001100_10000011_11001111_0;
      patterns[19590] = 25'b01001100_10000100_11010000_0;
      patterns[19591] = 25'b01001100_10000101_11010001_0;
      patterns[19592] = 25'b01001100_10000110_11010010_0;
      patterns[19593] = 25'b01001100_10000111_11010011_0;
      patterns[19594] = 25'b01001100_10001000_11010100_0;
      patterns[19595] = 25'b01001100_10001001_11010101_0;
      patterns[19596] = 25'b01001100_10001010_11010110_0;
      patterns[19597] = 25'b01001100_10001011_11010111_0;
      patterns[19598] = 25'b01001100_10001100_11011000_0;
      patterns[19599] = 25'b01001100_10001101_11011001_0;
      patterns[19600] = 25'b01001100_10001110_11011010_0;
      patterns[19601] = 25'b01001100_10001111_11011011_0;
      patterns[19602] = 25'b01001100_10010000_11011100_0;
      patterns[19603] = 25'b01001100_10010001_11011101_0;
      patterns[19604] = 25'b01001100_10010010_11011110_0;
      patterns[19605] = 25'b01001100_10010011_11011111_0;
      patterns[19606] = 25'b01001100_10010100_11100000_0;
      patterns[19607] = 25'b01001100_10010101_11100001_0;
      patterns[19608] = 25'b01001100_10010110_11100010_0;
      patterns[19609] = 25'b01001100_10010111_11100011_0;
      patterns[19610] = 25'b01001100_10011000_11100100_0;
      patterns[19611] = 25'b01001100_10011001_11100101_0;
      patterns[19612] = 25'b01001100_10011010_11100110_0;
      patterns[19613] = 25'b01001100_10011011_11100111_0;
      patterns[19614] = 25'b01001100_10011100_11101000_0;
      patterns[19615] = 25'b01001100_10011101_11101001_0;
      patterns[19616] = 25'b01001100_10011110_11101010_0;
      patterns[19617] = 25'b01001100_10011111_11101011_0;
      patterns[19618] = 25'b01001100_10100000_11101100_0;
      patterns[19619] = 25'b01001100_10100001_11101101_0;
      patterns[19620] = 25'b01001100_10100010_11101110_0;
      patterns[19621] = 25'b01001100_10100011_11101111_0;
      patterns[19622] = 25'b01001100_10100100_11110000_0;
      patterns[19623] = 25'b01001100_10100101_11110001_0;
      patterns[19624] = 25'b01001100_10100110_11110010_0;
      patterns[19625] = 25'b01001100_10100111_11110011_0;
      patterns[19626] = 25'b01001100_10101000_11110100_0;
      patterns[19627] = 25'b01001100_10101001_11110101_0;
      patterns[19628] = 25'b01001100_10101010_11110110_0;
      patterns[19629] = 25'b01001100_10101011_11110111_0;
      patterns[19630] = 25'b01001100_10101100_11111000_0;
      patterns[19631] = 25'b01001100_10101101_11111001_0;
      patterns[19632] = 25'b01001100_10101110_11111010_0;
      patterns[19633] = 25'b01001100_10101111_11111011_0;
      patterns[19634] = 25'b01001100_10110000_11111100_0;
      patterns[19635] = 25'b01001100_10110001_11111101_0;
      patterns[19636] = 25'b01001100_10110010_11111110_0;
      patterns[19637] = 25'b01001100_10110011_11111111_0;
      patterns[19638] = 25'b01001100_10110100_00000000_1;
      patterns[19639] = 25'b01001100_10110101_00000001_1;
      patterns[19640] = 25'b01001100_10110110_00000010_1;
      patterns[19641] = 25'b01001100_10110111_00000011_1;
      patterns[19642] = 25'b01001100_10111000_00000100_1;
      patterns[19643] = 25'b01001100_10111001_00000101_1;
      patterns[19644] = 25'b01001100_10111010_00000110_1;
      patterns[19645] = 25'b01001100_10111011_00000111_1;
      patterns[19646] = 25'b01001100_10111100_00001000_1;
      patterns[19647] = 25'b01001100_10111101_00001001_1;
      patterns[19648] = 25'b01001100_10111110_00001010_1;
      patterns[19649] = 25'b01001100_10111111_00001011_1;
      patterns[19650] = 25'b01001100_11000000_00001100_1;
      patterns[19651] = 25'b01001100_11000001_00001101_1;
      patterns[19652] = 25'b01001100_11000010_00001110_1;
      patterns[19653] = 25'b01001100_11000011_00001111_1;
      patterns[19654] = 25'b01001100_11000100_00010000_1;
      patterns[19655] = 25'b01001100_11000101_00010001_1;
      patterns[19656] = 25'b01001100_11000110_00010010_1;
      patterns[19657] = 25'b01001100_11000111_00010011_1;
      patterns[19658] = 25'b01001100_11001000_00010100_1;
      patterns[19659] = 25'b01001100_11001001_00010101_1;
      patterns[19660] = 25'b01001100_11001010_00010110_1;
      patterns[19661] = 25'b01001100_11001011_00010111_1;
      patterns[19662] = 25'b01001100_11001100_00011000_1;
      patterns[19663] = 25'b01001100_11001101_00011001_1;
      patterns[19664] = 25'b01001100_11001110_00011010_1;
      patterns[19665] = 25'b01001100_11001111_00011011_1;
      patterns[19666] = 25'b01001100_11010000_00011100_1;
      patterns[19667] = 25'b01001100_11010001_00011101_1;
      patterns[19668] = 25'b01001100_11010010_00011110_1;
      patterns[19669] = 25'b01001100_11010011_00011111_1;
      patterns[19670] = 25'b01001100_11010100_00100000_1;
      patterns[19671] = 25'b01001100_11010101_00100001_1;
      patterns[19672] = 25'b01001100_11010110_00100010_1;
      patterns[19673] = 25'b01001100_11010111_00100011_1;
      patterns[19674] = 25'b01001100_11011000_00100100_1;
      patterns[19675] = 25'b01001100_11011001_00100101_1;
      patterns[19676] = 25'b01001100_11011010_00100110_1;
      patterns[19677] = 25'b01001100_11011011_00100111_1;
      patterns[19678] = 25'b01001100_11011100_00101000_1;
      patterns[19679] = 25'b01001100_11011101_00101001_1;
      patterns[19680] = 25'b01001100_11011110_00101010_1;
      patterns[19681] = 25'b01001100_11011111_00101011_1;
      patterns[19682] = 25'b01001100_11100000_00101100_1;
      patterns[19683] = 25'b01001100_11100001_00101101_1;
      patterns[19684] = 25'b01001100_11100010_00101110_1;
      patterns[19685] = 25'b01001100_11100011_00101111_1;
      patterns[19686] = 25'b01001100_11100100_00110000_1;
      patterns[19687] = 25'b01001100_11100101_00110001_1;
      patterns[19688] = 25'b01001100_11100110_00110010_1;
      patterns[19689] = 25'b01001100_11100111_00110011_1;
      patterns[19690] = 25'b01001100_11101000_00110100_1;
      patterns[19691] = 25'b01001100_11101001_00110101_1;
      patterns[19692] = 25'b01001100_11101010_00110110_1;
      patterns[19693] = 25'b01001100_11101011_00110111_1;
      patterns[19694] = 25'b01001100_11101100_00111000_1;
      patterns[19695] = 25'b01001100_11101101_00111001_1;
      patterns[19696] = 25'b01001100_11101110_00111010_1;
      patterns[19697] = 25'b01001100_11101111_00111011_1;
      patterns[19698] = 25'b01001100_11110000_00111100_1;
      patterns[19699] = 25'b01001100_11110001_00111101_1;
      patterns[19700] = 25'b01001100_11110010_00111110_1;
      patterns[19701] = 25'b01001100_11110011_00111111_1;
      patterns[19702] = 25'b01001100_11110100_01000000_1;
      patterns[19703] = 25'b01001100_11110101_01000001_1;
      patterns[19704] = 25'b01001100_11110110_01000010_1;
      patterns[19705] = 25'b01001100_11110111_01000011_1;
      patterns[19706] = 25'b01001100_11111000_01000100_1;
      patterns[19707] = 25'b01001100_11111001_01000101_1;
      patterns[19708] = 25'b01001100_11111010_01000110_1;
      patterns[19709] = 25'b01001100_11111011_01000111_1;
      patterns[19710] = 25'b01001100_11111100_01001000_1;
      patterns[19711] = 25'b01001100_11111101_01001001_1;
      patterns[19712] = 25'b01001100_11111110_01001010_1;
      patterns[19713] = 25'b01001100_11111111_01001011_1;
      patterns[19714] = 25'b01001101_00000000_01001101_0;
      patterns[19715] = 25'b01001101_00000001_01001110_0;
      patterns[19716] = 25'b01001101_00000010_01001111_0;
      patterns[19717] = 25'b01001101_00000011_01010000_0;
      patterns[19718] = 25'b01001101_00000100_01010001_0;
      patterns[19719] = 25'b01001101_00000101_01010010_0;
      patterns[19720] = 25'b01001101_00000110_01010011_0;
      patterns[19721] = 25'b01001101_00000111_01010100_0;
      patterns[19722] = 25'b01001101_00001000_01010101_0;
      patterns[19723] = 25'b01001101_00001001_01010110_0;
      patterns[19724] = 25'b01001101_00001010_01010111_0;
      patterns[19725] = 25'b01001101_00001011_01011000_0;
      patterns[19726] = 25'b01001101_00001100_01011001_0;
      patterns[19727] = 25'b01001101_00001101_01011010_0;
      patterns[19728] = 25'b01001101_00001110_01011011_0;
      patterns[19729] = 25'b01001101_00001111_01011100_0;
      patterns[19730] = 25'b01001101_00010000_01011101_0;
      patterns[19731] = 25'b01001101_00010001_01011110_0;
      patterns[19732] = 25'b01001101_00010010_01011111_0;
      patterns[19733] = 25'b01001101_00010011_01100000_0;
      patterns[19734] = 25'b01001101_00010100_01100001_0;
      patterns[19735] = 25'b01001101_00010101_01100010_0;
      patterns[19736] = 25'b01001101_00010110_01100011_0;
      patterns[19737] = 25'b01001101_00010111_01100100_0;
      patterns[19738] = 25'b01001101_00011000_01100101_0;
      patterns[19739] = 25'b01001101_00011001_01100110_0;
      patterns[19740] = 25'b01001101_00011010_01100111_0;
      patterns[19741] = 25'b01001101_00011011_01101000_0;
      patterns[19742] = 25'b01001101_00011100_01101001_0;
      patterns[19743] = 25'b01001101_00011101_01101010_0;
      patterns[19744] = 25'b01001101_00011110_01101011_0;
      patterns[19745] = 25'b01001101_00011111_01101100_0;
      patterns[19746] = 25'b01001101_00100000_01101101_0;
      patterns[19747] = 25'b01001101_00100001_01101110_0;
      patterns[19748] = 25'b01001101_00100010_01101111_0;
      patterns[19749] = 25'b01001101_00100011_01110000_0;
      patterns[19750] = 25'b01001101_00100100_01110001_0;
      patterns[19751] = 25'b01001101_00100101_01110010_0;
      patterns[19752] = 25'b01001101_00100110_01110011_0;
      patterns[19753] = 25'b01001101_00100111_01110100_0;
      patterns[19754] = 25'b01001101_00101000_01110101_0;
      patterns[19755] = 25'b01001101_00101001_01110110_0;
      patterns[19756] = 25'b01001101_00101010_01110111_0;
      patterns[19757] = 25'b01001101_00101011_01111000_0;
      patterns[19758] = 25'b01001101_00101100_01111001_0;
      patterns[19759] = 25'b01001101_00101101_01111010_0;
      patterns[19760] = 25'b01001101_00101110_01111011_0;
      patterns[19761] = 25'b01001101_00101111_01111100_0;
      patterns[19762] = 25'b01001101_00110000_01111101_0;
      patterns[19763] = 25'b01001101_00110001_01111110_0;
      patterns[19764] = 25'b01001101_00110010_01111111_0;
      patterns[19765] = 25'b01001101_00110011_10000000_0;
      patterns[19766] = 25'b01001101_00110100_10000001_0;
      patterns[19767] = 25'b01001101_00110101_10000010_0;
      patterns[19768] = 25'b01001101_00110110_10000011_0;
      patterns[19769] = 25'b01001101_00110111_10000100_0;
      patterns[19770] = 25'b01001101_00111000_10000101_0;
      patterns[19771] = 25'b01001101_00111001_10000110_0;
      patterns[19772] = 25'b01001101_00111010_10000111_0;
      patterns[19773] = 25'b01001101_00111011_10001000_0;
      patterns[19774] = 25'b01001101_00111100_10001001_0;
      patterns[19775] = 25'b01001101_00111101_10001010_0;
      patterns[19776] = 25'b01001101_00111110_10001011_0;
      patterns[19777] = 25'b01001101_00111111_10001100_0;
      patterns[19778] = 25'b01001101_01000000_10001101_0;
      patterns[19779] = 25'b01001101_01000001_10001110_0;
      patterns[19780] = 25'b01001101_01000010_10001111_0;
      patterns[19781] = 25'b01001101_01000011_10010000_0;
      patterns[19782] = 25'b01001101_01000100_10010001_0;
      patterns[19783] = 25'b01001101_01000101_10010010_0;
      patterns[19784] = 25'b01001101_01000110_10010011_0;
      patterns[19785] = 25'b01001101_01000111_10010100_0;
      patterns[19786] = 25'b01001101_01001000_10010101_0;
      patterns[19787] = 25'b01001101_01001001_10010110_0;
      patterns[19788] = 25'b01001101_01001010_10010111_0;
      patterns[19789] = 25'b01001101_01001011_10011000_0;
      patterns[19790] = 25'b01001101_01001100_10011001_0;
      patterns[19791] = 25'b01001101_01001101_10011010_0;
      patterns[19792] = 25'b01001101_01001110_10011011_0;
      patterns[19793] = 25'b01001101_01001111_10011100_0;
      patterns[19794] = 25'b01001101_01010000_10011101_0;
      patterns[19795] = 25'b01001101_01010001_10011110_0;
      patterns[19796] = 25'b01001101_01010010_10011111_0;
      patterns[19797] = 25'b01001101_01010011_10100000_0;
      patterns[19798] = 25'b01001101_01010100_10100001_0;
      patterns[19799] = 25'b01001101_01010101_10100010_0;
      patterns[19800] = 25'b01001101_01010110_10100011_0;
      patterns[19801] = 25'b01001101_01010111_10100100_0;
      patterns[19802] = 25'b01001101_01011000_10100101_0;
      patterns[19803] = 25'b01001101_01011001_10100110_0;
      patterns[19804] = 25'b01001101_01011010_10100111_0;
      patterns[19805] = 25'b01001101_01011011_10101000_0;
      patterns[19806] = 25'b01001101_01011100_10101001_0;
      patterns[19807] = 25'b01001101_01011101_10101010_0;
      patterns[19808] = 25'b01001101_01011110_10101011_0;
      patterns[19809] = 25'b01001101_01011111_10101100_0;
      patterns[19810] = 25'b01001101_01100000_10101101_0;
      patterns[19811] = 25'b01001101_01100001_10101110_0;
      patterns[19812] = 25'b01001101_01100010_10101111_0;
      patterns[19813] = 25'b01001101_01100011_10110000_0;
      patterns[19814] = 25'b01001101_01100100_10110001_0;
      patterns[19815] = 25'b01001101_01100101_10110010_0;
      patterns[19816] = 25'b01001101_01100110_10110011_0;
      patterns[19817] = 25'b01001101_01100111_10110100_0;
      patterns[19818] = 25'b01001101_01101000_10110101_0;
      patterns[19819] = 25'b01001101_01101001_10110110_0;
      patterns[19820] = 25'b01001101_01101010_10110111_0;
      patterns[19821] = 25'b01001101_01101011_10111000_0;
      patterns[19822] = 25'b01001101_01101100_10111001_0;
      patterns[19823] = 25'b01001101_01101101_10111010_0;
      patterns[19824] = 25'b01001101_01101110_10111011_0;
      patterns[19825] = 25'b01001101_01101111_10111100_0;
      patterns[19826] = 25'b01001101_01110000_10111101_0;
      patterns[19827] = 25'b01001101_01110001_10111110_0;
      patterns[19828] = 25'b01001101_01110010_10111111_0;
      patterns[19829] = 25'b01001101_01110011_11000000_0;
      patterns[19830] = 25'b01001101_01110100_11000001_0;
      patterns[19831] = 25'b01001101_01110101_11000010_0;
      patterns[19832] = 25'b01001101_01110110_11000011_0;
      patterns[19833] = 25'b01001101_01110111_11000100_0;
      patterns[19834] = 25'b01001101_01111000_11000101_0;
      patterns[19835] = 25'b01001101_01111001_11000110_0;
      patterns[19836] = 25'b01001101_01111010_11000111_0;
      patterns[19837] = 25'b01001101_01111011_11001000_0;
      patterns[19838] = 25'b01001101_01111100_11001001_0;
      patterns[19839] = 25'b01001101_01111101_11001010_0;
      patterns[19840] = 25'b01001101_01111110_11001011_0;
      patterns[19841] = 25'b01001101_01111111_11001100_0;
      patterns[19842] = 25'b01001101_10000000_11001101_0;
      patterns[19843] = 25'b01001101_10000001_11001110_0;
      patterns[19844] = 25'b01001101_10000010_11001111_0;
      patterns[19845] = 25'b01001101_10000011_11010000_0;
      patterns[19846] = 25'b01001101_10000100_11010001_0;
      patterns[19847] = 25'b01001101_10000101_11010010_0;
      patterns[19848] = 25'b01001101_10000110_11010011_0;
      patterns[19849] = 25'b01001101_10000111_11010100_0;
      patterns[19850] = 25'b01001101_10001000_11010101_0;
      patterns[19851] = 25'b01001101_10001001_11010110_0;
      patterns[19852] = 25'b01001101_10001010_11010111_0;
      patterns[19853] = 25'b01001101_10001011_11011000_0;
      patterns[19854] = 25'b01001101_10001100_11011001_0;
      patterns[19855] = 25'b01001101_10001101_11011010_0;
      patterns[19856] = 25'b01001101_10001110_11011011_0;
      patterns[19857] = 25'b01001101_10001111_11011100_0;
      patterns[19858] = 25'b01001101_10010000_11011101_0;
      patterns[19859] = 25'b01001101_10010001_11011110_0;
      patterns[19860] = 25'b01001101_10010010_11011111_0;
      patterns[19861] = 25'b01001101_10010011_11100000_0;
      patterns[19862] = 25'b01001101_10010100_11100001_0;
      patterns[19863] = 25'b01001101_10010101_11100010_0;
      patterns[19864] = 25'b01001101_10010110_11100011_0;
      patterns[19865] = 25'b01001101_10010111_11100100_0;
      patterns[19866] = 25'b01001101_10011000_11100101_0;
      patterns[19867] = 25'b01001101_10011001_11100110_0;
      patterns[19868] = 25'b01001101_10011010_11100111_0;
      patterns[19869] = 25'b01001101_10011011_11101000_0;
      patterns[19870] = 25'b01001101_10011100_11101001_0;
      patterns[19871] = 25'b01001101_10011101_11101010_0;
      patterns[19872] = 25'b01001101_10011110_11101011_0;
      patterns[19873] = 25'b01001101_10011111_11101100_0;
      patterns[19874] = 25'b01001101_10100000_11101101_0;
      patterns[19875] = 25'b01001101_10100001_11101110_0;
      patterns[19876] = 25'b01001101_10100010_11101111_0;
      patterns[19877] = 25'b01001101_10100011_11110000_0;
      patterns[19878] = 25'b01001101_10100100_11110001_0;
      patterns[19879] = 25'b01001101_10100101_11110010_0;
      patterns[19880] = 25'b01001101_10100110_11110011_0;
      patterns[19881] = 25'b01001101_10100111_11110100_0;
      patterns[19882] = 25'b01001101_10101000_11110101_0;
      patterns[19883] = 25'b01001101_10101001_11110110_0;
      patterns[19884] = 25'b01001101_10101010_11110111_0;
      patterns[19885] = 25'b01001101_10101011_11111000_0;
      patterns[19886] = 25'b01001101_10101100_11111001_0;
      patterns[19887] = 25'b01001101_10101101_11111010_0;
      patterns[19888] = 25'b01001101_10101110_11111011_0;
      patterns[19889] = 25'b01001101_10101111_11111100_0;
      patterns[19890] = 25'b01001101_10110000_11111101_0;
      patterns[19891] = 25'b01001101_10110001_11111110_0;
      patterns[19892] = 25'b01001101_10110010_11111111_0;
      patterns[19893] = 25'b01001101_10110011_00000000_1;
      patterns[19894] = 25'b01001101_10110100_00000001_1;
      patterns[19895] = 25'b01001101_10110101_00000010_1;
      patterns[19896] = 25'b01001101_10110110_00000011_1;
      patterns[19897] = 25'b01001101_10110111_00000100_1;
      patterns[19898] = 25'b01001101_10111000_00000101_1;
      patterns[19899] = 25'b01001101_10111001_00000110_1;
      patterns[19900] = 25'b01001101_10111010_00000111_1;
      patterns[19901] = 25'b01001101_10111011_00001000_1;
      patterns[19902] = 25'b01001101_10111100_00001001_1;
      patterns[19903] = 25'b01001101_10111101_00001010_1;
      patterns[19904] = 25'b01001101_10111110_00001011_1;
      patterns[19905] = 25'b01001101_10111111_00001100_1;
      patterns[19906] = 25'b01001101_11000000_00001101_1;
      patterns[19907] = 25'b01001101_11000001_00001110_1;
      patterns[19908] = 25'b01001101_11000010_00001111_1;
      patterns[19909] = 25'b01001101_11000011_00010000_1;
      patterns[19910] = 25'b01001101_11000100_00010001_1;
      patterns[19911] = 25'b01001101_11000101_00010010_1;
      patterns[19912] = 25'b01001101_11000110_00010011_1;
      patterns[19913] = 25'b01001101_11000111_00010100_1;
      patterns[19914] = 25'b01001101_11001000_00010101_1;
      patterns[19915] = 25'b01001101_11001001_00010110_1;
      patterns[19916] = 25'b01001101_11001010_00010111_1;
      patterns[19917] = 25'b01001101_11001011_00011000_1;
      patterns[19918] = 25'b01001101_11001100_00011001_1;
      patterns[19919] = 25'b01001101_11001101_00011010_1;
      patterns[19920] = 25'b01001101_11001110_00011011_1;
      patterns[19921] = 25'b01001101_11001111_00011100_1;
      patterns[19922] = 25'b01001101_11010000_00011101_1;
      patterns[19923] = 25'b01001101_11010001_00011110_1;
      patterns[19924] = 25'b01001101_11010010_00011111_1;
      patterns[19925] = 25'b01001101_11010011_00100000_1;
      patterns[19926] = 25'b01001101_11010100_00100001_1;
      patterns[19927] = 25'b01001101_11010101_00100010_1;
      patterns[19928] = 25'b01001101_11010110_00100011_1;
      patterns[19929] = 25'b01001101_11010111_00100100_1;
      patterns[19930] = 25'b01001101_11011000_00100101_1;
      patterns[19931] = 25'b01001101_11011001_00100110_1;
      patterns[19932] = 25'b01001101_11011010_00100111_1;
      patterns[19933] = 25'b01001101_11011011_00101000_1;
      patterns[19934] = 25'b01001101_11011100_00101001_1;
      patterns[19935] = 25'b01001101_11011101_00101010_1;
      patterns[19936] = 25'b01001101_11011110_00101011_1;
      patterns[19937] = 25'b01001101_11011111_00101100_1;
      patterns[19938] = 25'b01001101_11100000_00101101_1;
      patterns[19939] = 25'b01001101_11100001_00101110_1;
      patterns[19940] = 25'b01001101_11100010_00101111_1;
      patterns[19941] = 25'b01001101_11100011_00110000_1;
      patterns[19942] = 25'b01001101_11100100_00110001_1;
      patterns[19943] = 25'b01001101_11100101_00110010_1;
      patterns[19944] = 25'b01001101_11100110_00110011_1;
      patterns[19945] = 25'b01001101_11100111_00110100_1;
      patterns[19946] = 25'b01001101_11101000_00110101_1;
      patterns[19947] = 25'b01001101_11101001_00110110_1;
      patterns[19948] = 25'b01001101_11101010_00110111_1;
      patterns[19949] = 25'b01001101_11101011_00111000_1;
      patterns[19950] = 25'b01001101_11101100_00111001_1;
      patterns[19951] = 25'b01001101_11101101_00111010_1;
      patterns[19952] = 25'b01001101_11101110_00111011_1;
      patterns[19953] = 25'b01001101_11101111_00111100_1;
      patterns[19954] = 25'b01001101_11110000_00111101_1;
      patterns[19955] = 25'b01001101_11110001_00111110_1;
      patterns[19956] = 25'b01001101_11110010_00111111_1;
      patterns[19957] = 25'b01001101_11110011_01000000_1;
      patterns[19958] = 25'b01001101_11110100_01000001_1;
      patterns[19959] = 25'b01001101_11110101_01000010_1;
      patterns[19960] = 25'b01001101_11110110_01000011_1;
      patterns[19961] = 25'b01001101_11110111_01000100_1;
      patterns[19962] = 25'b01001101_11111000_01000101_1;
      patterns[19963] = 25'b01001101_11111001_01000110_1;
      patterns[19964] = 25'b01001101_11111010_01000111_1;
      patterns[19965] = 25'b01001101_11111011_01001000_1;
      patterns[19966] = 25'b01001101_11111100_01001001_1;
      patterns[19967] = 25'b01001101_11111101_01001010_1;
      patterns[19968] = 25'b01001101_11111110_01001011_1;
      patterns[19969] = 25'b01001101_11111111_01001100_1;
      patterns[19970] = 25'b01001110_00000000_01001110_0;
      patterns[19971] = 25'b01001110_00000001_01001111_0;
      patterns[19972] = 25'b01001110_00000010_01010000_0;
      patterns[19973] = 25'b01001110_00000011_01010001_0;
      patterns[19974] = 25'b01001110_00000100_01010010_0;
      patterns[19975] = 25'b01001110_00000101_01010011_0;
      patterns[19976] = 25'b01001110_00000110_01010100_0;
      patterns[19977] = 25'b01001110_00000111_01010101_0;
      patterns[19978] = 25'b01001110_00001000_01010110_0;
      patterns[19979] = 25'b01001110_00001001_01010111_0;
      patterns[19980] = 25'b01001110_00001010_01011000_0;
      patterns[19981] = 25'b01001110_00001011_01011001_0;
      patterns[19982] = 25'b01001110_00001100_01011010_0;
      patterns[19983] = 25'b01001110_00001101_01011011_0;
      patterns[19984] = 25'b01001110_00001110_01011100_0;
      patterns[19985] = 25'b01001110_00001111_01011101_0;
      patterns[19986] = 25'b01001110_00010000_01011110_0;
      patterns[19987] = 25'b01001110_00010001_01011111_0;
      patterns[19988] = 25'b01001110_00010010_01100000_0;
      patterns[19989] = 25'b01001110_00010011_01100001_0;
      patterns[19990] = 25'b01001110_00010100_01100010_0;
      patterns[19991] = 25'b01001110_00010101_01100011_0;
      patterns[19992] = 25'b01001110_00010110_01100100_0;
      patterns[19993] = 25'b01001110_00010111_01100101_0;
      patterns[19994] = 25'b01001110_00011000_01100110_0;
      patterns[19995] = 25'b01001110_00011001_01100111_0;
      patterns[19996] = 25'b01001110_00011010_01101000_0;
      patterns[19997] = 25'b01001110_00011011_01101001_0;
      patterns[19998] = 25'b01001110_00011100_01101010_0;
      patterns[19999] = 25'b01001110_00011101_01101011_0;
      patterns[20000] = 25'b01001110_00011110_01101100_0;
      patterns[20001] = 25'b01001110_00011111_01101101_0;
      patterns[20002] = 25'b01001110_00100000_01101110_0;
      patterns[20003] = 25'b01001110_00100001_01101111_0;
      patterns[20004] = 25'b01001110_00100010_01110000_0;
      patterns[20005] = 25'b01001110_00100011_01110001_0;
      patterns[20006] = 25'b01001110_00100100_01110010_0;
      patterns[20007] = 25'b01001110_00100101_01110011_0;
      patterns[20008] = 25'b01001110_00100110_01110100_0;
      patterns[20009] = 25'b01001110_00100111_01110101_0;
      patterns[20010] = 25'b01001110_00101000_01110110_0;
      patterns[20011] = 25'b01001110_00101001_01110111_0;
      patterns[20012] = 25'b01001110_00101010_01111000_0;
      patterns[20013] = 25'b01001110_00101011_01111001_0;
      patterns[20014] = 25'b01001110_00101100_01111010_0;
      patterns[20015] = 25'b01001110_00101101_01111011_0;
      patterns[20016] = 25'b01001110_00101110_01111100_0;
      patterns[20017] = 25'b01001110_00101111_01111101_0;
      patterns[20018] = 25'b01001110_00110000_01111110_0;
      patterns[20019] = 25'b01001110_00110001_01111111_0;
      patterns[20020] = 25'b01001110_00110010_10000000_0;
      patterns[20021] = 25'b01001110_00110011_10000001_0;
      patterns[20022] = 25'b01001110_00110100_10000010_0;
      patterns[20023] = 25'b01001110_00110101_10000011_0;
      patterns[20024] = 25'b01001110_00110110_10000100_0;
      patterns[20025] = 25'b01001110_00110111_10000101_0;
      patterns[20026] = 25'b01001110_00111000_10000110_0;
      patterns[20027] = 25'b01001110_00111001_10000111_0;
      patterns[20028] = 25'b01001110_00111010_10001000_0;
      patterns[20029] = 25'b01001110_00111011_10001001_0;
      patterns[20030] = 25'b01001110_00111100_10001010_0;
      patterns[20031] = 25'b01001110_00111101_10001011_0;
      patterns[20032] = 25'b01001110_00111110_10001100_0;
      patterns[20033] = 25'b01001110_00111111_10001101_0;
      patterns[20034] = 25'b01001110_01000000_10001110_0;
      patterns[20035] = 25'b01001110_01000001_10001111_0;
      patterns[20036] = 25'b01001110_01000010_10010000_0;
      patterns[20037] = 25'b01001110_01000011_10010001_0;
      patterns[20038] = 25'b01001110_01000100_10010010_0;
      patterns[20039] = 25'b01001110_01000101_10010011_0;
      patterns[20040] = 25'b01001110_01000110_10010100_0;
      patterns[20041] = 25'b01001110_01000111_10010101_0;
      patterns[20042] = 25'b01001110_01001000_10010110_0;
      patterns[20043] = 25'b01001110_01001001_10010111_0;
      patterns[20044] = 25'b01001110_01001010_10011000_0;
      patterns[20045] = 25'b01001110_01001011_10011001_0;
      patterns[20046] = 25'b01001110_01001100_10011010_0;
      patterns[20047] = 25'b01001110_01001101_10011011_0;
      patterns[20048] = 25'b01001110_01001110_10011100_0;
      patterns[20049] = 25'b01001110_01001111_10011101_0;
      patterns[20050] = 25'b01001110_01010000_10011110_0;
      patterns[20051] = 25'b01001110_01010001_10011111_0;
      patterns[20052] = 25'b01001110_01010010_10100000_0;
      patterns[20053] = 25'b01001110_01010011_10100001_0;
      patterns[20054] = 25'b01001110_01010100_10100010_0;
      patterns[20055] = 25'b01001110_01010101_10100011_0;
      patterns[20056] = 25'b01001110_01010110_10100100_0;
      patterns[20057] = 25'b01001110_01010111_10100101_0;
      patterns[20058] = 25'b01001110_01011000_10100110_0;
      patterns[20059] = 25'b01001110_01011001_10100111_0;
      patterns[20060] = 25'b01001110_01011010_10101000_0;
      patterns[20061] = 25'b01001110_01011011_10101001_0;
      patterns[20062] = 25'b01001110_01011100_10101010_0;
      patterns[20063] = 25'b01001110_01011101_10101011_0;
      patterns[20064] = 25'b01001110_01011110_10101100_0;
      patterns[20065] = 25'b01001110_01011111_10101101_0;
      patterns[20066] = 25'b01001110_01100000_10101110_0;
      patterns[20067] = 25'b01001110_01100001_10101111_0;
      patterns[20068] = 25'b01001110_01100010_10110000_0;
      patterns[20069] = 25'b01001110_01100011_10110001_0;
      patterns[20070] = 25'b01001110_01100100_10110010_0;
      patterns[20071] = 25'b01001110_01100101_10110011_0;
      patterns[20072] = 25'b01001110_01100110_10110100_0;
      patterns[20073] = 25'b01001110_01100111_10110101_0;
      patterns[20074] = 25'b01001110_01101000_10110110_0;
      patterns[20075] = 25'b01001110_01101001_10110111_0;
      patterns[20076] = 25'b01001110_01101010_10111000_0;
      patterns[20077] = 25'b01001110_01101011_10111001_0;
      patterns[20078] = 25'b01001110_01101100_10111010_0;
      patterns[20079] = 25'b01001110_01101101_10111011_0;
      patterns[20080] = 25'b01001110_01101110_10111100_0;
      patterns[20081] = 25'b01001110_01101111_10111101_0;
      patterns[20082] = 25'b01001110_01110000_10111110_0;
      patterns[20083] = 25'b01001110_01110001_10111111_0;
      patterns[20084] = 25'b01001110_01110010_11000000_0;
      patterns[20085] = 25'b01001110_01110011_11000001_0;
      patterns[20086] = 25'b01001110_01110100_11000010_0;
      patterns[20087] = 25'b01001110_01110101_11000011_0;
      patterns[20088] = 25'b01001110_01110110_11000100_0;
      patterns[20089] = 25'b01001110_01110111_11000101_0;
      patterns[20090] = 25'b01001110_01111000_11000110_0;
      patterns[20091] = 25'b01001110_01111001_11000111_0;
      patterns[20092] = 25'b01001110_01111010_11001000_0;
      patterns[20093] = 25'b01001110_01111011_11001001_0;
      patterns[20094] = 25'b01001110_01111100_11001010_0;
      patterns[20095] = 25'b01001110_01111101_11001011_0;
      patterns[20096] = 25'b01001110_01111110_11001100_0;
      patterns[20097] = 25'b01001110_01111111_11001101_0;
      patterns[20098] = 25'b01001110_10000000_11001110_0;
      patterns[20099] = 25'b01001110_10000001_11001111_0;
      patterns[20100] = 25'b01001110_10000010_11010000_0;
      patterns[20101] = 25'b01001110_10000011_11010001_0;
      patterns[20102] = 25'b01001110_10000100_11010010_0;
      patterns[20103] = 25'b01001110_10000101_11010011_0;
      patterns[20104] = 25'b01001110_10000110_11010100_0;
      patterns[20105] = 25'b01001110_10000111_11010101_0;
      patterns[20106] = 25'b01001110_10001000_11010110_0;
      patterns[20107] = 25'b01001110_10001001_11010111_0;
      patterns[20108] = 25'b01001110_10001010_11011000_0;
      patterns[20109] = 25'b01001110_10001011_11011001_0;
      patterns[20110] = 25'b01001110_10001100_11011010_0;
      patterns[20111] = 25'b01001110_10001101_11011011_0;
      patterns[20112] = 25'b01001110_10001110_11011100_0;
      patterns[20113] = 25'b01001110_10001111_11011101_0;
      patterns[20114] = 25'b01001110_10010000_11011110_0;
      patterns[20115] = 25'b01001110_10010001_11011111_0;
      patterns[20116] = 25'b01001110_10010010_11100000_0;
      patterns[20117] = 25'b01001110_10010011_11100001_0;
      patterns[20118] = 25'b01001110_10010100_11100010_0;
      patterns[20119] = 25'b01001110_10010101_11100011_0;
      patterns[20120] = 25'b01001110_10010110_11100100_0;
      patterns[20121] = 25'b01001110_10010111_11100101_0;
      patterns[20122] = 25'b01001110_10011000_11100110_0;
      patterns[20123] = 25'b01001110_10011001_11100111_0;
      patterns[20124] = 25'b01001110_10011010_11101000_0;
      patterns[20125] = 25'b01001110_10011011_11101001_0;
      patterns[20126] = 25'b01001110_10011100_11101010_0;
      patterns[20127] = 25'b01001110_10011101_11101011_0;
      patterns[20128] = 25'b01001110_10011110_11101100_0;
      patterns[20129] = 25'b01001110_10011111_11101101_0;
      patterns[20130] = 25'b01001110_10100000_11101110_0;
      patterns[20131] = 25'b01001110_10100001_11101111_0;
      patterns[20132] = 25'b01001110_10100010_11110000_0;
      patterns[20133] = 25'b01001110_10100011_11110001_0;
      patterns[20134] = 25'b01001110_10100100_11110010_0;
      patterns[20135] = 25'b01001110_10100101_11110011_0;
      patterns[20136] = 25'b01001110_10100110_11110100_0;
      patterns[20137] = 25'b01001110_10100111_11110101_0;
      patterns[20138] = 25'b01001110_10101000_11110110_0;
      patterns[20139] = 25'b01001110_10101001_11110111_0;
      patterns[20140] = 25'b01001110_10101010_11111000_0;
      patterns[20141] = 25'b01001110_10101011_11111001_0;
      patterns[20142] = 25'b01001110_10101100_11111010_0;
      patterns[20143] = 25'b01001110_10101101_11111011_0;
      patterns[20144] = 25'b01001110_10101110_11111100_0;
      patterns[20145] = 25'b01001110_10101111_11111101_0;
      patterns[20146] = 25'b01001110_10110000_11111110_0;
      patterns[20147] = 25'b01001110_10110001_11111111_0;
      patterns[20148] = 25'b01001110_10110010_00000000_1;
      patterns[20149] = 25'b01001110_10110011_00000001_1;
      patterns[20150] = 25'b01001110_10110100_00000010_1;
      patterns[20151] = 25'b01001110_10110101_00000011_1;
      patterns[20152] = 25'b01001110_10110110_00000100_1;
      patterns[20153] = 25'b01001110_10110111_00000101_1;
      patterns[20154] = 25'b01001110_10111000_00000110_1;
      patterns[20155] = 25'b01001110_10111001_00000111_1;
      patterns[20156] = 25'b01001110_10111010_00001000_1;
      patterns[20157] = 25'b01001110_10111011_00001001_1;
      patterns[20158] = 25'b01001110_10111100_00001010_1;
      patterns[20159] = 25'b01001110_10111101_00001011_1;
      patterns[20160] = 25'b01001110_10111110_00001100_1;
      patterns[20161] = 25'b01001110_10111111_00001101_1;
      patterns[20162] = 25'b01001110_11000000_00001110_1;
      patterns[20163] = 25'b01001110_11000001_00001111_1;
      patterns[20164] = 25'b01001110_11000010_00010000_1;
      patterns[20165] = 25'b01001110_11000011_00010001_1;
      patterns[20166] = 25'b01001110_11000100_00010010_1;
      patterns[20167] = 25'b01001110_11000101_00010011_1;
      patterns[20168] = 25'b01001110_11000110_00010100_1;
      patterns[20169] = 25'b01001110_11000111_00010101_1;
      patterns[20170] = 25'b01001110_11001000_00010110_1;
      patterns[20171] = 25'b01001110_11001001_00010111_1;
      patterns[20172] = 25'b01001110_11001010_00011000_1;
      patterns[20173] = 25'b01001110_11001011_00011001_1;
      patterns[20174] = 25'b01001110_11001100_00011010_1;
      patterns[20175] = 25'b01001110_11001101_00011011_1;
      patterns[20176] = 25'b01001110_11001110_00011100_1;
      patterns[20177] = 25'b01001110_11001111_00011101_1;
      patterns[20178] = 25'b01001110_11010000_00011110_1;
      patterns[20179] = 25'b01001110_11010001_00011111_1;
      patterns[20180] = 25'b01001110_11010010_00100000_1;
      patterns[20181] = 25'b01001110_11010011_00100001_1;
      patterns[20182] = 25'b01001110_11010100_00100010_1;
      patterns[20183] = 25'b01001110_11010101_00100011_1;
      patterns[20184] = 25'b01001110_11010110_00100100_1;
      patterns[20185] = 25'b01001110_11010111_00100101_1;
      patterns[20186] = 25'b01001110_11011000_00100110_1;
      patterns[20187] = 25'b01001110_11011001_00100111_1;
      patterns[20188] = 25'b01001110_11011010_00101000_1;
      patterns[20189] = 25'b01001110_11011011_00101001_1;
      patterns[20190] = 25'b01001110_11011100_00101010_1;
      patterns[20191] = 25'b01001110_11011101_00101011_1;
      patterns[20192] = 25'b01001110_11011110_00101100_1;
      patterns[20193] = 25'b01001110_11011111_00101101_1;
      patterns[20194] = 25'b01001110_11100000_00101110_1;
      patterns[20195] = 25'b01001110_11100001_00101111_1;
      patterns[20196] = 25'b01001110_11100010_00110000_1;
      patterns[20197] = 25'b01001110_11100011_00110001_1;
      patterns[20198] = 25'b01001110_11100100_00110010_1;
      patterns[20199] = 25'b01001110_11100101_00110011_1;
      patterns[20200] = 25'b01001110_11100110_00110100_1;
      patterns[20201] = 25'b01001110_11100111_00110101_1;
      patterns[20202] = 25'b01001110_11101000_00110110_1;
      patterns[20203] = 25'b01001110_11101001_00110111_1;
      patterns[20204] = 25'b01001110_11101010_00111000_1;
      patterns[20205] = 25'b01001110_11101011_00111001_1;
      patterns[20206] = 25'b01001110_11101100_00111010_1;
      patterns[20207] = 25'b01001110_11101101_00111011_1;
      patterns[20208] = 25'b01001110_11101110_00111100_1;
      patterns[20209] = 25'b01001110_11101111_00111101_1;
      patterns[20210] = 25'b01001110_11110000_00111110_1;
      patterns[20211] = 25'b01001110_11110001_00111111_1;
      patterns[20212] = 25'b01001110_11110010_01000000_1;
      patterns[20213] = 25'b01001110_11110011_01000001_1;
      patterns[20214] = 25'b01001110_11110100_01000010_1;
      patterns[20215] = 25'b01001110_11110101_01000011_1;
      patterns[20216] = 25'b01001110_11110110_01000100_1;
      patterns[20217] = 25'b01001110_11110111_01000101_1;
      patterns[20218] = 25'b01001110_11111000_01000110_1;
      patterns[20219] = 25'b01001110_11111001_01000111_1;
      patterns[20220] = 25'b01001110_11111010_01001000_1;
      patterns[20221] = 25'b01001110_11111011_01001001_1;
      patterns[20222] = 25'b01001110_11111100_01001010_1;
      patterns[20223] = 25'b01001110_11111101_01001011_1;
      patterns[20224] = 25'b01001110_11111110_01001100_1;
      patterns[20225] = 25'b01001110_11111111_01001101_1;
      patterns[20226] = 25'b01001111_00000000_01001111_0;
      patterns[20227] = 25'b01001111_00000001_01010000_0;
      patterns[20228] = 25'b01001111_00000010_01010001_0;
      patterns[20229] = 25'b01001111_00000011_01010010_0;
      patterns[20230] = 25'b01001111_00000100_01010011_0;
      patterns[20231] = 25'b01001111_00000101_01010100_0;
      patterns[20232] = 25'b01001111_00000110_01010101_0;
      patterns[20233] = 25'b01001111_00000111_01010110_0;
      patterns[20234] = 25'b01001111_00001000_01010111_0;
      patterns[20235] = 25'b01001111_00001001_01011000_0;
      patterns[20236] = 25'b01001111_00001010_01011001_0;
      patterns[20237] = 25'b01001111_00001011_01011010_0;
      patterns[20238] = 25'b01001111_00001100_01011011_0;
      patterns[20239] = 25'b01001111_00001101_01011100_0;
      patterns[20240] = 25'b01001111_00001110_01011101_0;
      patterns[20241] = 25'b01001111_00001111_01011110_0;
      patterns[20242] = 25'b01001111_00010000_01011111_0;
      patterns[20243] = 25'b01001111_00010001_01100000_0;
      patterns[20244] = 25'b01001111_00010010_01100001_0;
      patterns[20245] = 25'b01001111_00010011_01100010_0;
      patterns[20246] = 25'b01001111_00010100_01100011_0;
      patterns[20247] = 25'b01001111_00010101_01100100_0;
      patterns[20248] = 25'b01001111_00010110_01100101_0;
      patterns[20249] = 25'b01001111_00010111_01100110_0;
      patterns[20250] = 25'b01001111_00011000_01100111_0;
      patterns[20251] = 25'b01001111_00011001_01101000_0;
      patterns[20252] = 25'b01001111_00011010_01101001_0;
      patterns[20253] = 25'b01001111_00011011_01101010_0;
      patterns[20254] = 25'b01001111_00011100_01101011_0;
      patterns[20255] = 25'b01001111_00011101_01101100_0;
      patterns[20256] = 25'b01001111_00011110_01101101_0;
      patterns[20257] = 25'b01001111_00011111_01101110_0;
      patterns[20258] = 25'b01001111_00100000_01101111_0;
      patterns[20259] = 25'b01001111_00100001_01110000_0;
      patterns[20260] = 25'b01001111_00100010_01110001_0;
      patterns[20261] = 25'b01001111_00100011_01110010_0;
      patterns[20262] = 25'b01001111_00100100_01110011_0;
      patterns[20263] = 25'b01001111_00100101_01110100_0;
      patterns[20264] = 25'b01001111_00100110_01110101_0;
      patterns[20265] = 25'b01001111_00100111_01110110_0;
      patterns[20266] = 25'b01001111_00101000_01110111_0;
      patterns[20267] = 25'b01001111_00101001_01111000_0;
      patterns[20268] = 25'b01001111_00101010_01111001_0;
      patterns[20269] = 25'b01001111_00101011_01111010_0;
      patterns[20270] = 25'b01001111_00101100_01111011_0;
      patterns[20271] = 25'b01001111_00101101_01111100_0;
      patterns[20272] = 25'b01001111_00101110_01111101_0;
      patterns[20273] = 25'b01001111_00101111_01111110_0;
      patterns[20274] = 25'b01001111_00110000_01111111_0;
      patterns[20275] = 25'b01001111_00110001_10000000_0;
      patterns[20276] = 25'b01001111_00110010_10000001_0;
      patterns[20277] = 25'b01001111_00110011_10000010_0;
      patterns[20278] = 25'b01001111_00110100_10000011_0;
      patterns[20279] = 25'b01001111_00110101_10000100_0;
      patterns[20280] = 25'b01001111_00110110_10000101_0;
      patterns[20281] = 25'b01001111_00110111_10000110_0;
      patterns[20282] = 25'b01001111_00111000_10000111_0;
      patterns[20283] = 25'b01001111_00111001_10001000_0;
      patterns[20284] = 25'b01001111_00111010_10001001_0;
      patterns[20285] = 25'b01001111_00111011_10001010_0;
      patterns[20286] = 25'b01001111_00111100_10001011_0;
      patterns[20287] = 25'b01001111_00111101_10001100_0;
      patterns[20288] = 25'b01001111_00111110_10001101_0;
      patterns[20289] = 25'b01001111_00111111_10001110_0;
      patterns[20290] = 25'b01001111_01000000_10001111_0;
      patterns[20291] = 25'b01001111_01000001_10010000_0;
      patterns[20292] = 25'b01001111_01000010_10010001_0;
      patterns[20293] = 25'b01001111_01000011_10010010_0;
      patterns[20294] = 25'b01001111_01000100_10010011_0;
      patterns[20295] = 25'b01001111_01000101_10010100_0;
      patterns[20296] = 25'b01001111_01000110_10010101_0;
      patterns[20297] = 25'b01001111_01000111_10010110_0;
      patterns[20298] = 25'b01001111_01001000_10010111_0;
      patterns[20299] = 25'b01001111_01001001_10011000_0;
      patterns[20300] = 25'b01001111_01001010_10011001_0;
      patterns[20301] = 25'b01001111_01001011_10011010_0;
      patterns[20302] = 25'b01001111_01001100_10011011_0;
      patterns[20303] = 25'b01001111_01001101_10011100_0;
      patterns[20304] = 25'b01001111_01001110_10011101_0;
      patterns[20305] = 25'b01001111_01001111_10011110_0;
      patterns[20306] = 25'b01001111_01010000_10011111_0;
      patterns[20307] = 25'b01001111_01010001_10100000_0;
      patterns[20308] = 25'b01001111_01010010_10100001_0;
      patterns[20309] = 25'b01001111_01010011_10100010_0;
      patterns[20310] = 25'b01001111_01010100_10100011_0;
      patterns[20311] = 25'b01001111_01010101_10100100_0;
      patterns[20312] = 25'b01001111_01010110_10100101_0;
      patterns[20313] = 25'b01001111_01010111_10100110_0;
      patterns[20314] = 25'b01001111_01011000_10100111_0;
      patterns[20315] = 25'b01001111_01011001_10101000_0;
      patterns[20316] = 25'b01001111_01011010_10101001_0;
      patterns[20317] = 25'b01001111_01011011_10101010_0;
      patterns[20318] = 25'b01001111_01011100_10101011_0;
      patterns[20319] = 25'b01001111_01011101_10101100_0;
      patterns[20320] = 25'b01001111_01011110_10101101_0;
      patterns[20321] = 25'b01001111_01011111_10101110_0;
      patterns[20322] = 25'b01001111_01100000_10101111_0;
      patterns[20323] = 25'b01001111_01100001_10110000_0;
      patterns[20324] = 25'b01001111_01100010_10110001_0;
      patterns[20325] = 25'b01001111_01100011_10110010_0;
      patterns[20326] = 25'b01001111_01100100_10110011_0;
      patterns[20327] = 25'b01001111_01100101_10110100_0;
      patterns[20328] = 25'b01001111_01100110_10110101_0;
      patterns[20329] = 25'b01001111_01100111_10110110_0;
      patterns[20330] = 25'b01001111_01101000_10110111_0;
      patterns[20331] = 25'b01001111_01101001_10111000_0;
      patterns[20332] = 25'b01001111_01101010_10111001_0;
      patterns[20333] = 25'b01001111_01101011_10111010_0;
      patterns[20334] = 25'b01001111_01101100_10111011_0;
      patterns[20335] = 25'b01001111_01101101_10111100_0;
      patterns[20336] = 25'b01001111_01101110_10111101_0;
      patterns[20337] = 25'b01001111_01101111_10111110_0;
      patterns[20338] = 25'b01001111_01110000_10111111_0;
      patterns[20339] = 25'b01001111_01110001_11000000_0;
      patterns[20340] = 25'b01001111_01110010_11000001_0;
      patterns[20341] = 25'b01001111_01110011_11000010_0;
      patterns[20342] = 25'b01001111_01110100_11000011_0;
      patterns[20343] = 25'b01001111_01110101_11000100_0;
      patterns[20344] = 25'b01001111_01110110_11000101_0;
      patterns[20345] = 25'b01001111_01110111_11000110_0;
      patterns[20346] = 25'b01001111_01111000_11000111_0;
      patterns[20347] = 25'b01001111_01111001_11001000_0;
      patterns[20348] = 25'b01001111_01111010_11001001_0;
      patterns[20349] = 25'b01001111_01111011_11001010_0;
      patterns[20350] = 25'b01001111_01111100_11001011_0;
      patterns[20351] = 25'b01001111_01111101_11001100_0;
      patterns[20352] = 25'b01001111_01111110_11001101_0;
      patterns[20353] = 25'b01001111_01111111_11001110_0;
      patterns[20354] = 25'b01001111_10000000_11001111_0;
      patterns[20355] = 25'b01001111_10000001_11010000_0;
      patterns[20356] = 25'b01001111_10000010_11010001_0;
      patterns[20357] = 25'b01001111_10000011_11010010_0;
      patterns[20358] = 25'b01001111_10000100_11010011_0;
      patterns[20359] = 25'b01001111_10000101_11010100_0;
      patterns[20360] = 25'b01001111_10000110_11010101_0;
      patterns[20361] = 25'b01001111_10000111_11010110_0;
      patterns[20362] = 25'b01001111_10001000_11010111_0;
      patterns[20363] = 25'b01001111_10001001_11011000_0;
      patterns[20364] = 25'b01001111_10001010_11011001_0;
      patterns[20365] = 25'b01001111_10001011_11011010_0;
      patterns[20366] = 25'b01001111_10001100_11011011_0;
      patterns[20367] = 25'b01001111_10001101_11011100_0;
      patterns[20368] = 25'b01001111_10001110_11011101_0;
      patterns[20369] = 25'b01001111_10001111_11011110_0;
      patterns[20370] = 25'b01001111_10010000_11011111_0;
      patterns[20371] = 25'b01001111_10010001_11100000_0;
      patterns[20372] = 25'b01001111_10010010_11100001_0;
      patterns[20373] = 25'b01001111_10010011_11100010_0;
      patterns[20374] = 25'b01001111_10010100_11100011_0;
      patterns[20375] = 25'b01001111_10010101_11100100_0;
      patterns[20376] = 25'b01001111_10010110_11100101_0;
      patterns[20377] = 25'b01001111_10010111_11100110_0;
      patterns[20378] = 25'b01001111_10011000_11100111_0;
      patterns[20379] = 25'b01001111_10011001_11101000_0;
      patterns[20380] = 25'b01001111_10011010_11101001_0;
      patterns[20381] = 25'b01001111_10011011_11101010_0;
      patterns[20382] = 25'b01001111_10011100_11101011_0;
      patterns[20383] = 25'b01001111_10011101_11101100_0;
      patterns[20384] = 25'b01001111_10011110_11101101_0;
      patterns[20385] = 25'b01001111_10011111_11101110_0;
      patterns[20386] = 25'b01001111_10100000_11101111_0;
      patterns[20387] = 25'b01001111_10100001_11110000_0;
      patterns[20388] = 25'b01001111_10100010_11110001_0;
      patterns[20389] = 25'b01001111_10100011_11110010_0;
      patterns[20390] = 25'b01001111_10100100_11110011_0;
      patterns[20391] = 25'b01001111_10100101_11110100_0;
      patterns[20392] = 25'b01001111_10100110_11110101_0;
      patterns[20393] = 25'b01001111_10100111_11110110_0;
      patterns[20394] = 25'b01001111_10101000_11110111_0;
      patterns[20395] = 25'b01001111_10101001_11111000_0;
      patterns[20396] = 25'b01001111_10101010_11111001_0;
      patterns[20397] = 25'b01001111_10101011_11111010_0;
      patterns[20398] = 25'b01001111_10101100_11111011_0;
      patterns[20399] = 25'b01001111_10101101_11111100_0;
      patterns[20400] = 25'b01001111_10101110_11111101_0;
      patterns[20401] = 25'b01001111_10101111_11111110_0;
      patterns[20402] = 25'b01001111_10110000_11111111_0;
      patterns[20403] = 25'b01001111_10110001_00000000_1;
      patterns[20404] = 25'b01001111_10110010_00000001_1;
      patterns[20405] = 25'b01001111_10110011_00000010_1;
      patterns[20406] = 25'b01001111_10110100_00000011_1;
      patterns[20407] = 25'b01001111_10110101_00000100_1;
      patterns[20408] = 25'b01001111_10110110_00000101_1;
      patterns[20409] = 25'b01001111_10110111_00000110_1;
      patterns[20410] = 25'b01001111_10111000_00000111_1;
      patterns[20411] = 25'b01001111_10111001_00001000_1;
      patterns[20412] = 25'b01001111_10111010_00001001_1;
      patterns[20413] = 25'b01001111_10111011_00001010_1;
      patterns[20414] = 25'b01001111_10111100_00001011_1;
      patterns[20415] = 25'b01001111_10111101_00001100_1;
      patterns[20416] = 25'b01001111_10111110_00001101_1;
      patterns[20417] = 25'b01001111_10111111_00001110_1;
      patterns[20418] = 25'b01001111_11000000_00001111_1;
      patterns[20419] = 25'b01001111_11000001_00010000_1;
      patterns[20420] = 25'b01001111_11000010_00010001_1;
      patterns[20421] = 25'b01001111_11000011_00010010_1;
      patterns[20422] = 25'b01001111_11000100_00010011_1;
      patterns[20423] = 25'b01001111_11000101_00010100_1;
      patterns[20424] = 25'b01001111_11000110_00010101_1;
      patterns[20425] = 25'b01001111_11000111_00010110_1;
      patterns[20426] = 25'b01001111_11001000_00010111_1;
      patterns[20427] = 25'b01001111_11001001_00011000_1;
      patterns[20428] = 25'b01001111_11001010_00011001_1;
      patterns[20429] = 25'b01001111_11001011_00011010_1;
      patterns[20430] = 25'b01001111_11001100_00011011_1;
      patterns[20431] = 25'b01001111_11001101_00011100_1;
      patterns[20432] = 25'b01001111_11001110_00011101_1;
      patterns[20433] = 25'b01001111_11001111_00011110_1;
      patterns[20434] = 25'b01001111_11010000_00011111_1;
      patterns[20435] = 25'b01001111_11010001_00100000_1;
      patterns[20436] = 25'b01001111_11010010_00100001_1;
      patterns[20437] = 25'b01001111_11010011_00100010_1;
      patterns[20438] = 25'b01001111_11010100_00100011_1;
      patterns[20439] = 25'b01001111_11010101_00100100_1;
      patterns[20440] = 25'b01001111_11010110_00100101_1;
      patterns[20441] = 25'b01001111_11010111_00100110_1;
      patterns[20442] = 25'b01001111_11011000_00100111_1;
      patterns[20443] = 25'b01001111_11011001_00101000_1;
      patterns[20444] = 25'b01001111_11011010_00101001_1;
      patterns[20445] = 25'b01001111_11011011_00101010_1;
      patterns[20446] = 25'b01001111_11011100_00101011_1;
      patterns[20447] = 25'b01001111_11011101_00101100_1;
      patterns[20448] = 25'b01001111_11011110_00101101_1;
      patterns[20449] = 25'b01001111_11011111_00101110_1;
      patterns[20450] = 25'b01001111_11100000_00101111_1;
      patterns[20451] = 25'b01001111_11100001_00110000_1;
      patterns[20452] = 25'b01001111_11100010_00110001_1;
      patterns[20453] = 25'b01001111_11100011_00110010_1;
      patterns[20454] = 25'b01001111_11100100_00110011_1;
      patterns[20455] = 25'b01001111_11100101_00110100_1;
      patterns[20456] = 25'b01001111_11100110_00110101_1;
      patterns[20457] = 25'b01001111_11100111_00110110_1;
      patterns[20458] = 25'b01001111_11101000_00110111_1;
      patterns[20459] = 25'b01001111_11101001_00111000_1;
      patterns[20460] = 25'b01001111_11101010_00111001_1;
      patterns[20461] = 25'b01001111_11101011_00111010_1;
      patterns[20462] = 25'b01001111_11101100_00111011_1;
      patterns[20463] = 25'b01001111_11101101_00111100_1;
      patterns[20464] = 25'b01001111_11101110_00111101_1;
      patterns[20465] = 25'b01001111_11101111_00111110_1;
      patterns[20466] = 25'b01001111_11110000_00111111_1;
      patterns[20467] = 25'b01001111_11110001_01000000_1;
      patterns[20468] = 25'b01001111_11110010_01000001_1;
      patterns[20469] = 25'b01001111_11110011_01000010_1;
      patterns[20470] = 25'b01001111_11110100_01000011_1;
      patterns[20471] = 25'b01001111_11110101_01000100_1;
      patterns[20472] = 25'b01001111_11110110_01000101_1;
      patterns[20473] = 25'b01001111_11110111_01000110_1;
      patterns[20474] = 25'b01001111_11111000_01000111_1;
      patterns[20475] = 25'b01001111_11111001_01001000_1;
      patterns[20476] = 25'b01001111_11111010_01001001_1;
      patterns[20477] = 25'b01001111_11111011_01001010_1;
      patterns[20478] = 25'b01001111_11111100_01001011_1;
      patterns[20479] = 25'b01001111_11111101_01001100_1;
      patterns[20480] = 25'b01001111_11111110_01001101_1;
      patterns[20481] = 25'b01001111_11111111_01001110_1;
      patterns[20482] = 25'b01010000_00000000_01010000_0;
      patterns[20483] = 25'b01010000_00000001_01010001_0;
      patterns[20484] = 25'b01010000_00000010_01010010_0;
      patterns[20485] = 25'b01010000_00000011_01010011_0;
      patterns[20486] = 25'b01010000_00000100_01010100_0;
      patterns[20487] = 25'b01010000_00000101_01010101_0;
      patterns[20488] = 25'b01010000_00000110_01010110_0;
      patterns[20489] = 25'b01010000_00000111_01010111_0;
      patterns[20490] = 25'b01010000_00001000_01011000_0;
      patterns[20491] = 25'b01010000_00001001_01011001_0;
      patterns[20492] = 25'b01010000_00001010_01011010_0;
      patterns[20493] = 25'b01010000_00001011_01011011_0;
      patterns[20494] = 25'b01010000_00001100_01011100_0;
      patterns[20495] = 25'b01010000_00001101_01011101_0;
      patterns[20496] = 25'b01010000_00001110_01011110_0;
      patterns[20497] = 25'b01010000_00001111_01011111_0;
      patterns[20498] = 25'b01010000_00010000_01100000_0;
      patterns[20499] = 25'b01010000_00010001_01100001_0;
      patterns[20500] = 25'b01010000_00010010_01100010_0;
      patterns[20501] = 25'b01010000_00010011_01100011_0;
      patterns[20502] = 25'b01010000_00010100_01100100_0;
      patterns[20503] = 25'b01010000_00010101_01100101_0;
      patterns[20504] = 25'b01010000_00010110_01100110_0;
      patterns[20505] = 25'b01010000_00010111_01100111_0;
      patterns[20506] = 25'b01010000_00011000_01101000_0;
      patterns[20507] = 25'b01010000_00011001_01101001_0;
      patterns[20508] = 25'b01010000_00011010_01101010_0;
      patterns[20509] = 25'b01010000_00011011_01101011_0;
      patterns[20510] = 25'b01010000_00011100_01101100_0;
      patterns[20511] = 25'b01010000_00011101_01101101_0;
      patterns[20512] = 25'b01010000_00011110_01101110_0;
      patterns[20513] = 25'b01010000_00011111_01101111_0;
      patterns[20514] = 25'b01010000_00100000_01110000_0;
      patterns[20515] = 25'b01010000_00100001_01110001_0;
      patterns[20516] = 25'b01010000_00100010_01110010_0;
      patterns[20517] = 25'b01010000_00100011_01110011_0;
      patterns[20518] = 25'b01010000_00100100_01110100_0;
      patterns[20519] = 25'b01010000_00100101_01110101_0;
      patterns[20520] = 25'b01010000_00100110_01110110_0;
      patterns[20521] = 25'b01010000_00100111_01110111_0;
      patterns[20522] = 25'b01010000_00101000_01111000_0;
      patterns[20523] = 25'b01010000_00101001_01111001_0;
      patterns[20524] = 25'b01010000_00101010_01111010_0;
      patterns[20525] = 25'b01010000_00101011_01111011_0;
      patterns[20526] = 25'b01010000_00101100_01111100_0;
      patterns[20527] = 25'b01010000_00101101_01111101_0;
      patterns[20528] = 25'b01010000_00101110_01111110_0;
      patterns[20529] = 25'b01010000_00101111_01111111_0;
      patterns[20530] = 25'b01010000_00110000_10000000_0;
      patterns[20531] = 25'b01010000_00110001_10000001_0;
      patterns[20532] = 25'b01010000_00110010_10000010_0;
      patterns[20533] = 25'b01010000_00110011_10000011_0;
      patterns[20534] = 25'b01010000_00110100_10000100_0;
      patterns[20535] = 25'b01010000_00110101_10000101_0;
      patterns[20536] = 25'b01010000_00110110_10000110_0;
      patterns[20537] = 25'b01010000_00110111_10000111_0;
      patterns[20538] = 25'b01010000_00111000_10001000_0;
      patterns[20539] = 25'b01010000_00111001_10001001_0;
      patterns[20540] = 25'b01010000_00111010_10001010_0;
      patterns[20541] = 25'b01010000_00111011_10001011_0;
      patterns[20542] = 25'b01010000_00111100_10001100_0;
      patterns[20543] = 25'b01010000_00111101_10001101_0;
      patterns[20544] = 25'b01010000_00111110_10001110_0;
      patterns[20545] = 25'b01010000_00111111_10001111_0;
      patterns[20546] = 25'b01010000_01000000_10010000_0;
      patterns[20547] = 25'b01010000_01000001_10010001_0;
      patterns[20548] = 25'b01010000_01000010_10010010_0;
      patterns[20549] = 25'b01010000_01000011_10010011_0;
      patterns[20550] = 25'b01010000_01000100_10010100_0;
      patterns[20551] = 25'b01010000_01000101_10010101_0;
      patterns[20552] = 25'b01010000_01000110_10010110_0;
      patterns[20553] = 25'b01010000_01000111_10010111_0;
      patterns[20554] = 25'b01010000_01001000_10011000_0;
      patterns[20555] = 25'b01010000_01001001_10011001_0;
      patterns[20556] = 25'b01010000_01001010_10011010_0;
      patterns[20557] = 25'b01010000_01001011_10011011_0;
      patterns[20558] = 25'b01010000_01001100_10011100_0;
      patterns[20559] = 25'b01010000_01001101_10011101_0;
      patterns[20560] = 25'b01010000_01001110_10011110_0;
      patterns[20561] = 25'b01010000_01001111_10011111_0;
      patterns[20562] = 25'b01010000_01010000_10100000_0;
      patterns[20563] = 25'b01010000_01010001_10100001_0;
      patterns[20564] = 25'b01010000_01010010_10100010_0;
      patterns[20565] = 25'b01010000_01010011_10100011_0;
      patterns[20566] = 25'b01010000_01010100_10100100_0;
      patterns[20567] = 25'b01010000_01010101_10100101_0;
      patterns[20568] = 25'b01010000_01010110_10100110_0;
      patterns[20569] = 25'b01010000_01010111_10100111_0;
      patterns[20570] = 25'b01010000_01011000_10101000_0;
      patterns[20571] = 25'b01010000_01011001_10101001_0;
      patterns[20572] = 25'b01010000_01011010_10101010_0;
      patterns[20573] = 25'b01010000_01011011_10101011_0;
      patterns[20574] = 25'b01010000_01011100_10101100_0;
      patterns[20575] = 25'b01010000_01011101_10101101_0;
      patterns[20576] = 25'b01010000_01011110_10101110_0;
      patterns[20577] = 25'b01010000_01011111_10101111_0;
      patterns[20578] = 25'b01010000_01100000_10110000_0;
      patterns[20579] = 25'b01010000_01100001_10110001_0;
      patterns[20580] = 25'b01010000_01100010_10110010_0;
      patterns[20581] = 25'b01010000_01100011_10110011_0;
      patterns[20582] = 25'b01010000_01100100_10110100_0;
      patterns[20583] = 25'b01010000_01100101_10110101_0;
      patterns[20584] = 25'b01010000_01100110_10110110_0;
      patterns[20585] = 25'b01010000_01100111_10110111_0;
      patterns[20586] = 25'b01010000_01101000_10111000_0;
      patterns[20587] = 25'b01010000_01101001_10111001_0;
      patterns[20588] = 25'b01010000_01101010_10111010_0;
      patterns[20589] = 25'b01010000_01101011_10111011_0;
      patterns[20590] = 25'b01010000_01101100_10111100_0;
      patterns[20591] = 25'b01010000_01101101_10111101_0;
      patterns[20592] = 25'b01010000_01101110_10111110_0;
      patterns[20593] = 25'b01010000_01101111_10111111_0;
      patterns[20594] = 25'b01010000_01110000_11000000_0;
      patterns[20595] = 25'b01010000_01110001_11000001_0;
      patterns[20596] = 25'b01010000_01110010_11000010_0;
      patterns[20597] = 25'b01010000_01110011_11000011_0;
      patterns[20598] = 25'b01010000_01110100_11000100_0;
      patterns[20599] = 25'b01010000_01110101_11000101_0;
      patterns[20600] = 25'b01010000_01110110_11000110_0;
      patterns[20601] = 25'b01010000_01110111_11000111_0;
      patterns[20602] = 25'b01010000_01111000_11001000_0;
      patterns[20603] = 25'b01010000_01111001_11001001_0;
      patterns[20604] = 25'b01010000_01111010_11001010_0;
      patterns[20605] = 25'b01010000_01111011_11001011_0;
      patterns[20606] = 25'b01010000_01111100_11001100_0;
      patterns[20607] = 25'b01010000_01111101_11001101_0;
      patterns[20608] = 25'b01010000_01111110_11001110_0;
      patterns[20609] = 25'b01010000_01111111_11001111_0;
      patterns[20610] = 25'b01010000_10000000_11010000_0;
      patterns[20611] = 25'b01010000_10000001_11010001_0;
      patterns[20612] = 25'b01010000_10000010_11010010_0;
      patterns[20613] = 25'b01010000_10000011_11010011_0;
      patterns[20614] = 25'b01010000_10000100_11010100_0;
      patterns[20615] = 25'b01010000_10000101_11010101_0;
      patterns[20616] = 25'b01010000_10000110_11010110_0;
      patterns[20617] = 25'b01010000_10000111_11010111_0;
      patterns[20618] = 25'b01010000_10001000_11011000_0;
      patterns[20619] = 25'b01010000_10001001_11011001_0;
      patterns[20620] = 25'b01010000_10001010_11011010_0;
      patterns[20621] = 25'b01010000_10001011_11011011_0;
      patterns[20622] = 25'b01010000_10001100_11011100_0;
      patterns[20623] = 25'b01010000_10001101_11011101_0;
      patterns[20624] = 25'b01010000_10001110_11011110_0;
      patterns[20625] = 25'b01010000_10001111_11011111_0;
      patterns[20626] = 25'b01010000_10010000_11100000_0;
      patterns[20627] = 25'b01010000_10010001_11100001_0;
      patterns[20628] = 25'b01010000_10010010_11100010_0;
      patterns[20629] = 25'b01010000_10010011_11100011_0;
      patterns[20630] = 25'b01010000_10010100_11100100_0;
      patterns[20631] = 25'b01010000_10010101_11100101_0;
      patterns[20632] = 25'b01010000_10010110_11100110_0;
      patterns[20633] = 25'b01010000_10010111_11100111_0;
      patterns[20634] = 25'b01010000_10011000_11101000_0;
      patterns[20635] = 25'b01010000_10011001_11101001_0;
      patterns[20636] = 25'b01010000_10011010_11101010_0;
      patterns[20637] = 25'b01010000_10011011_11101011_0;
      patterns[20638] = 25'b01010000_10011100_11101100_0;
      patterns[20639] = 25'b01010000_10011101_11101101_0;
      patterns[20640] = 25'b01010000_10011110_11101110_0;
      patterns[20641] = 25'b01010000_10011111_11101111_0;
      patterns[20642] = 25'b01010000_10100000_11110000_0;
      patterns[20643] = 25'b01010000_10100001_11110001_0;
      patterns[20644] = 25'b01010000_10100010_11110010_0;
      patterns[20645] = 25'b01010000_10100011_11110011_0;
      patterns[20646] = 25'b01010000_10100100_11110100_0;
      patterns[20647] = 25'b01010000_10100101_11110101_0;
      patterns[20648] = 25'b01010000_10100110_11110110_0;
      patterns[20649] = 25'b01010000_10100111_11110111_0;
      patterns[20650] = 25'b01010000_10101000_11111000_0;
      patterns[20651] = 25'b01010000_10101001_11111001_0;
      patterns[20652] = 25'b01010000_10101010_11111010_0;
      patterns[20653] = 25'b01010000_10101011_11111011_0;
      patterns[20654] = 25'b01010000_10101100_11111100_0;
      patterns[20655] = 25'b01010000_10101101_11111101_0;
      patterns[20656] = 25'b01010000_10101110_11111110_0;
      patterns[20657] = 25'b01010000_10101111_11111111_0;
      patterns[20658] = 25'b01010000_10110000_00000000_1;
      patterns[20659] = 25'b01010000_10110001_00000001_1;
      patterns[20660] = 25'b01010000_10110010_00000010_1;
      patterns[20661] = 25'b01010000_10110011_00000011_1;
      patterns[20662] = 25'b01010000_10110100_00000100_1;
      patterns[20663] = 25'b01010000_10110101_00000101_1;
      patterns[20664] = 25'b01010000_10110110_00000110_1;
      patterns[20665] = 25'b01010000_10110111_00000111_1;
      patterns[20666] = 25'b01010000_10111000_00001000_1;
      patterns[20667] = 25'b01010000_10111001_00001001_1;
      patterns[20668] = 25'b01010000_10111010_00001010_1;
      patterns[20669] = 25'b01010000_10111011_00001011_1;
      patterns[20670] = 25'b01010000_10111100_00001100_1;
      patterns[20671] = 25'b01010000_10111101_00001101_1;
      patterns[20672] = 25'b01010000_10111110_00001110_1;
      patterns[20673] = 25'b01010000_10111111_00001111_1;
      patterns[20674] = 25'b01010000_11000000_00010000_1;
      patterns[20675] = 25'b01010000_11000001_00010001_1;
      patterns[20676] = 25'b01010000_11000010_00010010_1;
      patterns[20677] = 25'b01010000_11000011_00010011_1;
      patterns[20678] = 25'b01010000_11000100_00010100_1;
      patterns[20679] = 25'b01010000_11000101_00010101_1;
      patterns[20680] = 25'b01010000_11000110_00010110_1;
      patterns[20681] = 25'b01010000_11000111_00010111_1;
      patterns[20682] = 25'b01010000_11001000_00011000_1;
      patterns[20683] = 25'b01010000_11001001_00011001_1;
      patterns[20684] = 25'b01010000_11001010_00011010_1;
      patterns[20685] = 25'b01010000_11001011_00011011_1;
      patterns[20686] = 25'b01010000_11001100_00011100_1;
      patterns[20687] = 25'b01010000_11001101_00011101_1;
      patterns[20688] = 25'b01010000_11001110_00011110_1;
      patterns[20689] = 25'b01010000_11001111_00011111_1;
      patterns[20690] = 25'b01010000_11010000_00100000_1;
      patterns[20691] = 25'b01010000_11010001_00100001_1;
      patterns[20692] = 25'b01010000_11010010_00100010_1;
      patterns[20693] = 25'b01010000_11010011_00100011_1;
      patterns[20694] = 25'b01010000_11010100_00100100_1;
      patterns[20695] = 25'b01010000_11010101_00100101_1;
      patterns[20696] = 25'b01010000_11010110_00100110_1;
      patterns[20697] = 25'b01010000_11010111_00100111_1;
      patterns[20698] = 25'b01010000_11011000_00101000_1;
      patterns[20699] = 25'b01010000_11011001_00101001_1;
      patterns[20700] = 25'b01010000_11011010_00101010_1;
      patterns[20701] = 25'b01010000_11011011_00101011_1;
      patterns[20702] = 25'b01010000_11011100_00101100_1;
      patterns[20703] = 25'b01010000_11011101_00101101_1;
      patterns[20704] = 25'b01010000_11011110_00101110_1;
      patterns[20705] = 25'b01010000_11011111_00101111_1;
      patterns[20706] = 25'b01010000_11100000_00110000_1;
      patterns[20707] = 25'b01010000_11100001_00110001_1;
      patterns[20708] = 25'b01010000_11100010_00110010_1;
      patterns[20709] = 25'b01010000_11100011_00110011_1;
      patterns[20710] = 25'b01010000_11100100_00110100_1;
      patterns[20711] = 25'b01010000_11100101_00110101_1;
      patterns[20712] = 25'b01010000_11100110_00110110_1;
      patterns[20713] = 25'b01010000_11100111_00110111_1;
      patterns[20714] = 25'b01010000_11101000_00111000_1;
      patterns[20715] = 25'b01010000_11101001_00111001_1;
      patterns[20716] = 25'b01010000_11101010_00111010_1;
      patterns[20717] = 25'b01010000_11101011_00111011_1;
      patterns[20718] = 25'b01010000_11101100_00111100_1;
      patterns[20719] = 25'b01010000_11101101_00111101_1;
      patterns[20720] = 25'b01010000_11101110_00111110_1;
      patterns[20721] = 25'b01010000_11101111_00111111_1;
      patterns[20722] = 25'b01010000_11110000_01000000_1;
      patterns[20723] = 25'b01010000_11110001_01000001_1;
      patterns[20724] = 25'b01010000_11110010_01000010_1;
      patterns[20725] = 25'b01010000_11110011_01000011_1;
      patterns[20726] = 25'b01010000_11110100_01000100_1;
      patterns[20727] = 25'b01010000_11110101_01000101_1;
      patterns[20728] = 25'b01010000_11110110_01000110_1;
      patterns[20729] = 25'b01010000_11110111_01000111_1;
      patterns[20730] = 25'b01010000_11111000_01001000_1;
      patterns[20731] = 25'b01010000_11111001_01001001_1;
      patterns[20732] = 25'b01010000_11111010_01001010_1;
      patterns[20733] = 25'b01010000_11111011_01001011_1;
      patterns[20734] = 25'b01010000_11111100_01001100_1;
      patterns[20735] = 25'b01010000_11111101_01001101_1;
      patterns[20736] = 25'b01010000_11111110_01001110_1;
      patterns[20737] = 25'b01010000_11111111_01001111_1;
      patterns[20738] = 25'b01010001_00000000_01010001_0;
      patterns[20739] = 25'b01010001_00000001_01010010_0;
      patterns[20740] = 25'b01010001_00000010_01010011_0;
      patterns[20741] = 25'b01010001_00000011_01010100_0;
      patterns[20742] = 25'b01010001_00000100_01010101_0;
      patterns[20743] = 25'b01010001_00000101_01010110_0;
      patterns[20744] = 25'b01010001_00000110_01010111_0;
      patterns[20745] = 25'b01010001_00000111_01011000_0;
      patterns[20746] = 25'b01010001_00001000_01011001_0;
      patterns[20747] = 25'b01010001_00001001_01011010_0;
      patterns[20748] = 25'b01010001_00001010_01011011_0;
      patterns[20749] = 25'b01010001_00001011_01011100_0;
      patterns[20750] = 25'b01010001_00001100_01011101_0;
      patterns[20751] = 25'b01010001_00001101_01011110_0;
      patterns[20752] = 25'b01010001_00001110_01011111_0;
      patterns[20753] = 25'b01010001_00001111_01100000_0;
      patterns[20754] = 25'b01010001_00010000_01100001_0;
      patterns[20755] = 25'b01010001_00010001_01100010_0;
      patterns[20756] = 25'b01010001_00010010_01100011_0;
      patterns[20757] = 25'b01010001_00010011_01100100_0;
      patterns[20758] = 25'b01010001_00010100_01100101_0;
      patterns[20759] = 25'b01010001_00010101_01100110_0;
      patterns[20760] = 25'b01010001_00010110_01100111_0;
      patterns[20761] = 25'b01010001_00010111_01101000_0;
      patterns[20762] = 25'b01010001_00011000_01101001_0;
      patterns[20763] = 25'b01010001_00011001_01101010_0;
      patterns[20764] = 25'b01010001_00011010_01101011_0;
      patterns[20765] = 25'b01010001_00011011_01101100_0;
      patterns[20766] = 25'b01010001_00011100_01101101_0;
      patterns[20767] = 25'b01010001_00011101_01101110_0;
      patterns[20768] = 25'b01010001_00011110_01101111_0;
      patterns[20769] = 25'b01010001_00011111_01110000_0;
      patterns[20770] = 25'b01010001_00100000_01110001_0;
      patterns[20771] = 25'b01010001_00100001_01110010_0;
      patterns[20772] = 25'b01010001_00100010_01110011_0;
      patterns[20773] = 25'b01010001_00100011_01110100_0;
      patterns[20774] = 25'b01010001_00100100_01110101_0;
      patterns[20775] = 25'b01010001_00100101_01110110_0;
      patterns[20776] = 25'b01010001_00100110_01110111_0;
      patterns[20777] = 25'b01010001_00100111_01111000_0;
      patterns[20778] = 25'b01010001_00101000_01111001_0;
      patterns[20779] = 25'b01010001_00101001_01111010_0;
      patterns[20780] = 25'b01010001_00101010_01111011_0;
      patterns[20781] = 25'b01010001_00101011_01111100_0;
      patterns[20782] = 25'b01010001_00101100_01111101_0;
      patterns[20783] = 25'b01010001_00101101_01111110_0;
      patterns[20784] = 25'b01010001_00101110_01111111_0;
      patterns[20785] = 25'b01010001_00101111_10000000_0;
      patterns[20786] = 25'b01010001_00110000_10000001_0;
      patterns[20787] = 25'b01010001_00110001_10000010_0;
      patterns[20788] = 25'b01010001_00110010_10000011_0;
      patterns[20789] = 25'b01010001_00110011_10000100_0;
      patterns[20790] = 25'b01010001_00110100_10000101_0;
      patterns[20791] = 25'b01010001_00110101_10000110_0;
      patterns[20792] = 25'b01010001_00110110_10000111_0;
      patterns[20793] = 25'b01010001_00110111_10001000_0;
      patterns[20794] = 25'b01010001_00111000_10001001_0;
      patterns[20795] = 25'b01010001_00111001_10001010_0;
      patterns[20796] = 25'b01010001_00111010_10001011_0;
      patterns[20797] = 25'b01010001_00111011_10001100_0;
      patterns[20798] = 25'b01010001_00111100_10001101_0;
      patterns[20799] = 25'b01010001_00111101_10001110_0;
      patterns[20800] = 25'b01010001_00111110_10001111_0;
      patterns[20801] = 25'b01010001_00111111_10010000_0;
      patterns[20802] = 25'b01010001_01000000_10010001_0;
      patterns[20803] = 25'b01010001_01000001_10010010_0;
      patterns[20804] = 25'b01010001_01000010_10010011_0;
      patterns[20805] = 25'b01010001_01000011_10010100_0;
      patterns[20806] = 25'b01010001_01000100_10010101_0;
      patterns[20807] = 25'b01010001_01000101_10010110_0;
      patterns[20808] = 25'b01010001_01000110_10010111_0;
      patterns[20809] = 25'b01010001_01000111_10011000_0;
      patterns[20810] = 25'b01010001_01001000_10011001_0;
      patterns[20811] = 25'b01010001_01001001_10011010_0;
      patterns[20812] = 25'b01010001_01001010_10011011_0;
      patterns[20813] = 25'b01010001_01001011_10011100_0;
      patterns[20814] = 25'b01010001_01001100_10011101_0;
      patterns[20815] = 25'b01010001_01001101_10011110_0;
      patterns[20816] = 25'b01010001_01001110_10011111_0;
      patterns[20817] = 25'b01010001_01001111_10100000_0;
      patterns[20818] = 25'b01010001_01010000_10100001_0;
      patterns[20819] = 25'b01010001_01010001_10100010_0;
      patterns[20820] = 25'b01010001_01010010_10100011_0;
      patterns[20821] = 25'b01010001_01010011_10100100_0;
      patterns[20822] = 25'b01010001_01010100_10100101_0;
      patterns[20823] = 25'b01010001_01010101_10100110_0;
      patterns[20824] = 25'b01010001_01010110_10100111_0;
      patterns[20825] = 25'b01010001_01010111_10101000_0;
      patterns[20826] = 25'b01010001_01011000_10101001_0;
      patterns[20827] = 25'b01010001_01011001_10101010_0;
      patterns[20828] = 25'b01010001_01011010_10101011_0;
      patterns[20829] = 25'b01010001_01011011_10101100_0;
      patterns[20830] = 25'b01010001_01011100_10101101_0;
      patterns[20831] = 25'b01010001_01011101_10101110_0;
      patterns[20832] = 25'b01010001_01011110_10101111_0;
      patterns[20833] = 25'b01010001_01011111_10110000_0;
      patterns[20834] = 25'b01010001_01100000_10110001_0;
      patterns[20835] = 25'b01010001_01100001_10110010_0;
      patterns[20836] = 25'b01010001_01100010_10110011_0;
      patterns[20837] = 25'b01010001_01100011_10110100_0;
      patterns[20838] = 25'b01010001_01100100_10110101_0;
      patterns[20839] = 25'b01010001_01100101_10110110_0;
      patterns[20840] = 25'b01010001_01100110_10110111_0;
      patterns[20841] = 25'b01010001_01100111_10111000_0;
      patterns[20842] = 25'b01010001_01101000_10111001_0;
      patterns[20843] = 25'b01010001_01101001_10111010_0;
      patterns[20844] = 25'b01010001_01101010_10111011_0;
      patterns[20845] = 25'b01010001_01101011_10111100_0;
      patterns[20846] = 25'b01010001_01101100_10111101_0;
      patterns[20847] = 25'b01010001_01101101_10111110_0;
      patterns[20848] = 25'b01010001_01101110_10111111_0;
      patterns[20849] = 25'b01010001_01101111_11000000_0;
      patterns[20850] = 25'b01010001_01110000_11000001_0;
      patterns[20851] = 25'b01010001_01110001_11000010_0;
      patterns[20852] = 25'b01010001_01110010_11000011_0;
      patterns[20853] = 25'b01010001_01110011_11000100_0;
      patterns[20854] = 25'b01010001_01110100_11000101_0;
      patterns[20855] = 25'b01010001_01110101_11000110_0;
      patterns[20856] = 25'b01010001_01110110_11000111_0;
      patterns[20857] = 25'b01010001_01110111_11001000_0;
      patterns[20858] = 25'b01010001_01111000_11001001_0;
      patterns[20859] = 25'b01010001_01111001_11001010_0;
      patterns[20860] = 25'b01010001_01111010_11001011_0;
      patterns[20861] = 25'b01010001_01111011_11001100_0;
      patterns[20862] = 25'b01010001_01111100_11001101_0;
      patterns[20863] = 25'b01010001_01111101_11001110_0;
      patterns[20864] = 25'b01010001_01111110_11001111_0;
      patterns[20865] = 25'b01010001_01111111_11010000_0;
      patterns[20866] = 25'b01010001_10000000_11010001_0;
      patterns[20867] = 25'b01010001_10000001_11010010_0;
      patterns[20868] = 25'b01010001_10000010_11010011_0;
      patterns[20869] = 25'b01010001_10000011_11010100_0;
      patterns[20870] = 25'b01010001_10000100_11010101_0;
      patterns[20871] = 25'b01010001_10000101_11010110_0;
      patterns[20872] = 25'b01010001_10000110_11010111_0;
      patterns[20873] = 25'b01010001_10000111_11011000_0;
      patterns[20874] = 25'b01010001_10001000_11011001_0;
      patterns[20875] = 25'b01010001_10001001_11011010_0;
      patterns[20876] = 25'b01010001_10001010_11011011_0;
      patterns[20877] = 25'b01010001_10001011_11011100_0;
      patterns[20878] = 25'b01010001_10001100_11011101_0;
      patterns[20879] = 25'b01010001_10001101_11011110_0;
      patterns[20880] = 25'b01010001_10001110_11011111_0;
      patterns[20881] = 25'b01010001_10001111_11100000_0;
      patterns[20882] = 25'b01010001_10010000_11100001_0;
      patterns[20883] = 25'b01010001_10010001_11100010_0;
      patterns[20884] = 25'b01010001_10010010_11100011_0;
      patterns[20885] = 25'b01010001_10010011_11100100_0;
      patterns[20886] = 25'b01010001_10010100_11100101_0;
      patterns[20887] = 25'b01010001_10010101_11100110_0;
      patterns[20888] = 25'b01010001_10010110_11100111_0;
      patterns[20889] = 25'b01010001_10010111_11101000_0;
      patterns[20890] = 25'b01010001_10011000_11101001_0;
      patterns[20891] = 25'b01010001_10011001_11101010_0;
      patterns[20892] = 25'b01010001_10011010_11101011_0;
      patterns[20893] = 25'b01010001_10011011_11101100_0;
      patterns[20894] = 25'b01010001_10011100_11101101_0;
      patterns[20895] = 25'b01010001_10011101_11101110_0;
      patterns[20896] = 25'b01010001_10011110_11101111_0;
      patterns[20897] = 25'b01010001_10011111_11110000_0;
      patterns[20898] = 25'b01010001_10100000_11110001_0;
      patterns[20899] = 25'b01010001_10100001_11110010_0;
      patterns[20900] = 25'b01010001_10100010_11110011_0;
      patterns[20901] = 25'b01010001_10100011_11110100_0;
      patterns[20902] = 25'b01010001_10100100_11110101_0;
      patterns[20903] = 25'b01010001_10100101_11110110_0;
      patterns[20904] = 25'b01010001_10100110_11110111_0;
      patterns[20905] = 25'b01010001_10100111_11111000_0;
      patterns[20906] = 25'b01010001_10101000_11111001_0;
      patterns[20907] = 25'b01010001_10101001_11111010_0;
      patterns[20908] = 25'b01010001_10101010_11111011_0;
      patterns[20909] = 25'b01010001_10101011_11111100_0;
      patterns[20910] = 25'b01010001_10101100_11111101_0;
      patterns[20911] = 25'b01010001_10101101_11111110_0;
      patterns[20912] = 25'b01010001_10101110_11111111_0;
      patterns[20913] = 25'b01010001_10101111_00000000_1;
      patterns[20914] = 25'b01010001_10110000_00000001_1;
      patterns[20915] = 25'b01010001_10110001_00000010_1;
      patterns[20916] = 25'b01010001_10110010_00000011_1;
      patterns[20917] = 25'b01010001_10110011_00000100_1;
      patterns[20918] = 25'b01010001_10110100_00000101_1;
      patterns[20919] = 25'b01010001_10110101_00000110_1;
      patterns[20920] = 25'b01010001_10110110_00000111_1;
      patterns[20921] = 25'b01010001_10110111_00001000_1;
      patterns[20922] = 25'b01010001_10111000_00001001_1;
      patterns[20923] = 25'b01010001_10111001_00001010_1;
      patterns[20924] = 25'b01010001_10111010_00001011_1;
      patterns[20925] = 25'b01010001_10111011_00001100_1;
      patterns[20926] = 25'b01010001_10111100_00001101_1;
      patterns[20927] = 25'b01010001_10111101_00001110_1;
      patterns[20928] = 25'b01010001_10111110_00001111_1;
      patterns[20929] = 25'b01010001_10111111_00010000_1;
      patterns[20930] = 25'b01010001_11000000_00010001_1;
      patterns[20931] = 25'b01010001_11000001_00010010_1;
      patterns[20932] = 25'b01010001_11000010_00010011_1;
      patterns[20933] = 25'b01010001_11000011_00010100_1;
      patterns[20934] = 25'b01010001_11000100_00010101_1;
      patterns[20935] = 25'b01010001_11000101_00010110_1;
      patterns[20936] = 25'b01010001_11000110_00010111_1;
      patterns[20937] = 25'b01010001_11000111_00011000_1;
      patterns[20938] = 25'b01010001_11001000_00011001_1;
      patterns[20939] = 25'b01010001_11001001_00011010_1;
      patterns[20940] = 25'b01010001_11001010_00011011_1;
      patterns[20941] = 25'b01010001_11001011_00011100_1;
      patterns[20942] = 25'b01010001_11001100_00011101_1;
      patterns[20943] = 25'b01010001_11001101_00011110_1;
      patterns[20944] = 25'b01010001_11001110_00011111_1;
      patterns[20945] = 25'b01010001_11001111_00100000_1;
      patterns[20946] = 25'b01010001_11010000_00100001_1;
      patterns[20947] = 25'b01010001_11010001_00100010_1;
      patterns[20948] = 25'b01010001_11010010_00100011_1;
      patterns[20949] = 25'b01010001_11010011_00100100_1;
      patterns[20950] = 25'b01010001_11010100_00100101_1;
      patterns[20951] = 25'b01010001_11010101_00100110_1;
      patterns[20952] = 25'b01010001_11010110_00100111_1;
      patterns[20953] = 25'b01010001_11010111_00101000_1;
      patterns[20954] = 25'b01010001_11011000_00101001_1;
      patterns[20955] = 25'b01010001_11011001_00101010_1;
      patterns[20956] = 25'b01010001_11011010_00101011_1;
      patterns[20957] = 25'b01010001_11011011_00101100_1;
      patterns[20958] = 25'b01010001_11011100_00101101_1;
      patterns[20959] = 25'b01010001_11011101_00101110_1;
      patterns[20960] = 25'b01010001_11011110_00101111_1;
      patterns[20961] = 25'b01010001_11011111_00110000_1;
      patterns[20962] = 25'b01010001_11100000_00110001_1;
      patterns[20963] = 25'b01010001_11100001_00110010_1;
      patterns[20964] = 25'b01010001_11100010_00110011_1;
      patterns[20965] = 25'b01010001_11100011_00110100_1;
      patterns[20966] = 25'b01010001_11100100_00110101_1;
      patterns[20967] = 25'b01010001_11100101_00110110_1;
      patterns[20968] = 25'b01010001_11100110_00110111_1;
      patterns[20969] = 25'b01010001_11100111_00111000_1;
      patterns[20970] = 25'b01010001_11101000_00111001_1;
      patterns[20971] = 25'b01010001_11101001_00111010_1;
      patterns[20972] = 25'b01010001_11101010_00111011_1;
      patterns[20973] = 25'b01010001_11101011_00111100_1;
      patterns[20974] = 25'b01010001_11101100_00111101_1;
      patterns[20975] = 25'b01010001_11101101_00111110_1;
      patterns[20976] = 25'b01010001_11101110_00111111_1;
      patterns[20977] = 25'b01010001_11101111_01000000_1;
      patterns[20978] = 25'b01010001_11110000_01000001_1;
      patterns[20979] = 25'b01010001_11110001_01000010_1;
      patterns[20980] = 25'b01010001_11110010_01000011_1;
      patterns[20981] = 25'b01010001_11110011_01000100_1;
      patterns[20982] = 25'b01010001_11110100_01000101_1;
      patterns[20983] = 25'b01010001_11110101_01000110_1;
      patterns[20984] = 25'b01010001_11110110_01000111_1;
      patterns[20985] = 25'b01010001_11110111_01001000_1;
      patterns[20986] = 25'b01010001_11111000_01001001_1;
      patterns[20987] = 25'b01010001_11111001_01001010_1;
      patterns[20988] = 25'b01010001_11111010_01001011_1;
      patterns[20989] = 25'b01010001_11111011_01001100_1;
      patterns[20990] = 25'b01010001_11111100_01001101_1;
      patterns[20991] = 25'b01010001_11111101_01001110_1;
      patterns[20992] = 25'b01010001_11111110_01001111_1;
      patterns[20993] = 25'b01010001_11111111_01010000_1;
      patterns[20994] = 25'b01010010_00000000_01010010_0;
      patterns[20995] = 25'b01010010_00000001_01010011_0;
      patterns[20996] = 25'b01010010_00000010_01010100_0;
      patterns[20997] = 25'b01010010_00000011_01010101_0;
      patterns[20998] = 25'b01010010_00000100_01010110_0;
      patterns[20999] = 25'b01010010_00000101_01010111_0;
      patterns[21000] = 25'b01010010_00000110_01011000_0;
      patterns[21001] = 25'b01010010_00000111_01011001_0;
      patterns[21002] = 25'b01010010_00001000_01011010_0;
      patterns[21003] = 25'b01010010_00001001_01011011_0;
      patterns[21004] = 25'b01010010_00001010_01011100_0;
      patterns[21005] = 25'b01010010_00001011_01011101_0;
      patterns[21006] = 25'b01010010_00001100_01011110_0;
      patterns[21007] = 25'b01010010_00001101_01011111_0;
      patterns[21008] = 25'b01010010_00001110_01100000_0;
      patterns[21009] = 25'b01010010_00001111_01100001_0;
      patterns[21010] = 25'b01010010_00010000_01100010_0;
      patterns[21011] = 25'b01010010_00010001_01100011_0;
      patterns[21012] = 25'b01010010_00010010_01100100_0;
      patterns[21013] = 25'b01010010_00010011_01100101_0;
      patterns[21014] = 25'b01010010_00010100_01100110_0;
      patterns[21015] = 25'b01010010_00010101_01100111_0;
      patterns[21016] = 25'b01010010_00010110_01101000_0;
      patterns[21017] = 25'b01010010_00010111_01101001_0;
      patterns[21018] = 25'b01010010_00011000_01101010_0;
      patterns[21019] = 25'b01010010_00011001_01101011_0;
      patterns[21020] = 25'b01010010_00011010_01101100_0;
      patterns[21021] = 25'b01010010_00011011_01101101_0;
      patterns[21022] = 25'b01010010_00011100_01101110_0;
      patterns[21023] = 25'b01010010_00011101_01101111_0;
      patterns[21024] = 25'b01010010_00011110_01110000_0;
      patterns[21025] = 25'b01010010_00011111_01110001_0;
      patterns[21026] = 25'b01010010_00100000_01110010_0;
      patterns[21027] = 25'b01010010_00100001_01110011_0;
      patterns[21028] = 25'b01010010_00100010_01110100_0;
      patterns[21029] = 25'b01010010_00100011_01110101_0;
      patterns[21030] = 25'b01010010_00100100_01110110_0;
      patterns[21031] = 25'b01010010_00100101_01110111_0;
      patterns[21032] = 25'b01010010_00100110_01111000_0;
      patterns[21033] = 25'b01010010_00100111_01111001_0;
      patterns[21034] = 25'b01010010_00101000_01111010_0;
      patterns[21035] = 25'b01010010_00101001_01111011_0;
      patterns[21036] = 25'b01010010_00101010_01111100_0;
      patterns[21037] = 25'b01010010_00101011_01111101_0;
      patterns[21038] = 25'b01010010_00101100_01111110_0;
      patterns[21039] = 25'b01010010_00101101_01111111_0;
      patterns[21040] = 25'b01010010_00101110_10000000_0;
      patterns[21041] = 25'b01010010_00101111_10000001_0;
      patterns[21042] = 25'b01010010_00110000_10000010_0;
      patterns[21043] = 25'b01010010_00110001_10000011_0;
      patterns[21044] = 25'b01010010_00110010_10000100_0;
      patterns[21045] = 25'b01010010_00110011_10000101_0;
      patterns[21046] = 25'b01010010_00110100_10000110_0;
      patterns[21047] = 25'b01010010_00110101_10000111_0;
      patterns[21048] = 25'b01010010_00110110_10001000_0;
      patterns[21049] = 25'b01010010_00110111_10001001_0;
      patterns[21050] = 25'b01010010_00111000_10001010_0;
      patterns[21051] = 25'b01010010_00111001_10001011_0;
      patterns[21052] = 25'b01010010_00111010_10001100_0;
      patterns[21053] = 25'b01010010_00111011_10001101_0;
      patterns[21054] = 25'b01010010_00111100_10001110_0;
      patterns[21055] = 25'b01010010_00111101_10001111_0;
      patterns[21056] = 25'b01010010_00111110_10010000_0;
      patterns[21057] = 25'b01010010_00111111_10010001_0;
      patterns[21058] = 25'b01010010_01000000_10010010_0;
      patterns[21059] = 25'b01010010_01000001_10010011_0;
      patterns[21060] = 25'b01010010_01000010_10010100_0;
      patterns[21061] = 25'b01010010_01000011_10010101_0;
      patterns[21062] = 25'b01010010_01000100_10010110_0;
      patterns[21063] = 25'b01010010_01000101_10010111_0;
      patterns[21064] = 25'b01010010_01000110_10011000_0;
      patterns[21065] = 25'b01010010_01000111_10011001_0;
      patterns[21066] = 25'b01010010_01001000_10011010_0;
      patterns[21067] = 25'b01010010_01001001_10011011_0;
      patterns[21068] = 25'b01010010_01001010_10011100_0;
      patterns[21069] = 25'b01010010_01001011_10011101_0;
      patterns[21070] = 25'b01010010_01001100_10011110_0;
      patterns[21071] = 25'b01010010_01001101_10011111_0;
      patterns[21072] = 25'b01010010_01001110_10100000_0;
      patterns[21073] = 25'b01010010_01001111_10100001_0;
      patterns[21074] = 25'b01010010_01010000_10100010_0;
      patterns[21075] = 25'b01010010_01010001_10100011_0;
      patterns[21076] = 25'b01010010_01010010_10100100_0;
      patterns[21077] = 25'b01010010_01010011_10100101_0;
      patterns[21078] = 25'b01010010_01010100_10100110_0;
      patterns[21079] = 25'b01010010_01010101_10100111_0;
      patterns[21080] = 25'b01010010_01010110_10101000_0;
      patterns[21081] = 25'b01010010_01010111_10101001_0;
      patterns[21082] = 25'b01010010_01011000_10101010_0;
      patterns[21083] = 25'b01010010_01011001_10101011_0;
      patterns[21084] = 25'b01010010_01011010_10101100_0;
      patterns[21085] = 25'b01010010_01011011_10101101_0;
      patterns[21086] = 25'b01010010_01011100_10101110_0;
      patterns[21087] = 25'b01010010_01011101_10101111_0;
      patterns[21088] = 25'b01010010_01011110_10110000_0;
      patterns[21089] = 25'b01010010_01011111_10110001_0;
      patterns[21090] = 25'b01010010_01100000_10110010_0;
      patterns[21091] = 25'b01010010_01100001_10110011_0;
      patterns[21092] = 25'b01010010_01100010_10110100_0;
      patterns[21093] = 25'b01010010_01100011_10110101_0;
      patterns[21094] = 25'b01010010_01100100_10110110_0;
      patterns[21095] = 25'b01010010_01100101_10110111_0;
      patterns[21096] = 25'b01010010_01100110_10111000_0;
      patterns[21097] = 25'b01010010_01100111_10111001_0;
      patterns[21098] = 25'b01010010_01101000_10111010_0;
      patterns[21099] = 25'b01010010_01101001_10111011_0;
      patterns[21100] = 25'b01010010_01101010_10111100_0;
      patterns[21101] = 25'b01010010_01101011_10111101_0;
      patterns[21102] = 25'b01010010_01101100_10111110_0;
      patterns[21103] = 25'b01010010_01101101_10111111_0;
      patterns[21104] = 25'b01010010_01101110_11000000_0;
      patterns[21105] = 25'b01010010_01101111_11000001_0;
      patterns[21106] = 25'b01010010_01110000_11000010_0;
      patterns[21107] = 25'b01010010_01110001_11000011_0;
      patterns[21108] = 25'b01010010_01110010_11000100_0;
      patterns[21109] = 25'b01010010_01110011_11000101_0;
      patterns[21110] = 25'b01010010_01110100_11000110_0;
      patterns[21111] = 25'b01010010_01110101_11000111_0;
      patterns[21112] = 25'b01010010_01110110_11001000_0;
      patterns[21113] = 25'b01010010_01110111_11001001_0;
      patterns[21114] = 25'b01010010_01111000_11001010_0;
      patterns[21115] = 25'b01010010_01111001_11001011_0;
      patterns[21116] = 25'b01010010_01111010_11001100_0;
      patterns[21117] = 25'b01010010_01111011_11001101_0;
      patterns[21118] = 25'b01010010_01111100_11001110_0;
      patterns[21119] = 25'b01010010_01111101_11001111_0;
      patterns[21120] = 25'b01010010_01111110_11010000_0;
      patterns[21121] = 25'b01010010_01111111_11010001_0;
      patterns[21122] = 25'b01010010_10000000_11010010_0;
      patterns[21123] = 25'b01010010_10000001_11010011_0;
      patterns[21124] = 25'b01010010_10000010_11010100_0;
      patterns[21125] = 25'b01010010_10000011_11010101_0;
      patterns[21126] = 25'b01010010_10000100_11010110_0;
      patterns[21127] = 25'b01010010_10000101_11010111_0;
      patterns[21128] = 25'b01010010_10000110_11011000_0;
      patterns[21129] = 25'b01010010_10000111_11011001_0;
      patterns[21130] = 25'b01010010_10001000_11011010_0;
      patterns[21131] = 25'b01010010_10001001_11011011_0;
      patterns[21132] = 25'b01010010_10001010_11011100_0;
      patterns[21133] = 25'b01010010_10001011_11011101_0;
      patterns[21134] = 25'b01010010_10001100_11011110_0;
      patterns[21135] = 25'b01010010_10001101_11011111_0;
      patterns[21136] = 25'b01010010_10001110_11100000_0;
      patterns[21137] = 25'b01010010_10001111_11100001_0;
      patterns[21138] = 25'b01010010_10010000_11100010_0;
      patterns[21139] = 25'b01010010_10010001_11100011_0;
      patterns[21140] = 25'b01010010_10010010_11100100_0;
      patterns[21141] = 25'b01010010_10010011_11100101_0;
      patterns[21142] = 25'b01010010_10010100_11100110_0;
      patterns[21143] = 25'b01010010_10010101_11100111_0;
      patterns[21144] = 25'b01010010_10010110_11101000_0;
      patterns[21145] = 25'b01010010_10010111_11101001_0;
      patterns[21146] = 25'b01010010_10011000_11101010_0;
      patterns[21147] = 25'b01010010_10011001_11101011_0;
      patterns[21148] = 25'b01010010_10011010_11101100_0;
      patterns[21149] = 25'b01010010_10011011_11101101_0;
      patterns[21150] = 25'b01010010_10011100_11101110_0;
      patterns[21151] = 25'b01010010_10011101_11101111_0;
      patterns[21152] = 25'b01010010_10011110_11110000_0;
      patterns[21153] = 25'b01010010_10011111_11110001_0;
      patterns[21154] = 25'b01010010_10100000_11110010_0;
      patterns[21155] = 25'b01010010_10100001_11110011_0;
      patterns[21156] = 25'b01010010_10100010_11110100_0;
      patterns[21157] = 25'b01010010_10100011_11110101_0;
      patterns[21158] = 25'b01010010_10100100_11110110_0;
      patterns[21159] = 25'b01010010_10100101_11110111_0;
      patterns[21160] = 25'b01010010_10100110_11111000_0;
      patterns[21161] = 25'b01010010_10100111_11111001_0;
      patterns[21162] = 25'b01010010_10101000_11111010_0;
      patterns[21163] = 25'b01010010_10101001_11111011_0;
      patterns[21164] = 25'b01010010_10101010_11111100_0;
      patterns[21165] = 25'b01010010_10101011_11111101_0;
      patterns[21166] = 25'b01010010_10101100_11111110_0;
      patterns[21167] = 25'b01010010_10101101_11111111_0;
      patterns[21168] = 25'b01010010_10101110_00000000_1;
      patterns[21169] = 25'b01010010_10101111_00000001_1;
      patterns[21170] = 25'b01010010_10110000_00000010_1;
      patterns[21171] = 25'b01010010_10110001_00000011_1;
      patterns[21172] = 25'b01010010_10110010_00000100_1;
      patterns[21173] = 25'b01010010_10110011_00000101_1;
      patterns[21174] = 25'b01010010_10110100_00000110_1;
      patterns[21175] = 25'b01010010_10110101_00000111_1;
      patterns[21176] = 25'b01010010_10110110_00001000_1;
      patterns[21177] = 25'b01010010_10110111_00001001_1;
      patterns[21178] = 25'b01010010_10111000_00001010_1;
      patterns[21179] = 25'b01010010_10111001_00001011_1;
      patterns[21180] = 25'b01010010_10111010_00001100_1;
      patterns[21181] = 25'b01010010_10111011_00001101_1;
      patterns[21182] = 25'b01010010_10111100_00001110_1;
      patterns[21183] = 25'b01010010_10111101_00001111_1;
      patterns[21184] = 25'b01010010_10111110_00010000_1;
      patterns[21185] = 25'b01010010_10111111_00010001_1;
      patterns[21186] = 25'b01010010_11000000_00010010_1;
      patterns[21187] = 25'b01010010_11000001_00010011_1;
      patterns[21188] = 25'b01010010_11000010_00010100_1;
      patterns[21189] = 25'b01010010_11000011_00010101_1;
      patterns[21190] = 25'b01010010_11000100_00010110_1;
      patterns[21191] = 25'b01010010_11000101_00010111_1;
      patterns[21192] = 25'b01010010_11000110_00011000_1;
      patterns[21193] = 25'b01010010_11000111_00011001_1;
      patterns[21194] = 25'b01010010_11001000_00011010_1;
      patterns[21195] = 25'b01010010_11001001_00011011_1;
      patterns[21196] = 25'b01010010_11001010_00011100_1;
      patterns[21197] = 25'b01010010_11001011_00011101_1;
      patterns[21198] = 25'b01010010_11001100_00011110_1;
      patterns[21199] = 25'b01010010_11001101_00011111_1;
      patterns[21200] = 25'b01010010_11001110_00100000_1;
      patterns[21201] = 25'b01010010_11001111_00100001_1;
      patterns[21202] = 25'b01010010_11010000_00100010_1;
      patterns[21203] = 25'b01010010_11010001_00100011_1;
      patterns[21204] = 25'b01010010_11010010_00100100_1;
      patterns[21205] = 25'b01010010_11010011_00100101_1;
      patterns[21206] = 25'b01010010_11010100_00100110_1;
      patterns[21207] = 25'b01010010_11010101_00100111_1;
      patterns[21208] = 25'b01010010_11010110_00101000_1;
      patterns[21209] = 25'b01010010_11010111_00101001_1;
      patterns[21210] = 25'b01010010_11011000_00101010_1;
      patterns[21211] = 25'b01010010_11011001_00101011_1;
      patterns[21212] = 25'b01010010_11011010_00101100_1;
      patterns[21213] = 25'b01010010_11011011_00101101_1;
      patterns[21214] = 25'b01010010_11011100_00101110_1;
      patterns[21215] = 25'b01010010_11011101_00101111_1;
      patterns[21216] = 25'b01010010_11011110_00110000_1;
      patterns[21217] = 25'b01010010_11011111_00110001_1;
      patterns[21218] = 25'b01010010_11100000_00110010_1;
      patterns[21219] = 25'b01010010_11100001_00110011_1;
      patterns[21220] = 25'b01010010_11100010_00110100_1;
      patterns[21221] = 25'b01010010_11100011_00110101_1;
      patterns[21222] = 25'b01010010_11100100_00110110_1;
      patterns[21223] = 25'b01010010_11100101_00110111_1;
      patterns[21224] = 25'b01010010_11100110_00111000_1;
      patterns[21225] = 25'b01010010_11100111_00111001_1;
      patterns[21226] = 25'b01010010_11101000_00111010_1;
      patterns[21227] = 25'b01010010_11101001_00111011_1;
      patterns[21228] = 25'b01010010_11101010_00111100_1;
      patterns[21229] = 25'b01010010_11101011_00111101_1;
      patterns[21230] = 25'b01010010_11101100_00111110_1;
      patterns[21231] = 25'b01010010_11101101_00111111_1;
      patterns[21232] = 25'b01010010_11101110_01000000_1;
      patterns[21233] = 25'b01010010_11101111_01000001_1;
      patterns[21234] = 25'b01010010_11110000_01000010_1;
      patterns[21235] = 25'b01010010_11110001_01000011_1;
      patterns[21236] = 25'b01010010_11110010_01000100_1;
      patterns[21237] = 25'b01010010_11110011_01000101_1;
      patterns[21238] = 25'b01010010_11110100_01000110_1;
      patterns[21239] = 25'b01010010_11110101_01000111_1;
      patterns[21240] = 25'b01010010_11110110_01001000_1;
      patterns[21241] = 25'b01010010_11110111_01001001_1;
      patterns[21242] = 25'b01010010_11111000_01001010_1;
      patterns[21243] = 25'b01010010_11111001_01001011_1;
      patterns[21244] = 25'b01010010_11111010_01001100_1;
      patterns[21245] = 25'b01010010_11111011_01001101_1;
      patterns[21246] = 25'b01010010_11111100_01001110_1;
      patterns[21247] = 25'b01010010_11111101_01001111_1;
      patterns[21248] = 25'b01010010_11111110_01010000_1;
      patterns[21249] = 25'b01010010_11111111_01010001_1;
      patterns[21250] = 25'b01010011_00000000_01010011_0;
      patterns[21251] = 25'b01010011_00000001_01010100_0;
      patterns[21252] = 25'b01010011_00000010_01010101_0;
      patterns[21253] = 25'b01010011_00000011_01010110_0;
      patterns[21254] = 25'b01010011_00000100_01010111_0;
      patterns[21255] = 25'b01010011_00000101_01011000_0;
      patterns[21256] = 25'b01010011_00000110_01011001_0;
      patterns[21257] = 25'b01010011_00000111_01011010_0;
      patterns[21258] = 25'b01010011_00001000_01011011_0;
      patterns[21259] = 25'b01010011_00001001_01011100_0;
      patterns[21260] = 25'b01010011_00001010_01011101_0;
      patterns[21261] = 25'b01010011_00001011_01011110_0;
      patterns[21262] = 25'b01010011_00001100_01011111_0;
      patterns[21263] = 25'b01010011_00001101_01100000_0;
      patterns[21264] = 25'b01010011_00001110_01100001_0;
      patterns[21265] = 25'b01010011_00001111_01100010_0;
      patterns[21266] = 25'b01010011_00010000_01100011_0;
      patterns[21267] = 25'b01010011_00010001_01100100_0;
      patterns[21268] = 25'b01010011_00010010_01100101_0;
      patterns[21269] = 25'b01010011_00010011_01100110_0;
      patterns[21270] = 25'b01010011_00010100_01100111_0;
      patterns[21271] = 25'b01010011_00010101_01101000_0;
      patterns[21272] = 25'b01010011_00010110_01101001_0;
      patterns[21273] = 25'b01010011_00010111_01101010_0;
      patterns[21274] = 25'b01010011_00011000_01101011_0;
      patterns[21275] = 25'b01010011_00011001_01101100_0;
      patterns[21276] = 25'b01010011_00011010_01101101_0;
      patterns[21277] = 25'b01010011_00011011_01101110_0;
      patterns[21278] = 25'b01010011_00011100_01101111_0;
      patterns[21279] = 25'b01010011_00011101_01110000_0;
      patterns[21280] = 25'b01010011_00011110_01110001_0;
      patterns[21281] = 25'b01010011_00011111_01110010_0;
      patterns[21282] = 25'b01010011_00100000_01110011_0;
      patterns[21283] = 25'b01010011_00100001_01110100_0;
      patterns[21284] = 25'b01010011_00100010_01110101_0;
      patterns[21285] = 25'b01010011_00100011_01110110_0;
      patterns[21286] = 25'b01010011_00100100_01110111_0;
      patterns[21287] = 25'b01010011_00100101_01111000_0;
      patterns[21288] = 25'b01010011_00100110_01111001_0;
      patterns[21289] = 25'b01010011_00100111_01111010_0;
      patterns[21290] = 25'b01010011_00101000_01111011_0;
      patterns[21291] = 25'b01010011_00101001_01111100_0;
      patterns[21292] = 25'b01010011_00101010_01111101_0;
      patterns[21293] = 25'b01010011_00101011_01111110_0;
      patterns[21294] = 25'b01010011_00101100_01111111_0;
      patterns[21295] = 25'b01010011_00101101_10000000_0;
      patterns[21296] = 25'b01010011_00101110_10000001_0;
      patterns[21297] = 25'b01010011_00101111_10000010_0;
      patterns[21298] = 25'b01010011_00110000_10000011_0;
      patterns[21299] = 25'b01010011_00110001_10000100_0;
      patterns[21300] = 25'b01010011_00110010_10000101_0;
      patterns[21301] = 25'b01010011_00110011_10000110_0;
      patterns[21302] = 25'b01010011_00110100_10000111_0;
      patterns[21303] = 25'b01010011_00110101_10001000_0;
      patterns[21304] = 25'b01010011_00110110_10001001_0;
      patterns[21305] = 25'b01010011_00110111_10001010_0;
      patterns[21306] = 25'b01010011_00111000_10001011_0;
      patterns[21307] = 25'b01010011_00111001_10001100_0;
      patterns[21308] = 25'b01010011_00111010_10001101_0;
      patterns[21309] = 25'b01010011_00111011_10001110_0;
      patterns[21310] = 25'b01010011_00111100_10001111_0;
      patterns[21311] = 25'b01010011_00111101_10010000_0;
      patterns[21312] = 25'b01010011_00111110_10010001_0;
      patterns[21313] = 25'b01010011_00111111_10010010_0;
      patterns[21314] = 25'b01010011_01000000_10010011_0;
      patterns[21315] = 25'b01010011_01000001_10010100_0;
      patterns[21316] = 25'b01010011_01000010_10010101_0;
      patterns[21317] = 25'b01010011_01000011_10010110_0;
      patterns[21318] = 25'b01010011_01000100_10010111_0;
      patterns[21319] = 25'b01010011_01000101_10011000_0;
      patterns[21320] = 25'b01010011_01000110_10011001_0;
      patterns[21321] = 25'b01010011_01000111_10011010_0;
      patterns[21322] = 25'b01010011_01001000_10011011_0;
      patterns[21323] = 25'b01010011_01001001_10011100_0;
      patterns[21324] = 25'b01010011_01001010_10011101_0;
      patterns[21325] = 25'b01010011_01001011_10011110_0;
      patterns[21326] = 25'b01010011_01001100_10011111_0;
      patterns[21327] = 25'b01010011_01001101_10100000_0;
      patterns[21328] = 25'b01010011_01001110_10100001_0;
      patterns[21329] = 25'b01010011_01001111_10100010_0;
      patterns[21330] = 25'b01010011_01010000_10100011_0;
      patterns[21331] = 25'b01010011_01010001_10100100_0;
      patterns[21332] = 25'b01010011_01010010_10100101_0;
      patterns[21333] = 25'b01010011_01010011_10100110_0;
      patterns[21334] = 25'b01010011_01010100_10100111_0;
      patterns[21335] = 25'b01010011_01010101_10101000_0;
      patterns[21336] = 25'b01010011_01010110_10101001_0;
      patterns[21337] = 25'b01010011_01010111_10101010_0;
      patterns[21338] = 25'b01010011_01011000_10101011_0;
      patterns[21339] = 25'b01010011_01011001_10101100_0;
      patterns[21340] = 25'b01010011_01011010_10101101_0;
      patterns[21341] = 25'b01010011_01011011_10101110_0;
      patterns[21342] = 25'b01010011_01011100_10101111_0;
      patterns[21343] = 25'b01010011_01011101_10110000_0;
      patterns[21344] = 25'b01010011_01011110_10110001_0;
      patterns[21345] = 25'b01010011_01011111_10110010_0;
      patterns[21346] = 25'b01010011_01100000_10110011_0;
      patterns[21347] = 25'b01010011_01100001_10110100_0;
      patterns[21348] = 25'b01010011_01100010_10110101_0;
      patterns[21349] = 25'b01010011_01100011_10110110_0;
      patterns[21350] = 25'b01010011_01100100_10110111_0;
      patterns[21351] = 25'b01010011_01100101_10111000_0;
      patterns[21352] = 25'b01010011_01100110_10111001_0;
      patterns[21353] = 25'b01010011_01100111_10111010_0;
      patterns[21354] = 25'b01010011_01101000_10111011_0;
      patterns[21355] = 25'b01010011_01101001_10111100_0;
      patterns[21356] = 25'b01010011_01101010_10111101_0;
      patterns[21357] = 25'b01010011_01101011_10111110_0;
      patterns[21358] = 25'b01010011_01101100_10111111_0;
      patterns[21359] = 25'b01010011_01101101_11000000_0;
      patterns[21360] = 25'b01010011_01101110_11000001_0;
      patterns[21361] = 25'b01010011_01101111_11000010_0;
      patterns[21362] = 25'b01010011_01110000_11000011_0;
      patterns[21363] = 25'b01010011_01110001_11000100_0;
      patterns[21364] = 25'b01010011_01110010_11000101_0;
      patterns[21365] = 25'b01010011_01110011_11000110_0;
      patterns[21366] = 25'b01010011_01110100_11000111_0;
      patterns[21367] = 25'b01010011_01110101_11001000_0;
      patterns[21368] = 25'b01010011_01110110_11001001_0;
      patterns[21369] = 25'b01010011_01110111_11001010_0;
      patterns[21370] = 25'b01010011_01111000_11001011_0;
      patterns[21371] = 25'b01010011_01111001_11001100_0;
      patterns[21372] = 25'b01010011_01111010_11001101_0;
      patterns[21373] = 25'b01010011_01111011_11001110_0;
      patterns[21374] = 25'b01010011_01111100_11001111_0;
      patterns[21375] = 25'b01010011_01111101_11010000_0;
      patterns[21376] = 25'b01010011_01111110_11010001_0;
      patterns[21377] = 25'b01010011_01111111_11010010_0;
      patterns[21378] = 25'b01010011_10000000_11010011_0;
      patterns[21379] = 25'b01010011_10000001_11010100_0;
      patterns[21380] = 25'b01010011_10000010_11010101_0;
      patterns[21381] = 25'b01010011_10000011_11010110_0;
      patterns[21382] = 25'b01010011_10000100_11010111_0;
      patterns[21383] = 25'b01010011_10000101_11011000_0;
      patterns[21384] = 25'b01010011_10000110_11011001_0;
      patterns[21385] = 25'b01010011_10000111_11011010_0;
      patterns[21386] = 25'b01010011_10001000_11011011_0;
      patterns[21387] = 25'b01010011_10001001_11011100_0;
      patterns[21388] = 25'b01010011_10001010_11011101_0;
      patterns[21389] = 25'b01010011_10001011_11011110_0;
      patterns[21390] = 25'b01010011_10001100_11011111_0;
      patterns[21391] = 25'b01010011_10001101_11100000_0;
      patterns[21392] = 25'b01010011_10001110_11100001_0;
      patterns[21393] = 25'b01010011_10001111_11100010_0;
      patterns[21394] = 25'b01010011_10010000_11100011_0;
      patterns[21395] = 25'b01010011_10010001_11100100_0;
      patterns[21396] = 25'b01010011_10010010_11100101_0;
      patterns[21397] = 25'b01010011_10010011_11100110_0;
      patterns[21398] = 25'b01010011_10010100_11100111_0;
      patterns[21399] = 25'b01010011_10010101_11101000_0;
      patterns[21400] = 25'b01010011_10010110_11101001_0;
      patterns[21401] = 25'b01010011_10010111_11101010_0;
      patterns[21402] = 25'b01010011_10011000_11101011_0;
      patterns[21403] = 25'b01010011_10011001_11101100_0;
      patterns[21404] = 25'b01010011_10011010_11101101_0;
      patterns[21405] = 25'b01010011_10011011_11101110_0;
      patterns[21406] = 25'b01010011_10011100_11101111_0;
      patterns[21407] = 25'b01010011_10011101_11110000_0;
      patterns[21408] = 25'b01010011_10011110_11110001_0;
      patterns[21409] = 25'b01010011_10011111_11110010_0;
      patterns[21410] = 25'b01010011_10100000_11110011_0;
      patterns[21411] = 25'b01010011_10100001_11110100_0;
      patterns[21412] = 25'b01010011_10100010_11110101_0;
      patterns[21413] = 25'b01010011_10100011_11110110_0;
      patterns[21414] = 25'b01010011_10100100_11110111_0;
      patterns[21415] = 25'b01010011_10100101_11111000_0;
      patterns[21416] = 25'b01010011_10100110_11111001_0;
      patterns[21417] = 25'b01010011_10100111_11111010_0;
      patterns[21418] = 25'b01010011_10101000_11111011_0;
      patterns[21419] = 25'b01010011_10101001_11111100_0;
      patterns[21420] = 25'b01010011_10101010_11111101_0;
      patterns[21421] = 25'b01010011_10101011_11111110_0;
      patterns[21422] = 25'b01010011_10101100_11111111_0;
      patterns[21423] = 25'b01010011_10101101_00000000_1;
      patterns[21424] = 25'b01010011_10101110_00000001_1;
      patterns[21425] = 25'b01010011_10101111_00000010_1;
      patterns[21426] = 25'b01010011_10110000_00000011_1;
      patterns[21427] = 25'b01010011_10110001_00000100_1;
      patterns[21428] = 25'b01010011_10110010_00000101_1;
      patterns[21429] = 25'b01010011_10110011_00000110_1;
      patterns[21430] = 25'b01010011_10110100_00000111_1;
      patterns[21431] = 25'b01010011_10110101_00001000_1;
      patterns[21432] = 25'b01010011_10110110_00001001_1;
      patterns[21433] = 25'b01010011_10110111_00001010_1;
      patterns[21434] = 25'b01010011_10111000_00001011_1;
      patterns[21435] = 25'b01010011_10111001_00001100_1;
      patterns[21436] = 25'b01010011_10111010_00001101_1;
      patterns[21437] = 25'b01010011_10111011_00001110_1;
      patterns[21438] = 25'b01010011_10111100_00001111_1;
      patterns[21439] = 25'b01010011_10111101_00010000_1;
      patterns[21440] = 25'b01010011_10111110_00010001_1;
      patterns[21441] = 25'b01010011_10111111_00010010_1;
      patterns[21442] = 25'b01010011_11000000_00010011_1;
      patterns[21443] = 25'b01010011_11000001_00010100_1;
      patterns[21444] = 25'b01010011_11000010_00010101_1;
      patterns[21445] = 25'b01010011_11000011_00010110_1;
      patterns[21446] = 25'b01010011_11000100_00010111_1;
      patterns[21447] = 25'b01010011_11000101_00011000_1;
      patterns[21448] = 25'b01010011_11000110_00011001_1;
      patterns[21449] = 25'b01010011_11000111_00011010_1;
      patterns[21450] = 25'b01010011_11001000_00011011_1;
      patterns[21451] = 25'b01010011_11001001_00011100_1;
      patterns[21452] = 25'b01010011_11001010_00011101_1;
      patterns[21453] = 25'b01010011_11001011_00011110_1;
      patterns[21454] = 25'b01010011_11001100_00011111_1;
      patterns[21455] = 25'b01010011_11001101_00100000_1;
      patterns[21456] = 25'b01010011_11001110_00100001_1;
      patterns[21457] = 25'b01010011_11001111_00100010_1;
      patterns[21458] = 25'b01010011_11010000_00100011_1;
      patterns[21459] = 25'b01010011_11010001_00100100_1;
      patterns[21460] = 25'b01010011_11010010_00100101_1;
      patterns[21461] = 25'b01010011_11010011_00100110_1;
      patterns[21462] = 25'b01010011_11010100_00100111_1;
      patterns[21463] = 25'b01010011_11010101_00101000_1;
      patterns[21464] = 25'b01010011_11010110_00101001_1;
      patterns[21465] = 25'b01010011_11010111_00101010_1;
      patterns[21466] = 25'b01010011_11011000_00101011_1;
      patterns[21467] = 25'b01010011_11011001_00101100_1;
      patterns[21468] = 25'b01010011_11011010_00101101_1;
      patterns[21469] = 25'b01010011_11011011_00101110_1;
      patterns[21470] = 25'b01010011_11011100_00101111_1;
      patterns[21471] = 25'b01010011_11011101_00110000_1;
      patterns[21472] = 25'b01010011_11011110_00110001_1;
      patterns[21473] = 25'b01010011_11011111_00110010_1;
      patterns[21474] = 25'b01010011_11100000_00110011_1;
      patterns[21475] = 25'b01010011_11100001_00110100_1;
      patterns[21476] = 25'b01010011_11100010_00110101_1;
      patterns[21477] = 25'b01010011_11100011_00110110_1;
      patterns[21478] = 25'b01010011_11100100_00110111_1;
      patterns[21479] = 25'b01010011_11100101_00111000_1;
      patterns[21480] = 25'b01010011_11100110_00111001_1;
      patterns[21481] = 25'b01010011_11100111_00111010_1;
      patterns[21482] = 25'b01010011_11101000_00111011_1;
      patterns[21483] = 25'b01010011_11101001_00111100_1;
      patterns[21484] = 25'b01010011_11101010_00111101_1;
      patterns[21485] = 25'b01010011_11101011_00111110_1;
      patterns[21486] = 25'b01010011_11101100_00111111_1;
      patterns[21487] = 25'b01010011_11101101_01000000_1;
      patterns[21488] = 25'b01010011_11101110_01000001_1;
      patterns[21489] = 25'b01010011_11101111_01000010_1;
      patterns[21490] = 25'b01010011_11110000_01000011_1;
      patterns[21491] = 25'b01010011_11110001_01000100_1;
      patterns[21492] = 25'b01010011_11110010_01000101_1;
      patterns[21493] = 25'b01010011_11110011_01000110_1;
      patterns[21494] = 25'b01010011_11110100_01000111_1;
      patterns[21495] = 25'b01010011_11110101_01001000_1;
      patterns[21496] = 25'b01010011_11110110_01001001_1;
      patterns[21497] = 25'b01010011_11110111_01001010_1;
      patterns[21498] = 25'b01010011_11111000_01001011_1;
      patterns[21499] = 25'b01010011_11111001_01001100_1;
      patterns[21500] = 25'b01010011_11111010_01001101_1;
      patterns[21501] = 25'b01010011_11111011_01001110_1;
      patterns[21502] = 25'b01010011_11111100_01001111_1;
      patterns[21503] = 25'b01010011_11111101_01010000_1;
      patterns[21504] = 25'b01010011_11111110_01010001_1;
      patterns[21505] = 25'b01010011_11111111_01010010_1;
      patterns[21506] = 25'b01010100_00000000_01010100_0;
      patterns[21507] = 25'b01010100_00000001_01010101_0;
      patterns[21508] = 25'b01010100_00000010_01010110_0;
      patterns[21509] = 25'b01010100_00000011_01010111_0;
      patterns[21510] = 25'b01010100_00000100_01011000_0;
      patterns[21511] = 25'b01010100_00000101_01011001_0;
      patterns[21512] = 25'b01010100_00000110_01011010_0;
      patterns[21513] = 25'b01010100_00000111_01011011_0;
      patterns[21514] = 25'b01010100_00001000_01011100_0;
      patterns[21515] = 25'b01010100_00001001_01011101_0;
      patterns[21516] = 25'b01010100_00001010_01011110_0;
      patterns[21517] = 25'b01010100_00001011_01011111_0;
      patterns[21518] = 25'b01010100_00001100_01100000_0;
      patterns[21519] = 25'b01010100_00001101_01100001_0;
      patterns[21520] = 25'b01010100_00001110_01100010_0;
      patterns[21521] = 25'b01010100_00001111_01100011_0;
      patterns[21522] = 25'b01010100_00010000_01100100_0;
      patterns[21523] = 25'b01010100_00010001_01100101_0;
      patterns[21524] = 25'b01010100_00010010_01100110_0;
      patterns[21525] = 25'b01010100_00010011_01100111_0;
      patterns[21526] = 25'b01010100_00010100_01101000_0;
      patterns[21527] = 25'b01010100_00010101_01101001_0;
      patterns[21528] = 25'b01010100_00010110_01101010_0;
      patterns[21529] = 25'b01010100_00010111_01101011_0;
      patterns[21530] = 25'b01010100_00011000_01101100_0;
      patterns[21531] = 25'b01010100_00011001_01101101_0;
      patterns[21532] = 25'b01010100_00011010_01101110_0;
      patterns[21533] = 25'b01010100_00011011_01101111_0;
      patterns[21534] = 25'b01010100_00011100_01110000_0;
      patterns[21535] = 25'b01010100_00011101_01110001_0;
      patterns[21536] = 25'b01010100_00011110_01110010_0;
      patterns[21537] = 25'b01010100_00011111_01110011_0;
      patterns[21538] = 25'b01010100_00100000_01110100_0;
      patterns[21539] = 25'b01010100_00100001_01110101_0;
      patterns[21540] = 25'b01010100_00100010_01110110_0;
      patterns[21541] = 25'b01010100_00100011_01110111_0;
      patterns[21542] = 25'b01010100_00100100_01111000_0;
      patterns[21543] = 25'b01010100_00100101_01111001_0;
      patterns[21544] = 25'b01010100_00100110_01111010_0;
      patterns[21545] = 25'b01010100_00100111_01111011_0;
      patterns[21546] = 25'b01010100_00101000_01111100_0;
      patterns[21547] = 25'b01010100_00101001_01111101_0;
      patterns[21548] = 25'b01010100_00101010_01111110_0;
      patterns[21549] = 25'b01010100_00101011_01111111_0;
      patterns[21550] = 25'b01010100_00101100_10000000_0;
      patterns[21551] = 25'b01010100_00101101_10000001_0;
      patterns[21552] = 25'b01010100_00101110_10000010_0;
      patterns[21553] = 25'b01010100_00101111_10000011_0;
      patterns[21554] = 25'b01010100_00110000_10000100_0;
      patterns[21555] = 25'b01010100_00110001_10000101_0;
      patterns[21556] = 25'b01010100_00110010_10000110_0;
      patterns[21557] = 25'b01010100_00110011_10000111_0;
      patterns[21558] = 25'b01010100_00110100_10001000_0;
      patterns[21559] = 25'b01010100_00110101_10001001_0;
      patterns[21560] = 25'b01010100_00110110_10001010_0;
      patterns[21561] = 25'b01010100_00110111_10001011_0;
      patterns[21562] = 25'b01010100_00111000_10001100_0;
      patterns[21563] = 25'b01010100_00111001_10001101_0;
      patterns[21564] = 25'b01010100_00111010_10001110_0;
      patterns[21565] = 25'b01010100_00111011_10001111_0;
      patterns[21566] = 25'b01010100_00111100_10010000_0;
      patterns[21567] = 25'b01010100_00111101_10010001_0;
      patterns[21568] = 25'b01010100_00111110_10010010_0;
      patterns[21569] = 25'b01010100_00111111_10010011_0;
      patterns[21570] = 25'b01010100_01000000_10010100_0;
      patterns[21571] = 25'b01010100_01000001_10010101_0;
      patterns[21572] = 25'b01010100_01000010_10010110_0;
      patterns[21573] = 25'b01010100_01000011_10010111_0;
      patterns[21574] = 25'b01010100_01000100_10011000_0;
      patterns[21575] = 25'b01010100_01000101_10011001_0;
      patterns[21576] = 25'b01010100_01000110_10011010_0;
      patterns[21577] = 25'b01010100_01000111_10011011_0;
      patterns[21578] = 25'b01010100_01001000_10011100_0;
      patterns[21579] = 25'b01010100_01001001_10011101_0;
      patterns[21580] = 25'b01010100_01001010_10011110_0;
      patterns[21581] = 25'b01010100_01001011_10011111_0;
      patterns[21582] = 25'b01010100_01001100_10100000_0;
      patterns[21583] = 25'b01010100_01001101_10100001_0;
      patterns[21584] = 25'b01010100_01001110_10100010_0;
      patterns[21585] = 25'b01010100_01001111_10100011_0;
      patterns[21586] = 25'b01010100_01010000_10100100_0;
      patterns[21587] = 25'b01010100_01010001_10100101_0;
      patterns[21588] = 25'b01010100_01010010_10100110_0;
      patterns[21589] = 25'b01010100_01010011_10100111_0;
      patterns[21590] = 25'b01010100_01010100_10101000_0;
      patterns[21591] = 25'b01010100_01010101_10101001_0;
      patterns[21592] = 25'b01010100_01010110_10101010_0;
      patterns[21593] = 25'b01010100_01010111_10101011_0;
      patterns[21594] = 25'b01010100_01011000_10101100_0;
      patterns[21595] = 25'b01010100_01011001_10101101_0;
      patterns[21596] = 25'b01010100_01011010_10101110_0;
      patterns[21597] = 25'b01010100_01011011_10101111_0;
      patterns[21598] = 25'b01010100_01011100_10110000_0;
      patterns[21599] = 25'b01010100_01011101_10110001_0;
      patterns[21600] = 25'b01010100_01011110_10110010_0;
      patterns[21601] = 25'b01010100_01011111_10110011_0;
      patterns[21602] = 25'b01010100_01100000_10110100_0;
      patterns[21603] = 25'b01010100_01100001_10110101_0;
      patterns[21604] = 25'b01010100_01100010_10110110_0;
      patterns[21605] = 25'b01010100_01100011_10110111_0;
      patterns[21606] = 25'b01010100_01100100_10111000_0;
      patterns[21607] = 25'b01010100_01100101_10111001_0;
      patterns[21608] = 25'b01010100_01100110_10111010_0;
      patterns[21609] = 25'b01010100_01100111_10111011_0;
      patterns[21610] = 25'b01010100_01101000_10111100_0;
      patterns[21611] = 25'b01010100_01101001_10111101_0;
      patterns[21612] = 25'b01010100_01101010_10111110_0;
      patterns[21613] = 25'b01010100_01101011_10111111_0;
      patterns[21614] = 25'b01010100_01101100_11000000_0;
      patterns[21615] = 25'b01010100_01101101_11000001_0;
      patterns[21616] = 25'b01010100_01101110_11000010_0;
      patterns[21617] = 25'b01010100_01101111_11000011_0;
      patterns[21618] = 25'b01010100_01110000_11000100_0;
      patterns[21619] = 25'b01010100_01110001_11000101_0;
      patterns[21620] = 25'b01010100_01110010_11000110_0;
      patterns[21621] = 25'b01010100_01110011_11000111_0;
      patterns[21622] = 25'b01010100_01110100_11001000_0;
      patterns[21623] = 25'b01010100_01110101_11001001_0;
      patterns[21624] = 25'b01010100_01110110_11001010_0;
      patterns[21625] = 25'b01010100_01110111_11001011_0;
      patterns[21626] = 25'b01010100_01111000_11001100_0;
      patterns[21627] = 25'b01010100_01111001_11001101_0;
      patterns[21628] = 25'b01010100_01111010_11001110_0;
      patterns[21629] = 25'b01010100_01111011_11001111_0;
      patterns[21630] = 25'b01010100_01111100_11010000_0;
      patterns[21631] = 25'b01010100_01111101_11010001_0;
      patterns[21632] = 25'b01010100_01111110_11010010_0;
      patterns[21633] = 25'b01010100_01111111_11010011_0;
      patterns[21634] = 25'b01010100_10000000_11010100_0;
      patterns[21635] = 25'b01010100_10000001_11010101_0;
      patterns[21636] = 25'b01010100_10000010_11010110_0;
      patterns[21637] = 25'b01010100_10000011_11010111_0;
      patterns[21638] = 25'b01010100_10000100_11011000_0;
      patterns[21639] = 25'b01010100_10000101_11011001_0;
      patterns[21640] = 25'b01010100_10000110_11011010_0;
      patterns[21641] = 25'b01010100_10000111_11011011_0;
      patterns[21642] = 25'b01010100_10001000_11011100_0;
      patterns[21643] = 25'b01010100_10001001_11011101_0;
      patterns[21644] = 25'b01010100_10001010_11011110_0;
      patterns[21645] = 25'b01010100_10001011_11011111_0;
      patterns[21646] = 25'b01010100_10001100_11100000_0;
      patterns[21647] = 25'b01010100_10001101_11100001_0;
      patterns[21648] = 25'b01010100_10001110_11100010_0;
      patterns[21649] = 25'b01010100_10001111_11100011_0;
      patterns[21650] = 25'b01010100_10010000_11100100_0;
      patterns[21651] = 25'b01010100_10010001_11100101_0;
      patterns[21652] = 25'b01010100_10010010_11100110_0;
      patterns[21653] = 25'b01010100_10010011_11100111_0;
      patterns[21654] = 25'b01010100_10010100_11101000_0;
      patterns[21655] = 25'b01010100_10010101_11101001_0;
      patterns[21656] = 25'b01010100_10010110_11101010_0;
      patterns[21657] = 25'b01010100_10010111_11101011_0;
      patterns[21658] = 25'b01010100_10011000_11101100_0;
      patterns[21659] = 25'b01010100_10011001_11101101_0;
      patterns[21660] = 25'b01010100_10011010_11101110_0;
      patterns[21661] = 25'b01010100_10011011_11101111_0;
      patterns[21662] = 25'b01010100_10011100_11110000_0;
      patterns[21663] = 25'b01010100_10011101_11110001_0;
      patterns[21664] = 25'b01010100_10011110_11110010_0;
      patterns[21665] = 25'b01010100_10011111_11110011_0;
      patterns[21666] = 25'b01010100_10100000_11110100_0;
      patterns[21667] = 25'b01010100_10100001_11110101_0;
      patterns[21668] = 25'b01010100_10100010_11110110_0;
      patterns[21669] = 25'b01010100_10100011_11110111_0;
      patterns[21670] = 25'b01010100_10100100_11111000_0;
      patterns[21671] = 25'b01010100_10100101_11111001_0;
      patterns[21672] = 25'b01010100_10100110_11111010_0;
      patterns[21673] = 25'b01010100_10100111_11111011_0;
      patterns[21674] = 25'b01010100_10101000_11111100_0;
      patterns[21675] = 25'b01010100_10101001_11111101_0;
      patterns[21676] = 25'b01010100_10101010_11111110_0;
      patterns[21677] = 25'b01010100_10101011_11111111_0;
      patterns[21678] = 25'b01010100_10101100_00000000_1;
      patterns[21679] = 25'b01010100_10101101_00000001_1;
      patterns[21680] = 25'b01010100_10101110_00000010_1;
      patterns[21681] = 25'b01010100_10101111_00000011_1;
      patterns[21682] = 25'b01010100_10110000_00000100_1;
      patterns[21683] = 25'b01010100_10110001_00000101_1;
      patterns[21684] = 25'b01010100_10110010_00000110_1;
      patterns[21685] = 25'b01010100_10110011_00000111_1;
      patterns[21686] = 25'b01010100_10110100_00001000_1;
      patterns[21687] = 25'b01010100_10110101_00001001_1;
      patterns[21688] = 25'b01010100_10110110_00001010_1;
      patterns[21689] = 25'b01010100_10110111_00001011_1;
      patterns[21690] = 25'b01010100_10111000_00001100_1;
      patterns[21691] = 25'b01010100_10111001_00001101_1;
      patterns[21692] = 25'b01010100_10111010_00001110_1;
      patterns[21693] = 25'b01010100_10111011_00001111_1;
      patterns[21694] = 25'b01010100_10111100_00010000_1;
      patterns[21695] = 25'b01010100_10111101_00010001_1;
      patterns[21696] = 25'b01010100_10111110_00010010_1;
      patterns[21697] = 25'b01010100_10111111_00010011_1;
      patterns[21698] = 25'b01010100_11000000_00010100_1;
      patterns[21699] = 25'b01010100_11000001_00010101_1;
      patterns[21700] = 25'b01010100_11000010_00010110_1;
      patterns[21701] = 25'b01010100_11000011_00010111_1;
      patterns[21702] = 25'b01010100_11000100_00011000_1;
      patterns[21703] = 25'b01010100_11000101_00011001_1;
      patterns[21704] = 25'b01010100_11000110_00011010_1;
      patterns[21705] = 25'b01010100_11000111_00011011_1;
      patterns[21706] = 25'b01010100_11001000_00011100_1;
      patterns[21707] = 25'b01010100_11001001_00011101_1;
      patterns[21708] = 25'b01010100_11001010_00011110_1;
      patterns[21709] = 25'b01010100_11001011_00011111_1;
      patterns[21710] = 25'b01010100_11001100_00100000_1;
      patterns[21711] = 25'b01010100_11001101_00100001_1;
      patterns[21712] = 25'b01010100_11001110_00100010_1;
      patterns[21713] = 25'b01010100_11001111_00100011_1;
      patterns[21714] = 25'b01010100_11010000_00100100_1;
      patterns[21715] = 25'b01010100_11010001_00100101_1;
      patterns[21716] = 25'b01010100_11010010_00100110_1;
      patterns[21717] = 25'b01010100_11010011_00100111_1;
      patterns[21718] = 25'b01010100_11010100_00101000_1;
      patterns[21719] = 25'b01010100_11010101_00101001_1;
      patterns[21720] = 25'b01010100_11010110_00101010_1;
      patterns[21721] = 25'b01010100_11010111_00101011_1;
      patterns[21722] = 25'b01010100_11011000_00101100_1;
      patterns[21723] = 25'b01010100_11011001_00101101_1;
      patterns[21724] = 25'b01010100_11011010_00101110_1;
      patterns[21725] = 25'b01010100_11011011_00101111_1;
      patterns[21726] = 25'b01010100_11011100_00110000_1;
      patterns[21727] = 25'b01010100_11011101_00110001_1;
      patterns[21728] = 25'b01010100_11011110_00110010_1;
      patterns[21729] = 25'b01010100_11011111_00110011_1;
      patterns[21730] = 25'b01010100_11100000_00110100_1;
      patterns[21731] = 25'b01010100_11100001_00110101_1;
      patterns[21732] = 25'b01010100_11100010_00110110_1;
      patterns[21733] = 25'b01010100_11100011_00110111_1;
      patterns[21734] = 25'b01010100_11100100_00111000_1;
      patterns[21735] = 25'b01010100_11100101_00111001_1;
      patterns[21736] = 25'b01010100_11100110_00111010_1;
      patterns[21737] = 25'b01010100_11100111_00111011_1;
      patterns[21738] = 25'b01010100_11101000_00111100_1;
      patterns[21739] = 25'b01010100_11101001_00111101_1;
      patterns[21740] = 25'b01010100_11101010_00111110_1;
      patterns[21741] = 25'b01010100_11101011_00111111_1;
      patterns[21742] = 25'b01010100_11101100_01000000_1;
      patterns[21743] = 25'b01010100_11101101_01000001_1;
      patterns[21744] = 25'b01010100_11101110_01000010_1;
      patterns[21745] = 25'b01010100_11101111_01000011_1;
      patterns[21746] = 25'b01010100_11110000_01000100_1;
      patterns[21747] = 25'b01010100_11110001_01000101_1;
      patterns[21748] = 25'b01010100_11110010_01000110_1;
      patterns[21749] = 25'b01010100_11110011_01000111_1;
      patterns[21750] = 25'b01010100_11110100_01001000_1;
      patterns[21751] = 25'b01010100_11110101_01001001_1;
      patterns[21752] = 25'b01010100_11110110_01001010_1;
      patterns[21753] = 25'b01010100_11110111_01001011_1;
      patterns[21754] = 25'b01010100_11111000_01001100_1;
      patterns[21755] = 25'b01010100_11111001_01001101_1;
      patterns[21756] = 25'b01010100_11111010_01001110_1;
      patterns[21757] = 25'b01010100_11111011_01001111_1;
      patterns[21758] = 25'b01010100_11111100_01010000_1;
      patterns[21759] = 25'b01010100_11111101_01010001_1;
      patterns[21760] = 25'b01010100_11111110_01010010_1;
      patterns[21761] = 25'b01010100_11111111_01010011_1;
      patterns[21762] = 25'b01010101_00000000_01010101_0;
      patterns[21763] = 25'b01010101_00000001_01010110_0;
      patterns[21764] = 25'b01010101_00000010_01010111_0;
      patterns[21765] = 25'b01010101_00000011_01011000_0;
      patterns[21766] = 25'b01010101_00000100_01011001_0;
      patterns[21767] = 25'b01010101_00000101_01011010_0;
      patterns[21768] = 25'b01010101_00000110_01011011_0;
      patterns[21769] = 25'b01010101_00000111_01011100_0;
      patterns[21770] = 25'b01010101_00001000_01011101_0;
      patterns[21771] = 25'b01010101_00001001_01011110_0;
      patterns[21772] = 25'b01010101_00001010_01011111_0;
      patterns[21773] = 25'b01010101_00001011_01100000_0;
      patterns[21774] = 25'b01010101_00001100_01100001_0;
      patterns[21775] = 25'b01010101_00001101_01100010_0;
      patterns[21776] = 25'b01010101_00001110_01100011_0;
      patterns[21777] = 25'b01010101_00001111_01100100_0;
      patterns[21778] = 25'b01010101_00010000_01100101_0;
      patterns[21779] = 25'b01010101_00010001_01100110_0;
      patterns[21780] = 25'b01010101_00010010_01100111_0;
      patterns[21781] = 25'b01010101_00010011_01101000_0;
      patterns[21782] = 25'b01010101_00010100_01101001_0;
      patterns[21783] = 25'b01010101_00010101_01101010_0;
      patterns[21784] = 25'b01010101_00010110_01101011_0;
      patterns[21785] = 25'b01010101_00010111_01101100_0;
      patterns[21786] = 25'b01010101_00011000_01101101_0;
      patterns[21787] = 25'b01010101_00011001_01101110_0;
      patterns[21788] = 25'b01010101_00011010_01101111_0;
      patterns[21789] = 25'b01010101_00011011_01110000_0;
      patterns[21790] = 25'b01010101_00011100_01110001_0;
      patterns[21791] = 25'b01010101_00011101_01110010_0;
      patterns[21792] = 25'b01010101_00011110_01110011_0;
      patterns[21793] = 25'b01010101_00011111_01110100_0;
      patterns[21794] = 25'b01010101_00100000_01110101_0;
      patterns[21795] = 25'b01010101_00100001_01110110_0;
      patterns[21796] = 25'b01010101_00100010_01110111_0;
      patterns[21797] = 25'b01010101_00100011_01111000_0;
      patterns[21798] = 25'b01010101_00100100_01111001_0;
      patterns[21799] = 25'b01010101_00100101_01111010_0;
      patterns[21800] = 25'b01010101_00100110_01111011_0;
      patterns[21801] = 25'b01010101_00100111_01111100_0;
      patterns[21802] = 25'b01010101_00101000_01111101_0;
      patterns[21803] = 25'b01010101_00101001_01111110_0;
      patterns[21804] = 25'b01010101_00101010_01111111_0;
      patterns[21805] = 25'b01010101_00101011_10000000_0;
      patterns[21806] = 25'b01010101_00101100_10000001_0;
      patterns[21807] = 25'b01010101_00101101_10000010_0;
      patterns[21808] = 25'b01010101_00101110_10000011_0;
      patterns[21809] = 25'b01010101_00101111_10000100_0;
      patterns[21810] = 25'b01010101_00110000_10000101_0;
      patterns[21811] = 25'b01010101_00110001_10000110_0;
      patterns[21812] = 25'b01010101_00110010_10000111_0;
      patterns[21813] = 25'b01010101_00110011_10001000_0;
      patterns[21814] = 25'b01010101_00110100_10001001_0;
      patterns[21815] = 25'b01010101_00110101_10001010_0;
      patterns[21816] = 25'b01010101_00110110_10001011_0;
      patterns[21817] = 25'b01010101_00110111_10001100_0;
      patterns[21818] = 25'b01010101_00111000_10001101_0;
      patterns[21819] = 25'b01010101_00111001_10001110_0;
      patterns[21820] = 25'b01010101_00111010_10001111_0;
      patterns[21821] = 25'b01010101_00111011_10010000_0;
      patterns[21822] = 25'b01010101_00111100_10010001_0;
      patterns[21823] = 25'b01010101_00111101_10010010_0;
      patterns[21824] = 25'b01010101_00111110_10010011_0;
      patterns[21825] = 25'b01010101_00111111_10010100_0;
      patterns[21826] = 25'b01010101_01000000_10010101_0;
      patterns[21827] = 25'b01010101_01000001_10010110_0;
      patterns[21828] = 25'b01010101_01000010_10010111_0;
      patterns[21829] = 25'b01010101_01000011_10011000_0;
      patterns[21830] = 25'b01010101_01000100_10011001_0;
      patterns[21831] = 25'b01010101_01000101_10011010_0;
      patterns[21832] = 25'b01010101_01000110_10011011_0;
      patterns[21833] = 25'b01010101_01000111_10011100_0;
      patterns[21834] = 25'b01010101_01001000_10011101_0;
      patterns[21835] = 25'b01010101_01001001_10011110_0;
      patterns[21836] = 25'b01010101_01001010_10011111_0;
      patterns[21837] = 25'b01010101_01001011_10100000_0;
      patterns[21838] = 25'b01010101_01001100_10100001_0;
      patterns[21839] = 25'b01010101_01001101_10100010_0;
      patterns[21840] = 25'b01010101_01001110_10100011_0;
      patterns[21841] = 25'b01010101_01001111_10100100_0;
      patterns[21842] = 25'b01010101_01010000_10100101_0;
      patterns[21843] = 25'b01010101_01010001_10100110_0;
      patterns[21844] = 25'b01010101_01010010_10100111_0;
      patterns[21845] = 25'b01010101_01010011_10101000_0;
      patterns[21846] = 25'b01010101_01010100_10101001_0;
      patterns[21847] = 25'b01010101_01010101_10101010_0;
      patterns[21848] = 25'b01010101_01010110_10101011_0;
      patterns[21849] = 25'b01010101_01010111_10101100_0;
      patterns[21850] = 25'b01010101_01011000_10101101_0;
      patterns[21851] = 25'b01010101_01011001_10101110_0;
      patterns[21852] = 25'b01010101_01011010_10101111_0;
      patterns[21853] = 25'b01010101_01011011_10110000_0;
      patterns[21854] = 25'b01010101_01011100_10110001_0;
      patterns[21855] = 25'b01010101_01011101_10110010_0;
      patterns[21856] = 25'b01010101_01011110_10110011_0;
      patterns[21857] = 25'b01010101_01011111_10110100_0;
      patterns[21858] = 25'b01010101_01100000_10110101_0;
      patterns[21859] = 25'b01010101_01100001_10110110_0;
      patterns[21860] = 25'b01010101_01100010_10110111_0;
      patterns[21861] = 25'b01010101_01100011_10111000_0;
      patterns[21862] = 25'b01010101_01100100_10111001_0;
      patterns[21863] = 25'b01010101_01100101_10111010_0;
      patterns[21864] = 25'b01010101_01100110_10111011_0;
      patterns[21865] = 25'b01010101_01100111_10111100_0;
      patterns[21866] = 25'b01010101_01101000_10111101_0;
      patterns[21867] = 25'b01010101_01101001_10111110_0;
      patterns[21868] = 25'b01010101_01101010_10111111_0;
      patterns[21869] = 25'b01010101_01101011_11000000_0;
      patterns[21870] = 25'b01010101_01101100_11000001_0;
      patterns[21871] = 25'b01010101_01101101_11000010_0;
      patterns[21872] = 25'b01010101_01101110_11000011_0;
      patterns[21873] = 25'b01010101_01101111_11000100_0;
      patterns[21874] = 25'b01010101_01110000_11000101_0;
      patterns[21875] = 25'b01010101_01110001_11000110_0;
      patterns[21876] = 25'b01010101_01110010_11000111_0;
      patterns[21877] = 25'b01010101_01110011_11001000_0;
      patterns[21878] = 25'b01010101_01110100_11001001_0;
      patterns[21879] = 25'b01010101_01110101_11001010_0;
      patterns[21880] = 25'b01010101_01110110_11001011_0;
      patterns[21881] = 25'b01010101_01110111_11001100_0;
      patterns[21882] = 25'b01010101_01111000_11001101_0;
      patterns[21883] = 25'b01010101_01111001_11001110_0;
      patterns[21884] = 25'b01010101_01111010_11001111_0;
      patterns[21885] = 25'b01010101_01111011_11010000_0;
      patterns[21886] = 25'b01010101_01111100_11010001_0;
      patterns[21887] = 25'b01010101_01111101_11010010_0;
      patterns[21888] = 25'b01010101_01111110_11010011_0;
      patterns[21889] = 25'b01010101_01111111_11010100_0;
      patterns[21890] = 25'b01010101_10000000_11010101_0;
      patterns[21891] = 25'b01010101_10000001_11010110_0;
      patterns[21892] = 25'b01010101_10000010_11010111_0;
      patterns[21893] = 25'b01010101_10000011_11011000_0;
      patterns[21894] = 25'b01010101_10000100_11011001_0;
      patterns[21895] = 25'b01010101_10000101_11011010_0;
      patterns[21896] = 25'b01010101_10000110_11011011_0;
      patterns[21897] = 25'b01010101_10000111_11011100_0;
      patterns[21898] = 25'b01010101_10001000_11011101_0;
      patterns[21899] = 25'b01010101_10001001_11011110_0;
      patterns[21900] = 25'b01010101_10001010_11011111_0;
      patterns[21901] = 25'b01010101_10001011_11100000_0;
      patterns[21902] = 25'b01010101_10001100_11100001_0;
      patterns[21903] = 25'b01010101_10001101_11100010_0;
      patterns[21904] = 25'b01010101_10001110_11100011_0;
      patterns[21905] = 25'b01010101_10001111_11100100_0;
      patterns[21906] = 25'b01010101_10010000_11100101_0;
      patterns[21907] = 25'b01010101_10010001_11100110_0;
      patterns[21908] = 25'b01010101_10010010_11100111_0;
      patterns[21909] = 25'b01010101_10010011_11101000_0;
      patterns[21910] = 25'b01010101_10010100_11101001_0;
      patterns[21911] = 25'b01010101_10010101_11101010_0;
      patterns[21912] = 25'b01010101_10010110_11101011_0;
      patterns[21913] = 25'b01010101_10010111_11101100_0;
      patterns[21914] = 25'b01010101_10011000_11101101_0;
      patterns[21915] = 25'b01010101_10011001_11101110_0;
      patterns[21916] = 25'b01010101_10011010_11101111_0;
      patterns[21917] = 25'b01010101_10011011_11110000_0;
      patterns[21918] = 25'b01010101_10011100_11110001_0;
      patterns[21919] = 25'b01010101_10011101_11110010_0;
      patterns[21920] = 25'b01010101_10011110_11110011_0;
      patterns[21921] = 25'b01010101_10011111_11110100_0;
      patterns[21922] = 25'b01010101_10100000_11110101_0;
      patterns[21923] = 25'b01010101_10100001_11110110_0;
      patterns[21924] = 25'b01010101_10100010_11110111_0;
      patterns[21925] = 25'b01010101_10100011_11111000_0;
      patterns[21926] = 25'b01010101_10100100_11111001_0;
      patterns[21927] = 25'b01010101_10100101_11111010_0;
      patterns[21928] = 25'b01010101_10100110_11111011_0;
      patterns[21929] = 25'b01010101_10100111_11111100_0;
      patterns[21930] = 25'b01010101_10101000_11111101_0;
      patterns[21931] = 25'b01010101_10101001_11111110_0;
      patterns[21932] = 25'b01010101_10101010_11111111_0;
      patterns[21933] = 25'b01010101_10101011_00000000_1;
      patterns[21934] = 25'b01010101_10101100_00000001_1;
      patterns[21935] = 25'b01010101_10101101_00000010_1;
      patterns[21936] = 25'b01010101_10101110_00000011_1;
      patterns[21937] = 25'b01010101_10101111_00000100_1;
      patterns[21938] = 25'b01010101_10110000_00000101_1;
      patterns[21939] = 25'b01010101_10110001_00000110_1;
      patterns[21940] = 25'b01010101_10110010_00000111_1;
      patterns[21941] = 25'b01010101_10110011_00001000_1;
      patterns[21942] = 25'b01010101_10110100_00001001_1;
      patterns[21943] = 25'b01010101_10110101_00001010_1;
      patterns[21944] = 25'b01010101_10110110_00001011_1;
      patterns[21945] = 25'b01010101_10110111_00001100_1;
      patterns[21946] = 25'b01010101_10111000_00001101_1;
      patterns[21947] = 25'b01010101_10111001_00001110_1;
      patterns[21948] = 25'b01010101_10111010_00001111_1;
      patterns[21949] = 25'b01010101_10111011_00010000_1;
      patterns[21950] = 25'b01010101_10111100_00010001_1;
      patterns[21951] = 25'b01010101_10111101_00010010_1;
      patterns[21952] = 25'b01010101_10111110_00010011_1;
      patterns[21953] = 25'b01010101_10111111_00010100_1;
      patterns[21954] = 25'b01010101_11000000_00010101_1;
      patterns[21955] = 25'b01010101_11000001_00010110_1;
      patterns[21956] = 25'b01010101_11000010_00010111_1;
      patterns[21957] = 25'b01010101_11000011_00011000_1;
      patterns[21958] = 25'b01010101_11000100_00011001_1;
      patterns[21959] = 25'b01010101_11000101_00011010_1;
      patterns[21960] = 25'b01010101_11000110_00011011_1;
      patterns[21961] = 25'b01010101_11000111_00011100_1;
      patterns[21962] = 25'b01010101_11001000_00011101_1;
      patterns[21963] = 25'b01010101_11001001_00011110_1;
      patterns[21964] = 25'b01010101_11001010_00011111_1;
      patterns[21965] = 25'b01010101_11001011_00100000_1;
      patterns[21966] = 25'b01010101_11001100_00100001_1;
      patterns[21967] = 25'b01010101_11001101_00100010_1;
      patterns[21968] = 25'b01010101_11001110_00100011_1;
      patterns[21969] = 25'b01010101_11001111_00100100_1;
      patterns[21970] = 25'b01010101_11010000_00100101_1;
      patterns[21971] = 25'b01010101_11010001_00100110_1;
      patterns[21972] = 25'b01010101_11010010_00100111_1;
      patterns[21973] = 25'b01010101_11010011_00101000_1;
      patterns[21974] = 25'b01010101_11010100_00101001_1;
      patterns[21975] = 25'b01010101_11010101_00101010_1;
      patterns[21976] = 25'b01010101_11010110_00101011_1;
      patterns[21977] = 25'b01010101_11010111_00101100_1;
      patterns[21978] = 25'b01010101_11011000_00101101_1;
      patterns[21979] = 25'b01010101_11011001_00101110_1;
      patterns[21980] = 25'b01010101_11011010_00101111_1;
      patterns[21981] = 25'b01010101_11011011_00110000_1;
      patterns[21982] = 25'b01010101_11011100_00110001_1;
      patterns[21983] = 25'b01010101_11011101_00110010_1;
      patterns[21984] = 25'b01010101_11011110_00110011_1;
      patterns[21985] = 25'b01010101_11011111_00110100_1;
      patterns[21986] = 25'b01010101_11100000_00110101_1;
      patterns[21987] = 25'b01010101_11100001_00110110_1;
      patterns[21988] = 25'b01010101_11100010_00110111_1;
      patterns[21989] = 25'b01010101_11100011_00111000_1;
      patterns[21990] = 25'b01010101_11100100_00111001_1;
      patterns[21991] = 25'b01010101_11100101_00111010_1;
      patterns[21992] = 25'b01010101_11100110_00111011_1;
      patterns[21993] = 25'b01010101_11100111_00111100_1;
      patterns[21994] = 25'b01010101_11101000_00111101_1;
      patterns[21995] = 25'b01010101_11101001_00111110_1;
      patterns[21996] = 25'b01010101_11101010_00111111_1;
      patterns[21997] = 25'b01010101_11101011_01000000_1;
      patterns[21998] = 25'b01010101_11101100_01000001_1;
      patterns[21999] = 25'b01010101_11101101_01000010_1;
      patterns[22000] = 25'b01010101_11101110_01000011_1;
      patterns[22001] = 25'b01010101_11101111_01000100_1;
      patterns[22002] = 25'b01010101_11110000_01000101_1;
      patterns[22003] = 25'b01010101_11110001_01000110_1;
      patterns[22004] = 25'b01010101_11110010_01000111_1;
      patterns[22005] = 25'b01010101_11110011_01001000_1;
      patterns[22006] = 25'b01010101_11110100_01001001_1;
      patterns[22007] = 25'b01010101_11110101_01001010_1;
      patterns[22008] = 25'b01010101_11110110_01001011_1;
      patterns[22009] = 25'b01010101_11110111_01001100_1;
      patterns[22010] = 25'b01010101_11111000_01001101_1;
      patterns[22011] = 25'b01010101_11111001_01001110_1;
      patterns[22012] = 25'b01010101_11111010_01001111_1;
      patterns[22013] = 25'b01010101_11111011_01010000_1;
      patterns[22014] = 25'b01010101_11111100_01010001_1;
      patterns[22015] = 25'b01010101_11111101_01010010_1;
      patterns[22016] = 25'b01010101_11111110_01010011_1;
      patterns[22017] = 25'b01010101_11111111_01010100_1;
      patterns[22018] = 25'b01010110_00000000_01010110_0;
      patterns[22019] = 25'b01010110_00000001_01010111_0;
      patterns[22020] = 25'b01010110_00000010_01011000_0;
      patterns[22021] = 25'b01010110_00000011_01011001_0;
      patterns[22022] = 25'b01010110_00000100_01011010_0;
      patterns[22023] = 25'b01010110_00000101_01011011_0;
      patterns[22024] = 25'b01010110_00000110_01011100_0;
      patterns[22025] = 25'b01010110_00000111_01011101_0;
      patterns[22026] = 25'b01010110_00001000_01011110_0;
      patterns[22027] = 25'b01010110_00001001_01011111_0;
      patterns[22028] = 25'b01010110_00001010_01100000_0;
      patterns[22029] = 25'b01010110_00001011_01100001_0;
      patterns[22030] = 25'b01010110_00001100_01100010_0;
      patterns[22031] = 25'b01010110_00001101_01100011_0;
      patterns[22032] = 25'b01010110_00001110_01100100_0;
      patterns[22033] = 25'b01010110_00001111_01100101_0;
      patterns[22034] = 25'b01010110_00010000_01100110_0;
      patterns[22035] = 25'b01010110_00010001_01100111_0;
      patterns[22036] = 25'b01010110_00010010_01101000_0;
      patterns[22037] = 25'b01010110_00010011_01101001_0;
      patterns[22038] = 25'b01010110_00010100_01101010_0;
      patterns[22039] = 25'b01010110_00010101_01101011_0;
      patterns[22040] = 25'b01010110_00010110_01101100_0;
      patterns[22041] = 25'b01010110_00010111_01101101_0;
      patterns[22042] = 25'b01010110_00011000_01101110_0;
      patterns[22043] = 25'b01010110_00011001_01101111_0;
      patterns[22044] = 25'b01010110_00011010_01110000_0;
      patterns[22045] = 25'b01010110_00011011_01110001_0;
      patterns[22046] = 25'b01010110_00011100_01110010_0;
      patterns[22047] = 25'b01010110_00011101_01110011_0;
      patterns[22048] = 25'b01010110_00011110_01110100_0;
      patterns[22049] = 25'b01010110_00011111_01110101_0;
      patterns[22050] = 25'b01010110_00100000_01110110_0;
      patterns[22051] = 25'b01010110_00100001_01110111_0;
      patterns[22052] = 25'b01010110_00100010_01111000_0;
      patterns[22053] = 25'b01010110_00100011_01111001_0;
      patterns[22054] = 25'b01010110_00100100_01111010_0;
      patterns[22055] = 25'b01010110_00100101_01111011_0;
      patterns[22056] = 25'b01010110_00100110_01111100_0;
      patterns[22057] = 25'b01010110_00100111_01111101_0;
      patterns[22058] = 25'b01010110_00101000_01111110_0;
      patterns[22059] = 25'b01010110_00101001_01111111_0;
      patterns[22060] = 25'b01010110_00101010_10000000_0;
      patterns[22061] = 25'b01010110_00101011_10000001_0;
      patterns[22062] = 25'b01010110_00101100_10000010_0;
      patterns[22063] = 25'b01010110_00101101_10000011_0;
      patterns[22064] = 25'b01010110_00101110_10000100_0;
      patterns[22065] = 25'b01010110_00101111_10000101_0;
      patterns[22066] = 25'b01010110_00110000_10000110_0;
      patterns[22067] = 25'b01010110_00110001_10000111_0;
      patterns[22068] = 25'b01010110_00110010_10001000_0;
      patterns[22069] = 25'b01010110_00110011_10001001_0;
      patterns[22070] = 25'b01010110_00110100_10001010_0;
      patterns[22071] = 25'b01010110_00110101_10001011_0;
      patterns[22072] = 25'b01010110_00110110_10001100_0;
      patterns[22073] = 25'b01010110_00110111_10001101_0;
      patterns[22074] = 25'b01010110_00111000_10001110_0;
      patterns[22075] = 25'b01010110_00111001_10001111_0;
      patterns[22076] = 25'b01010110_00111010_10010000_0;
      patterns[22077] = 25'b01010110_00111011_10010001_0;
      patterns[22078] = 25'b01010110_00111100_10010010_0;
      patterns[22079] = 25'b01010110_00111101_10010011_0;
      patterns[22080] = 25'b01010110_00111110_10010100_0;
      patterns[22081] = 25'b01010110_00111111_10010101_0;
      patterns[22082] = 25'b01010110_01000000_10010110_0;
      patterns[22083] = 25'b01010110_01000001_10010111_0;
      patterns[22084] = 25'b01010110_01000010_10011000_0;
      patterns[22085] = 25'b01010110_01000011_10011001_0;
      patterns[22086] = 25'b01010110_01000100_10011010_0;
      patterns[22087] = 25'b01010110_01000101_10011011_0;
      patterns[22088] = 25'b01010110_01000110_10011100_0;
      patterns[22089] = 25'b01010110_01000111_10011101_0;
      patterns[22090] = 25'b01010110_01001000_10011110_0;
      patterns[22091] = 25'b01010110_01001001_10011111_0;
      patterns[22092] = 25'b01010110_01001010_10100000_0;
      patterns[22093] = 25'b01010110_01001011_10100001_0;
      patterns[22094] = 25'b01010110_01001100_10100010_0;
      patterns[22095] = 25'b01010110_01001101_10100011_0;
      patterns[22096] = 25'b01010110_01001110_10100100_0;
      patterns[22097] = 25'b01010110_01001111_10100101_0;
      patterns[22098] = 25'b01010110_01010000_10100110_0;
      patterns[22099] = 25'b01010110_01010001_10100111_0;
      patterns[22100] = 25'b01010110_01010010_10101000_0;
      patterns[22101] = 25'b01010110_01010011_10101001_0;
      patterns[22102] = 25'b01010110_01010100_10101010_0;
      patterns[22103] = 25'b01010110_01010101_10101011_0;
      patterns[22104] = 25'b01010110_01010110_10101100_0;
      patterns[22105] = 25'b01010110_01010111_10101101_0;
      patterns[22106] = 25'b01010110_01011000_10101110_0;
      patterns[22107] = 25'b01010110_01011001_10101111_0;
      patterns[22108] = 25'b01010110_01011010_10110000_0;
      patterns[22109] = 25'b01010110_01011011_10110001_0;
      patterns[22110] = 25'b01010110_01011100_10110010_0;
      patterns[22111] = 25'b01010110_01011101_10110011_0;
      patterns[22112] = 25'b01010110_01011110_10110100_0;
      patterns[22113] = 25'b01010110_01011111_10110101_0;
      patterns[22114] = 25'b01010110_01100000_10110110_0;
      patterns[22115] = 25'b01010110_01100001_10110111_0;
      patterns[22116] = 25'b01010110_01100010_10111000_0;
      patterns[22117] = 25'b01010110_01100011_10111001_0;
      patterns[22118] = 25'b01010110_01100100_10111010_0;
      patterns[22119] = 25'b01010110_01100101_10111011_0;
      patterns[22120] = 25'b01010110_01100110_10111100_0;
      patterns[22121] = 25'b01010110_01100111_10111101_0;
      patterns[22122] = 25'b01010110_01101000_10111110_0;
      patterns[22123] = 25'b01010110_01101001_10111111_0;
      patterns[22124] = 25'b01010110_01101010_11000000_0;
      patterns[22125] = 25'b01010110_01101011_11000001_0;
      patterns[22126] = 25'b01010110_01101100_11000010_0;
      patterns[22127] = 25'b01010110_01101101_11000011_0;
      patterns[22128] = 25'b01010110_01101110_11000100_0;
      patterns[22129] = 25'b01010110_01101111_11000101_0;
      patterns[22130] = 25'b01010110_01110000_11000110_0;
      patterns[22131] = 25'b01010110_01110001_11000111_0;
      patterns[22132] = 25'b01010110_01110010_11001000_0;
      patterns[22133] = 25'b01010110_01110011_11001001_0;
      patterns[22134] = 25'b01010110_01110100_11001010_0;
      patterns[22135] = 25'b01010110_01110101_11001011_0;
      patterns[22136] = 25'b01010110_01110110_11001100_0;
      patterns[22137] = 25'b01010110_01110111_11001101_0;
      patterns[22138] = 25'b01010110_01111000_11001110_0;
      patterns[22139] = 25'b01010110_01111001_11001111_0;
      patterns[22140] = 25'b01010110_01111010_11010000_0;
      patterns[22141] = 25'b01010110_01111011_11010001_0;
      patterns[22142] = 25'b01010110_01111100_11010010_0;
      patterns[22143] = 25'b01010110_01111101_11010011_0;
      patterns[22144] = 25'b01010110_01111110_11010100_0;
      patterns[22145] = 25'b01010110_01111111_11010101_0;
      patterns[22146] = 25'b01010110_10000000_11010110_0;
      patterns[22147] = 25'b01010110_10000001_11010111_0;
      patterns[22148] = 25'b01010110_10000010_11011000_0;
      patterns[22149] = 25'b01010110_10000011_11011001_0;
      patterns[22150] = 25'b01010110_10000100_11011010_0;
      patterns[22151] = 25'b01010110_10000101_11011011_0;
      patterns[22152] = 25'b01010110_10000110_11011100_0;
      patterns[22153] = 25'b01010110_10000111_11011101_0;
      patterns[22154] = 25'b01010110_10001000_11011110_0;
      patterns[22155] = 25'b01010110_10001001_11011111_0;
      patterns[22156] = 25'b01010110_10001010_11100000_0;
      patterns[22157] = 25'b01010110_10001011_11100001_0;
      patterns[22158] = 25'b01010110_10001100_11100010_0;
      patterns[22159] = 25'b01010110_10001101_11100011_0;
      patterns[22160] = 25'b01010110_10001110_11100100_0;
      patterns[22161] = 25'b01010110_10001111_11100101_0;
      patterns[22162] = 25'b01010110_10010000_11100110_0;
      patterns[22163] = 25'b01010110_10010001_11100111_0;
      patterns[22164] = 25'b01010110_10010010_11101000_0;
      patterns[22165] = 25'b01010110_10010011_11101001_0;
      patterns[22166] = 25'b01010110_10010100_11101010_0;
      patterns[22167] = 25'b01010110_10010101_11101011_0;
      patterns[22168] = 25'b01010110_10010110_11101100_0;
      patterns[22169] = 25'b01010110_10010111_11101101_0;
      patterns[22170] = 25'b01010110_10011000_11101110_0;
      patterns[22171] = 25'b01010110_10011001_11101111_0;
      patterns[22172] = 25'b01010110_10011010_11110000_0;
      patterns[22173] = 25'b01010110_10011011_11110001_0;
      patterns[22174] = 25'b01010110_10011100_11110010_0;
      patterns[22175] = 25'b01010110_10011101_11110011_0;
      patterns[22176] = 25'b01010110_10011110_11110100_0;
      patterns[22177] = 25'b01010110_10011111_11110101_0;
      patterns[22178] = 25'b01010110_10100000_11110110_0;
      patterns[22179] = 25'b01010110_10100001_11110111_0;
      patterns[22180] = 25'b01010110_10100010_11111000_0;
      patterns[22181] = 25'b01010110_10100011_11111001_0;
      patterns[22182] = 25'b01010110_10100100_11111010_0;
      patterns[22183] = 25'b01010110_10100101_11111011_0;
      patterns[22184] = 25'b01010110_10100110_11111100_0;
      patterns[22185] = 25'b01010110_10100111_11111101_0;
      patterns[22186] = 25'b01010110_10101000_11111110_0;
      patterns[22187] = 25'b01010110_10101001_11111111_0;
      patterns[22188] = 25'b01010110_10101010_00000000_1;
      patterns[22189] = 25'b01010110_10101011_00000001_1;
      patterns[22190] = 25'b01010110_10101100_00000010_1;
      patterns[22191] = 25'b01010110_10101101_00000011_1;
      patterns[22192] = 25'b01010110_10101110_00000100_1;
      patterns[22193] = 25'b01010110_10101111_00000101_1;
      patterns[22194] = 25'b01010110_10110000_00000110_1;
      patterns[22195] = 25'b01010110_10110001_00000111_1;
      patterns[22196] = 25'b01010110_10110010_00001000_1;
      patterns[22197] = 25'b01010110_10110011_00001001_1;
      patterns[22198] = 25'b01010110_10110100_00001010_1;
      patterns[22199] = 25'b01010110_10110101_00001011_1;
      patterns[22200] = 25'b01010110_10110110_00001100_1;
      patterns[22201] = 25'b01010110_10110111_00001101_1;
      patterns[22202] = 25'b01010110_10111000_00001110_1;
      patterns[22203] = 25'b01010110_10111001_00001111_1;
      patterns[22204] = 25'b01010110_10111010_00010000_1;
      patterns[22205] = 25'b01010110_10111011_00010001_1;
      patterns[22206] = 25'b01010110_10111100_00010010_1;
      patterns[22207] = 25'b01010110_10111101_00010011_1;
      patterns[22208] = 25'b01010110_10111110_00010100_1;
      patterns[22209] = 25'b01010110_10111111_00010101_1;
      patterns[22210] = 25'b01010110_11000000_00010110_1;
      patterns[22211] = 25'b01010110_11000001_00010111_1;
      patterns[22212] = 25'b01010110_11000010_00011000_1;
      patterns[22213] = 25'b01010110_11000011_00011001_1;
      patterns[22214] = 25'b01010110_11000100_00011010_1;
      patterns[22215] = 25'b01010110_11000101_00011011_1;
      patterns[22216] = 25'b01010110_11000110_00011100_1;
      patterns[22217] = 25'b01010110_11000111_00011101_1;
      patterns[22218] = 25'b01010110_11001000_00011110_1;
      patterns[22219] = 25'b01010110_11001001_00011111_1;
      patterns[22220] = 25'b01010110_11001010_00100000_1;
      patterns[22221] = 25'b01010110_11001011_00100001_1;
      patterns[22222] = 25'b01010110_11001100_00100010_1;
      patterns[22223] = 25'b01010110_11001101_00100011_1;
      patterns[22224] = 25'b01010110_11001110_00100100_1;
      patterns[22225] = 25'b01010110_11001111_00100101_1;
      patterns[22226] = 25'b01010110_11010000_00100110_1;
      patterns[22227] = 25'b01010110_11010001_00100111_1;
      patterns[22228] = 25'b01010110_11010010_00101000_1;
      patterns[22229] = 25'b01010110_11010011_00101001_1;
      patterns[22230] = 25'b01010110_11010100_00101010_1;
      patterns[22231] = 25'b01010110_11010101_00101011_1;
      patterns[22232] = 25'b01010110_11010110_00101100_1;
      patterns[22233] = 25'b01010110_11010111_00101101_1;
      patterns[22234] = 25'b01010110_11011000_00101110_1;
      patterns[22235] = 25'b01010110_11011001_00101111_1;
      patterns[22236] = 25'b01010110_11011010_00110000_1;
      patterns[22237] = 25'b01010110_11011011_00110001_1;
      patterns[22238] = 25'b01010110_11011100_00110010_1;
      patterns[22239] = 25'b01010110_11011101_00110011_1;
      patterns[22240] = 25'b01010110_11011110_00110100_1;
      patterns[22241] = 25'b01010110_11011111_00110101_1;
      patterns[22242] = 25'b01010110_11100000_00110110_1;
      patterns[22243] = 25'b01010110_11100001_00110111_1;
      patterns[22244] = 25'b01010110_11100010_00111000_1;
      patterns[22245] = 25'b01010110_11100011_00111001_1;
      patterns[22246] = 25'b01010110_11100100_00111010_1;
      patterns[22247] = 25'b01010110_11100101_00111011_1;
      patterns[22248] = 25'b01010110_11100110_00111100_1;
      patterns[22249] = 25'b01010110_11100111_00111101_1;
      patterns[22250] = 25'b01010110_11101000_00111110_1;
      patterns[22251] = 25'b01010110_11101001_00111111_1;
      patterns[22252] = 25'b01010110_11101010_01000000_1;
      patterns[22253] = 25'b01010110_11101011_01000001_1;
      patterns[22254] = 25'b01010110_11101100_01000010_1;
      patterns[22255] = 25'b01010110_11101101_01000011_1;
      patterns[22256] = 25'b01010110_11101110_01000100_1;
      patterns[22257] = 25'b01010110_11101111_01000101_1;
      patterns[22258] = 25'b01010110_11110000_01000110_1;
      patterns[22259] = 25'b01010110_11110001_01000111_1;
      patterns[22260] = 25'b01010110_11110010_01001000_1;
      patterns[22261] = 25'b01010110_11110011_01001001_1;
      patterns[22262] = 25'b01010110_11110100_01001010_1;
      patterns[22263] = 25'b01010110_11110101_01001011_1;
      patterns[22264] = 25'b01010110_11110110_01001100_1;
      patterns[22265] = 25'b01010110_11110111_01001101_1;
      patterns[22266] = 25'b01010110_11111000_01001110_1;
      patterns[22267] = 25'b01010110_11111001_01001111_1;
      patterns[22268] = 25'b01010110_11111010_01010000_1;
      patterns[22269] = 25'b01010110_11111011_01010001_1;
      patterns[22270] = 25'b01010110_11111100_01010010_1;
      patterns[22271] = 25'b01010110_11111101_01010011_1;
      patterns[22272] = 25'b01010110_11111110_01010100_1;
      patterns[22273] = 25'b01010110_11111111_01010101_1;
      patterns[22274] = 25'b01010111_00000000_01010111_0;
      patterns[22275] = 25'b01010111_00000001_01011000_0;
      patterns[22276] = 25'b01010111_00000010_01011001_0;
      patterns[22277] = 25'b01010111_00000011_01011010_0;
      patterns[22278] = 25'b01010111_00000100_01011011_0;
      patterns[22279] = 25'b01010111_00000101_01011100_0;
      patterns[22280] = 25'b01010111_00000110_01011101_0;
      patterns[22281] = 25'b01010111_00000111_01011110_0;
      patterns[22282] = 25'b01010111_00001000_01011111_0;
      patterns[22283] = 25'b01010111_00001001_01100000_0;
      patterns[22284] = 25'b01010111_00001010_01100001_0;
      patterns[22285] = 25'b01010111_00001011_01100010_0;
      patterns[22286] = 25'b01010111_00001100_01100011_0;
      patterns[22287] = 25'b01010111_00001101_01100100_0;
      patterns[22288] = 25'b01010111_00001110_01100101_0;
      patterns[22289] = 25'b01010111_00001111_01100110_0;
      patterns[22290] = 25'b01010111_00010000_01100111_0;
      patterns[22291] = 25'b01010111_00010001_01101000_0;
      patterns[22292] = 25'b01010111_00010010_01101001_0;
      patterns[22293] = 25'b01010111_00010011_01101010_0;
      patterns[22294] = 25'b01010111_00010100_01101011_0;
      patterns[22295] = 25'b01010111_00010101_01101100_0;
      patterns[22296] = 25'b01010111_00010110_01101101_0;
      patterns[22297] = 25'b01010111_00010111_01101110_0;
      patterns[22298] = 25'b01010111_00011000_01101111_0;
      patterns[22299] = 25'b01010111_00011001_01110000_0;
      patterns[22300] = 25'b01010111_00011010_01110001_0;
      patterns[22301] = 25'b01010111_00011011_01110010_0;
      patterns[22302] = 25'b01010111_00011100_01110011_0;
      patterns[22303] = 25'b01010111_00011101_01110100_0;
      patterns[22304] = 25'b01010111_00011110_01110101_0;
      patterns[22305] = 25'b01010111_00011111_01110110_0;
      patterns[22306] = 25'b01010111_00100000_01110111_0;
      patterns[22307] = 25'b01010111_00100001_01111000_0;
      patterns[22308] = 25'b01010111_00100010_01111001_0;
      patterns[22309] = 25'b01010111_00100011_01111010_0;
      patterns[22310] = 25'b01010111_00100100_01111011_0;
      patterns[22311] = 25'b01010111_00100101_01111100_0;
      patterns[22312] = 25'b01010111_00100110_01111101_0;
      patterns[22313] = 25'b01010111_00100111_01111110_0;
      patterns[22314] = 25'b01010111_00101000_01111111_0;
      patterns[22315] = 25'b01010111_00101001_10000000_0;
      patterns[22316] = 25'b01010111_00101010_10000001_0;
      patterns[22317] = 25'b01010111_00101011_10000010_0;
      patterns[22318] = 25'b01010111_00101100_10000011_0;
      patterns[22319] = 25'b01010111_00101101_10000100_0;
      patterns[22320] = 25'b01010111_00101110_10000101_0;
      patterns[22321] = 25'b01010111_00101111_10000110_0;
      patterns[22322] = 25'b01010111_00110000_10000111_0;
      patterns[22323] = 25'b01010111_00110001_10001000_0;
      patterns[22324] = 25'b01010111_00110010_10001001_0;
      patterns[22325] = 25'b01010111_00110011_10001010_0;
      patterns[22326] = 25'b01010111_00110100_10001011_0;
      patterns[22327] = 25'b01010111_00110101_10001100_0;
      patterns[22328] = 25'b01010111_00110110_10001101_0;
      patterns[22329] = 25'b01010111_00110111_10001110_0;
      patterns[22330] = 25'b01010111_00111000_10001111_0;
      patterns[22331] = 25'b01010111_00111001_10010000_0;
      patterns[22332] = 25'b01010111_00111010_10010001_0;
      patterns[22333] = 25'b01010111_00111011_10010010_0;
      patterns[22334] = 25'b01010111_00111100_10010011_0;
      patterns[22335] = 25'b01010111_00111101_10010100_0;
      patterns[22336] = 25'b01010111_00111110_10010101_0;
      patterns[22337] = 25'b01010111_00111111_10010110_0;
      patterns[22338] = 25'b01010111_01000000_10010111_0;
      patterns[22339] = 25'b01010111_01000001_10011000_0;
      patterns[22340] = 25'b01010111_01000010_10011001_0;
      patterns[22341] = 25'b01010111_01000011_10011010_0;
      patterns[22342] = 25'b01010111_01000100_10011011_0;
      patterns[22343] = 25'b01010111_01000101_10011100_0;
      patterns[22344] = 25'b01010111_01000110_10011101_0;
      patterns[22345] = 25'b01010111_01000111_10011110_0;
      patterns[22346] = 25'b01010111_01001000_10011111_0;
      patterns[22347] = 25'b01010111_01001001_10100000_0;
      patterns[22348] = 25'b01010111_01001010_10100001_0;
      patterns[22349] = 25'b01010111_01001011_10100010_0;
      patterns[22350] = 25'b01010111_01001100_10100011_0;
      patterns[22351] = 25'b01010111_01001101_10100100_0;
      patterns[22352] = 25'b01010111_01001110_10100101_0;
      patterns[22353] = 25'b01010111_01001111_10100110_0;
      patterns[22354] = 25'b01010111_01010000_10100111_0;
      patterns[22355] = 25'b01010111_01010001_10101000_0;
      patterns[22356] = 25'b01010111_01010010_10101001_0;
      patterns[22357] = 25'b01010111_01010011_10101010_0;
      patterns[22358] = 25'b01010111_01010100_10101011_0;
      patterns[22359] = 25'b01010111_01010101_10101100_0;
      patterns[22360] = 25'b01010111_01010110_10101101_0;
      patterns[22361] = 25'b01010111_01010111_10101110_0;
      patterns[22362] = 25'b01010111_01011000_10101111_0;
      patterns[22363] = 25'b01010111_01011001_10110000_0;
      patterns[22364] = 25'b01010111_01011010_10110001_0;
      patterns[22365] = 25'b01010111_01011011_10110010_0;
      patterns[22366] = 25'b01010111_01011100_10110011_0;
      patterns[22367] = 25'b01010111_01011101_10110100_0;
      patterns[22368] = 25'b01010111_01011110_10110101_0;
      patterns[22369] = 25'b01010111_01011111_10110110_0;
      patterns[22370] = 25'b01010111_01100000_10110111_0;
      patterns[22371] = 25'b01010111_01100001_10111000_0;
      patterns[22372] = 25'b01010111_01100010_10111001_0;
      patterns[22373] = 25'b01010111_01100011_10111010_0;
      patterns[22374] = 25'b01010111_01100100_10111011_0;
      patterns[22375] = 25'b01010111_01100101_10111100_0;
      patterns[22376] = 25'b01010111_01100110_10111101_0;
      patterns[22377] = 25'b01010111_01100111_10111110_0;
      patterns[22378] = 25'b01010111_01101000_10111111_0;
      patterns[22379] = 25'b01010111_01101001_11000000_0;
      patterns[22380] = 25'b01010111_01101010_11000001_0;
      patterns[22381] = 25'b01010111_01101011_11000010_0;
      patterns[22382] = 25'b01010111_01101100_11000011_0;
      patterns[22383] = 25'b01010111_01101101_11000100_0;
      patterns[22384] = 25'b01010111_01101110_11000101_0;
      patterns[22385] = 25'b01010111_01101111_11000110_0;
      patterns[22386] = 25'b01010111_01110000_11000111_0;
      patterns[22387] = 25'b01010111_01110001_11001000_0;
      patterns[22388] = 25'b01010111_01110010_11001001_0;
      patterns[22389] = 25'b01010111_01110011_11001010_0;
      patterns[22390] = 25'b01010111_01110100_11001011_0;
      patterns[22391] = 25'b01010111_01110101_11001100_0;
      patterns[22392] = 25'b01010111_01110110_11001101_0;
      patterns[22393] = 25'b01010111_01110111_11001110_0;
      patterns[22394] = 25'b01010111_01111000_11001111_0;
      patterns[22395] = 25'b01010111_01111001_11010000_0;
      patterns[22396] = 25'b01010111_01111010_11010001_0;
      patterns[22397] = 25'b01010111_01111011_11010010_0;
      patterns[22398] = 25'b01010111_01111100_11010011_0;
      patterns[22399] = 25'b01010111_01111101_11010100_0;
      patterns[22400] = 25'b01010111_01111110_11010101_0;
      patterns[22401] = 25'b01010111_01111111_11010110_0;
      patterns[22402] = 25'b01010111_10000000_11010111_0;
      patterns[22403] = 25'b01010111_10000001_11011000_0;
      patterns[22404] = 25'b01010111_10000010_11011001_0;
      patterns[22405] = 25'b01010111_10000011_11011010_0;
      patterns[22406] = 25'b01010111_10000100_11011011_0;
      patterns[22407] = 25'b01010111_10000101_11011100_0;
      patterns[22408] = 25'b01010111_10000110_11011101_0;
      patterns[22409] = 25'b01010111_10000111_11011110_0;
      patterns[22410] = 25'b01010111_10001000_11011111_0;
      patterns[22411] = 25'b01010111_10001001_11100000_0;
      patterns[22412] = 25'b01010111_10001010_11100001_0;
      patterns[22413] = 25'b01010111_10001011_11100010_0;
      patterns[22414] = 25'b01010111_10001100_11100011_0;
      patterns[22415] = 25'b01010111_10001101_11100100_0;
      patterns[22416] = 25'b01010111_10001110_11100101_0;
      patterns[22417] = 25'b01010111_10001111_11100110_0;
      patterns[22418] = 25'b01010111_10010000_11100111_0;
      patterns[22419] = 25'b01010111_10010001_11101000_0;
      patterns[22420] = 25'b01010111_10010010_11101001_0;
      patterns[22421] = 25'b01010111_10010011_11101010_0;
      patterns[22422] = 25'b01010111_10010100_11101011_0;
      patterns[22423] = 25'b01010111_10010101_11101100_0;
      patterns[22424] = 25'b01010111_10010110_11101101_0;
      patterns[22425] = 25'b01010111_10010111_11101110_0;
      patterns[22426] = 25'b01010111_10011000_11101111_0;
      patterns[22427] = 25'b01010111_10011001_11110000_0;
      patterns[22428] = 25'b01010111_10011010_11110001_0;
      patterns[22429] = 25'b01010111_10011011_11110010_0;
      patterns[22430] = 25'b01010111_10011100_11110011_0;
      patterns[22431] = 25'b01010111_10011101_11110100_0;
      patterns[22432] = 25'b01010111_10011110_11110101_0;
      patterns[22433] = 25'b01010111_10011111_11110110_0;
      patterns[22434] = 25'b01010111_10100000_11110111_0;
      patterns[22435] = 25'b01010111_10100001_11111000_0;
      patterns[22436] = 25'b01010111_10100010_11111001_0;
      patterns[22437] = 25'b01010111_10100011_11111010_0;
      patterns[22438] = 25'b01010111_10100100_11111011_0;
      patterns[22439] = 25'b01010111_10100101_11111100_0;
      patterns[22440] = 25'b01010111_10100110_11111101_0;
      patterns[22441] = 25'b01010111_10100111_11111110_0;
      patterns[22442] = 25'b01010111_10101000_11111111_0;
      patterns[22443] = 25'b01010111_10101001_00000000_1;
      patterns[22444] = 25'b01010111_10101010_00000001_1;
      patterns[22445] = 25'b01010111_10101011_00000010_1;
      patterns[22446] = 25'b01010111_10101100_00000011_1;
      patterns[22447] = 25'b01010111_10101101_00000100_1;
      patterns[22448] = 25'b01010111_10101110_00000101_1;
      patterns[22449] = 25'b01010111_10101111_00000110_1;
      patterns[22450] = 25'b01010111_10110000_00000111_1;
      patterns[22451] = 25'b01010111_10110001_00001000_1;
      patterns[22452] = 25'b01010111_10110010_00001001_1;
      patterns[22453] = 25'b01010111_10110011_00001010_1;
      patterns[22454] = 25'b01010111_10110100_00001011_1;
      patterns[22455] = 25'b01010111_10110101_00001100_1;
      patterns[22456] = 25'b01010111_10110110_00001101_1;
      patterns[22457] = 25'b01010111_10110111_00001110_1;
      patterns[22458] = 25'b01010111_10111000_00001111_1;
      patterns[22459] = 25'b01010111_10111001_00010000_1;
      patterns[22460] = 25'b01010111_10111010_00010001_1;
      patterns[22461] = 25'b01010111_10111011_00010010_1;
      patterns[22462] = 25'b01010111_10111100_00010011_1;
      patterns[22463] = 25'b01010111_10111101_00010100_1;
      patterns[22464] = 25'b01010111_10111110_00010101_1;
      patterns[22465] = 25'b01010111_10111111_00010110_1;
      patterns[22466] = 25'b01010111_11000000_00010111_1;
      patterns[22467] = 25'b01010111_11000001_00011000_1;
      patterns[22468] = 25'b01010111_11000010_00011001_1;
      patterns[22469] = 25'b01010111_11000011_00011010_1;
      patterns[22470] = 25'b01010111_11000100_00011011_1;
      patterns[22471] = 25'b01010111_11000101_00011100_1;
      patterns[22472] = 25'b01010111_11000110_00011101_1;
      patterns[22473] = 25'b01010111_11000111_00011110_1;
      patterns[22474] = 25'b01010111_11001000_00011111_1;
      patterns[22475] = 25'b01010111_11001001_00100000_1;
      patterns[22476] = 25'b01010111_11001010_00100001_1;
      patterns[22477] = 25'b01010111_11001011_00100010_1;
      patterns[22478] = 25'b01010111_11001100_00100011_1;
      patterns[22479] = 25'b01010111_11001101_00100100_1;
      patterns[22480] = 25'b01010111_11001110_00100101_1;
      patterns[22481] = 25'b01010111_11001111_00100110_1;
      patterns[22482] = 25'b01010111_11010000_00100111_1;
      patterns[22483] = 25'b01010111_11010001_00101000_1;
      patterns[22484] = 25'b01010111_11010010_00101001_1;
      patterns[22485] = 25'b01010111_11010011_00101010_1;
      patterns[22486] = 25'b01010111_11010100_00101011_1;
      patterns[22487] = 25'b01010111_11010101_00101100_1;
      patterns[22488] = 25'b01010111_11010110_00101101_1;
      patterns[22489] = 25'b01010111_11010111_00101110_1;
      patterns[22490] = 25'b01010111_11011000_00101111_1;
      patterns[22491] = 25'b01010111_11011001_00110000_1;
      patterns[22492] = 25'b01010111_11011010_00110001_1;
      patterns[22493] = 25'b01010111_11011011_00110010_1;
      patterns[22494] = 25'b01010111_11011100_00110011_1;
      patterns[22495] = 25'b01010111_11011101_00110100_1;
      patterns[22496] = 25'b01010111_11011110_00110101_1;
      patterns[22497] = 25'b01010111_11011111_00110110_1;
      patterns[22498] = 25'b01010111_11100000_00110111_1;
      patterns[22499] = 25'b01010111_11100001_00111000_1;
      patterns[22500] = 25'b01010111_11100010_00111001_1;
      patterns[22501] = 25'b01010111_11100011_00111010_1;
      patterns[22502] = 25'b01010111_11100100_00111011_1;
      patterns[22503] = 25'b01010111_11100101_00111100_1;
      patterns[22504] = 25'b01010111_11100110_00111101_1;
      patterns[22505] = 25'b01010111_11100111_00111110_1;
      patterns[22506] = 25'b01010111_11101000_00111111_1;
      patterns[22507] = 25'b01010111_11101001_01000000_1;
      patterns[22508] = 25'b01010111_11101010_01000001_1;
      patterns[22509] = 25'b01010111_11101011_01000010_1;
      patterns[22510] = 25'b01010111_11101100_01000011_1;
      patterns[22511] = 25'b01010111_11101101_01000100_1;
      patterns[22512] = 25'b01010111_11101110_01000101_1;
      patterns[22513] = 25'b01010111_11101111_01000110_1;
      patterns[22514] = 25'b01010111_11110000_01000111_1;
      patterns[22515] = 25'b01010111_11110001_01001000_1;
      patterns[22516] = 25'b01010111_11110010_01001001_1;
      patterns[22517] = 25'b01010111_11110011_01001010_1;
      patterns[22518] = 25'b01010111_11110100_01001011_1;
      patterns[22519] = 25'b01010111_11110101_01001100_1;
      patterns[22520] = 25'b01010111_11110110_01001101_1;
      patterns[22521] = 25'b01010111_11110111_01001110_1;
      patterns[22522] = 25'b01010111_11111000_01001111_1;
      patterns[22523] = 25'b01010111_11111001_01010000_1;
      patterns[22524] = 25'b01010111_11111010_01010001_1;
      patterns[22525] = 25'b01010111_11111011_01010010_1;
      patterns[22526] = 25'b01010111_11111100_01010011_1;
      patterns[22527] = 25'b01010111_11111101_01010100_1;
      patterns[22528] = 25'b01010111_11111110_01010101_1;
      patterns[22529] = 25'b01010111_11111111_01010110_1;
      patterns[22530] = 25'b01011000_00000000_01011000_0;
      patterns[22531] = 25'b01011000_00000001_01011001_0;
      patterns[22532] = 25'b01011000_00000010_01011010_0;
      patterns[22533] = 25'b01011000_00000011_01011011_0;
      patterns[22534] = 25'b01011000_00000100_01011100_0;
      patterns[22535] = 25'b01011000_00000101_01011101_0;
      patterns[22536] = 25'b01011000_00000110_01011110_0;
      patterns[22537] = 25'b01011000_00000111_01011111_0;
      patterns[22538] = 25'b01011000_00001000_01100000_0;
      patterns[22539] = 25'b01011000_00001001_01100001_0;
      patterns[22540] = 25'b01011000_00001010_01100010_0;
      patterns[22541] = 25'b01011000_00001011_01100011_0;
      patterns[22542] = 25'b01011000_00001100_01100100_0;
      patterns[22543] = 25'b01011000_00001101_01100101_0;
      patterns[22544] = 25'b01011000_00001110_01100110_0;
      patterns[22545] = 25'b01011000_00001111_01100111_0;
      patterns[22546] = 25'b01011000_00010000_01101000_0;
      patterns[22547] = 25'b01011000_00010001_01101001_0;
      patterns[22548] = 25'b01011000_00010010_01101010_0;
      patterns[22549] = 25'b01011000_00010011_01101011_0;
      patterns[22550] = 25'b01011000_00010100_01101100_0;
      patterns[22551] = 25'b01011000_00010101_01101101_0;
      patterns[22552] = 25'b01011000_00010110_01101110_0;
      patterns[22553] = 25'b01011000_00010111_01101111_0;
      patterns[22554] = 25'b01011000_00011000_01110000_0;
      patterns[22555] = 25'b01011000_00011001_01110001_0;
      patterns[22556] = 25'b01011000_00011010_01110010_0;
      patterns[22557] = 25'b01011000_00011011_01110011_0;
      patterns[22558] = 25'b01011000_00011100_01110100_0;
      patterns[22559] = 25'b01011000_00011101_01110101_0;
      patterns[22560] = 25'b01011000_00011110_01110110_0;
      patterns[22561] = 25'b01011000_00011111_01110111_0;
      patterns[22562] = 25'b01011000_00100000_01111000_0;
      patterns[22563] = 25'b01011000_00100001_01111001_0;
      patterns[22564] = 25'b01011000_00100010_01111010_0;
      patterns[22565] = 25'b01011000_00100011_01111011_0;
      patterns[22566] = 25'b01011000_00100100_01111100_0;
      patterns[22567] = 25'b01011000_00100101_01111101_0;
      patterns[22568] = 25'b01011000_00100110_01111110_0;
      patterns[22569] = 25'b01011000_00100111_01111111_0;
      patterns[22570] = 25'b01011000_00101000_10000000_0;
      patterns[22571] = 25'b01011000_00101001_10000001_0;
      patterns[22572] = 25'b01011000_00101010_10000010_0;
      patterns[22573] = 25'b01011000_00101011_10000011_0;
      patterns[22574] = 25'b01011000_00101100_10000100_0;
      patterns[22575] = 25'b01011000_00101101_10000101_0;
      patterns[22576] = 25'b01011000_00101110_10000110_0;
      patterns[22577] = 25'b01011000_00101111_10000111_0;
      patterns[22578] = 25'b01011000_00110000_10001000_0;
      patterns[22579] = 25'b01011000_00110001_10001001_0;
      patterns[22580] = 25'b01011000_00110010_10001010_0;
      patterns[22581] = 25'b01011000_00110011_10001011_0;
      patterns[22582] = 25'b01011000_00110100_10001100_0;
      patterns[22583] = 25'b01011000_00110101_10001101_0;
      patterns[22584] = 25'b01011000_00110110_10001110_0;
      patterns[22585] = 25'b01011000_00110111_10001111_0;
      patterns[22586] = 25'b01011000_00111000_10010000_0;
      patterns[22587] = 25'b01011000_00111001_10010001_0;
      patterns[22588] = 25'b01011000_00111010_10010010_0;
      patterns[22589] = 25'b01011000_00111011_10010011_0;
      patterns[22590] = 25'b01011000_00111100_10010100_0;
      patterns[22591] = 25'b01011000_00111101_10010101_0;
      patterns[22592] = 25'b01011000_00111110_10010110_0;
      patterns[22593] = 25'b01011000_00111111_10010111_0;
      patterns[22594] = 25'b01011000_01000000_10011000_0;
      patterns[22595] = 25'b01011000_01000001_10011001_0;
      patterns[22596] = 25'b01011000_01000010_10011010_0;
      patterns[22597] = 25'b01011000_01000011_10011011_0;
      patterns[22598] = 25'b01011000_01000100_10011100_0;
      patterns[22599] = 25'b01011000_01000101_10011101_0;
      patterns[22600] = 25'b01011000_01000110_10011110_0;
      patterns[22601] = 25'b01011000_01000111_10011111_0;
      patterns[22602] = 25'b01011000_01001000_10100000_0;
      patterns[22603] = 25'b01011000_01001001_10100001_0;
      patterns[22604] = 25'b01011000_01001010_10100010_0;
      patterns[22605] = 25'b01011000_01001011_10100011_0;
      patterns[22606] = 25'b01011000_01001100_10100100_0;
      patterns[22607] = 25'b01011000_01001101_10100101_0;
      patterns[22608] = 25'b01011000_01001110_10100110_0;
      patterns[22609] = 25'b01011000_01001111_10100111_0;
      patterns[22610] = 25'b01011000_01010000_10101000_0;
      patterns[22611] = 25'b01011000_01010001_10101001_0;
      patterns[22612] = 25'b01011000_01010010_10101010_0;
      patterns[22613] = 25'b01011000_01010011_10101011_0;
      patterns[22614] = 25'b01011000_01010100_10101100_0;
      patterns[22615] = 25'b01011000_01010101_10101101_0;
      patterns[22616] = 25'b01011000_01010110_10101110_0;
      patterns[22617] = 25'b01011000_01010111_10101111_0;
      patterns[22618] = 25'b01011000_01011000_10110000_0;
      patterns[22619] = 25'b01011000_01011001_10110001_0;
      patterns[22620] = 25'b01011000_01011010_10110010_0;
      patterns[22621] = 25'b01011000_01011011_10110011_0;
      patterns[22622] = 25'b01011000_01011100_10110100_0;
      patterns[22623] = 25'b01011000_01011101_10110101_0;
      patterns[22624] = 25'b01011000_01011110_10110110_0;
      patterns[22625] = 25'b01011000_01011111_10110111_0;
      patterns[22626] = 25'b01011000_01100000_10111000_0;
      patterns[22627] = 25'b01011000_01100001_10111001_0;
      patterns[22628] = 25'b01011000_01100010_10111010_0;
      patterns[22629] = 25'b01011000_01100011_10111011_0;
      patterns[22630] = 25'b01011000_01100100_10111100_0;
      patterns[22631] = 25'b01011000_01100101_10111101_0;
      patterns[22632] = 25'b01011000_01100110_10111110_0;
      patterns[22633] = 25'b01011000_01100111_10111111_0;
      patterns[22634] = 25'b01011000_01101000_11000000_0;
      patterns[22635] = 25'b01011000_01101001_11000001_0;
      patterns[22636] = 25'b01011000_01101010_11000010_0;
      patterns[22637] = 25'b01011000_01101011_11000011_0;
      patterns[22638] = 25'b01011000_01101100_11000100_0;
      patterns[22639] = 25'b01011000_01101101_11000101_0;
      patterns[22640] = 25'b01011000_01101110_11000110_0;
      patterns[22641] = 25'b01011000_01101111_11000111_0;
      patterns[22642] = 25'b01011000_01110000_11001000_0;
      patterns[22643] = 25'b01011000_01110001_11001001_0;
      patterns[22644] = 25'b01011000_01110010_11001010_0;
      patterns[22645] = 25'b01011000_01110011_11001011_0;
      patterns[22646] = 25'b01011000_01110100_11001100_0;
      patterns[22647] = 25'b01011000_01110101_11001101_0;
      patterns[22648] = 25'b01011000_01110110_11001110_0;
      patterns[22649] = 25'b01011000_01110111_11001111_0;
      patterns[22650] = 25'b01011000_01111000_11010000_0;
      patterns[22651] = 25'b01011000_01111001_11010001_0;
      patterns[22652] = 25'b01011000_01111010_11010010_0;
      patterns[22653] = 25'b01011000_01111011_11010011_0;
      patterns[22654] = 25'b01011000_01111100_11010100_0;
      patterns[22655] = 25'b01011000_01111101_11010101_0;
      patterns[22656] = 25'b01011000_01111110_11010110_0;
      patterns[22657] = 25'b01011000_01111111_11010111_0;
      patterns[22658] = 25'b01011000_10000000_11011000_0;
      patterns[22659] = 25'b01011000_10000001_11011001_0;
      patterns[22660] = 25'b01011000_10000010_11011010_0;
      patterns[22661] = 25'b01011000_10000011_11011011_0;
      patterns[22662] = 25'b01011000_10000100_11011100_0;
      patterns[22663] = 25'b01011000_10000101_11011101_0;
      patterns[22664] = 25'b01011000_10000110_11011110_0;
      patterns[22665] = 25'b01011000_10000111_11011111_0;
      patterns[22666] = 25'b01011000_10001000_11100000_0;
      patterns[22667] = 25'b01011000_10001001_11100001_0;
      patterns[22668] = 25'b01011000_10001010_11100010_0;
      patterns[22669] = 25'b01011000_10001011_11100011_0;
      patterns[22670] = 25'b01011000_10001100_11100100_0;
      patterns[22671] = 25'b01011000_10001101_11100101_0;
      patterns[22672] = 25'b01011000_10001110_11100110_0;
      patterns[22673] = 25'b01011000_10001111_11100111_0;
      patterns[22674] = 25'b01011000_10010000_11101000_0;
      patterns[22675] = 25'b01011000_10010001_11101001_0;
      patterns[22676] = 25'b01011000_10010010_11101010_0;
      patterns[22677] = 25'b01011000_10010011_11101011_0;
      patterns[22678] = 25'b01011000_10010100_11101100_0;
      patterns[22679] = 25'b01011000_10010101_11101101_0;
      patterns[22680] = 25'b01011000_10010110_11101110_0;
      patterns[22681] = 25'b01011000_10010111_11101111_0;
      patterns[22682] = 25'b01011000_10011000_11110000_0;
      patterns[22683] = 25'b01011000_10011001_11110001_0;
      patterns[22684] = 25'b01011000_10011010_11110010_0;
      patterns[22685] = 25'b01011000_10011011_11110011_0;
      patterns[22686] = 25'b01011000_10011100_11110100_0;
      patterns[22687] = 25'b01011000_10011101_11110101_0;
      patterns[22688] = 25'b01011000_10011110_11110110_0;
      patterns[22689] = 25'b01011000_10011111_11110111_0;
      patterns[22690] = 25'b01011000_10100000_11111000_0;
      patterns[22691] = 25'b01011000_10100001_11111001_0;
      patterns[22692] = 25'b01011000_10100010_11111010_0;
      patterns[22693] = 25'b01011000_10100011_11111011_0;
      patterns[22694] = 25'b01011000_10100100_11111100_0;
      patterns[22695] = 25'b01011000_10100101_11111101_0;
      patterns[22696] = 25'b01011000_10100110_11111110_0;
      patterns[22697] = 25'b01011000_10100111_11111111_0;
      patterns[22698] = 25'b01011000_10101000_00000000_1;
      patterns[22699] = 25'b01011000_10101001_00000001_1;
      patterns[22700] = 25'b01011000_10101010_00000010_1;
      patterns[22701] = 25'b01011000_10101011_00000011_1;
      patterns[22702] = 25'b01011000_10101100_00000100_1;
      patterns[22703] = 25'b01011000_10101101_00000101_1;
      patterns[22704] = 25'b01011000_10101110_00000110_1;
      patterns[22705] = 25'b01011000_10101111_00000111_1;
      patterns[22706] = 25'b01011000_10110000_00001000_1;
      patterns[22707] = 25'b01011000_10110001_00001001_1;
      patterns[22708] = 25'b01011000_10110010_00001010_1;
      patterns[22709] = 25'b01011000_10110011_00001011_1;
      patterns[22710] = 25'b01011000_10110100_00001100_1;
      patterns[22711] = 25'b01011000_10110101_00001101_1;
      patterns[22712] = 25'b01011000_10110110_00001110_1;
      patterns[22713] = 25'b01011000_10110111_00001111_1;
      patterns[22714] = 25'b01011000_10111000_00010000_1;
      patterns[22715] = 25'b01011000_10111001_00010001_1;
      patterns[22716] = 25'b01011000_10111010_00010010_1;
      patterns[22717] = 25'b01011000_10111011_00010011_1;
      patterns[22718] = 25'b01011000_10111100_00010100_1;
      patterns[22719] = 25'b01011000_10111101_00010101_1;
      patterns[22720] = 25'b01011000_10111110_00010110_1;
      patterns[22721] = 25'b01011000_10111111_00010111_1;
      patterns[22722] = 25'b01011000_11000000_00011000_1;
      patterns[22723] = 25'b01011000_11000001_00011001_1;
      patterns[22724] = 25'b01011000_11000010_00011010_1;
      patterns[22725] = 25'b01011000_11000011_00011011_1;
      patterns[22726] = 25'b01011000_11000100_00011100_1;
      patterns[22727] = 25'b01011000_11000101_00011101_1;
      patterns[22728] = 25'b01011000_11000110_00011110_1;
      patterns[22729] = 25'b01011000_11000111_00011111_1;
      patterns[22730] = 25'b01011000_11001000_00100000_1;
      patterns[22731] = 25'b01011000_11001001_00100001_1;
      patterns[22732] = 25'b01011000_11001010_00100010_1;
      patterns[22733] = 25'b01011000_11001011_00100011_1;
      patterns[22734] = 25'b01011000_11001100_00100100_1;
      patterns[22735] = 25'b01011000_11001101_00100101_1;
      patterns[22736] = 25'b01011000_11001110_00100110_1;
      patterns[22737] = 25'b01011000_11001111_00100111_1;
      patterns[22738] = 25'b01011000_11010000_00101000_1;
      patterns[22739] = 25'b01011000_11010001_00101001_1;
      patterns[22740] = 25'b01011000_11010010_00101010_1;
      patterns[22741] = 25'b01011000_11010011_00101011_1;
      patterns[22742] = 25'b01011000_11010100_00101100_1;
      patterns[22743] = 25'b01011000_11010101_00101101_1;
      patterns[22744] = 25'b01011000_11010110_00101110_1;
      patterns[22745] = 25'b01011000_11010111_00101111_1;
      patterns[22746] = 25'b01011000_11011000_00110000_1;
      patterns[22747] = 25'b01011000_11011001_00110001_1;
      patterns[22748] = 25'b01011000_11011010_00110010_1;
      patterns[22749] = 25'b01011000_11011011_00110011_1;
      patterns[22750] = 25'b01011000_11011100_00110100_1;
      patterns[22751] = 25'b01011000_11011101_00110101_1;
      patterns[22752] = 25'b01011000_11011110_00110110_1;
      patterns[22753] = 25'b01011000_11011111_00110111_1;
      patterns[22754] = 25'b01011000_11100000_00111000_1;
      patterns[22755] = 25'b01011000_11100001_00111001_1;
      patterns[22756] = 25'b01011000_11100010_00111010_1;
      patterns[22757] = 25'b01011000_11100011_00111011_1;
      patterns[22758] = 25'b01011000_11100100_00111100_1;
      patterns[22759] = 25'b01011000_11100101_00111101_1;
      patterns[22760] = 25'b01011000_11100110_00111110_1;
      patterns[22761] = 25'b01011000_11100111_00111111_1;
      patterns[22762] = 25'b01011000_11101000_01000000_1;
      patterns[22763] = 25'b01011000_11101001_01000001_1;
      patterns[22764] = 25'b01011000_11101010_01000010_1;
      patterns[22765] = 25'b01011000_11101011_01000011_1;
      patterns[22766] = 25'b01011000_11101100_01000100_1;
      patterns[22767] = 25'b01011000_11101101_01000101_1;
      patterns[22768] = 25'b01011000_11101110_01000110_1;
      patterns[22769] = 25'b01011000_11101111_01000111_1;
      patterns[22770] = 25'b01011000_11110000_01001000_1;
      patterns[22771] = 25'b01011000_11110001_01001001_1;
      patterns[22772] = 25'b01011000_11110010_01001010_1;
      patterns[22773] = 25'b01011000_11110011_01001011_1;
      patterns[22774] = 25'b01011000_11110100_01001100_1;
      patterns[22775] = 25'b01011000_11110101_01001101_1;
      patterns[22776] = 25'b01011000_11110110_01001110_1;
      patterns[22777] = 25'b01011000_11110111_01001111_1;
      patterns[22778] = 25'b01011000_11111000_01010000_1;
      patterns[22779] = 25'b01011000_11111001_01010001_1;
      patterns[22780] = 25'b01011000_11111010_01010010_1;
      patterns[22781] = 25'b01011000_11111011_01010011_1;
      patterns[22782] = 25'b01011000_11111100_01010100_1;
      patterns[22783] = 25'b01011000_11111101_01010101_1;
      patterns[22784] = 25'b01011000_11111110_01010110_1;
      patterns[22785] = 25'b01011000_11111111_01010111_1;
      patterns[22786] = 25'b01011001_00000000_01011001_0;
      patterns[22787] = 25'b01011001_00000001_01011010_0;
      patterns[22788] = 25'b01011001_00000010_01011011_0;
      patterns[22789] = 25'b01011001_00000011_01011100_0;
      patterns[22790] = 25'b01011001_00000100_01011101_0;
      patterns[22791] = 25'b01011001_00000101_01011110_0;
      patterns[22792] = 25'b01011001_00000110_01011111_0;
      patterns[22793] = 25'b01011001_00000111_01100000_0;
      patterns[22794] = 25'b01011001_00001000_01100001_0;
      patterns[22795] = 25'b01011001_00001001_01100010_0;
      patterns[22796] = 25'b01011001_00001010_01100011_0;
      patterns[22797] = 25'b01011001_00001011_01100100_0;
      patterns[22798] = 25'b01011001_00001100_01100101_0;
      patterns[22799] = 25'b01011001_00001101_01100110_0;
      patterns[22800] = 25'b01011001_00001110_01100111_0;
      patterns[22801] = 25'b01011001_00001111_01101000_0;
      patterns[22802] = 25'b01011001_00010000_01101001_0;
      patterns[22803] = 25'b01011001_00010001_01101010_0;
      patterns[22804] = 25'b01011001_00010010_01101011_0;
      patterns[22805] = 25'b01011001_00010011_01101100_0;
      patterns[22806] = 25'b01011001_00010100_01101101_0;
      patterns[22807] = 25'b01011001_00010101_01101110_0;
      patterns[22808] = 25'b01011001_00010110_01101111_0;
      patterns[22809] = 25'b01011001_00010111_01110000_0;
      patterns[22810] = 25'b01011001_00011000_01110001_0;
      patterns[22811] = 25'b01011001_00011001_01110010_0;
      patterns[22812] = 25'b01011001_00011010_01110011_0;
      patterns[22813] = 25'b01011001_00011011_01110100_0;
      patterns[22814] = 25'b01011001_00011100_01110101_0;
      patterns[22815] = 25'b01011001_00011101_01110110_0;
      patterns[22816] = 25'b01011001_00011110_01110111_0;
      patterns[22817] = 25'b01011001_00011111_01111000_0;
      patterns[22818] = 25'b01011001_00100000_01111001_0;
      patterns[22819] = 25'b01011001_00100001_01111010_0;
      patterns[22820] = 25'b01011001_00100010_01111011_0;
      patterns[22821] = 25'b01011001_00100011_01111100_0;
      patterns[22822] = 25'b01011001_00100100_01111101_0;
      patterns[22823] = 25'b01011001_00100101_01111110_0;
      patterns[22824] = 25'b01011001_00100110_01111111_0;
      patterns[22825] = 25'b01011001_00100111_10000000_0;
      patterns[22826] = 25'b01011001_00101000_10000001_0;
      patterns[22827] = 25'b01011001_00101001_10000010_0;
      patterns[22828] = 25'b01011001_00101010_10000011_0;
      patterns[22829] = 25'b01011001_00101011_10000100_0;
      patterns[22830] = 25'b01011001_00101100_10000101_0;
      patterns[22831] = 25'b01011001_00101101_10000110_0;
      patterns[22832] = 25'b01011001_00101110_10000111_0;
      patterns[22833] = 25'b01011001_00101111_10001000_0;
      patterns[22834] = 25'b01011001_00110000_10001001_0;
      patterns[22835] = 25'b01011001_00110001_10001010_0;
      patterns[22836] = 25'b01011001_00110010_10001011_0;
      patterns[22837] = 25'b01011001_00110011_10001100_0;
      patterns[22838] = 25'b01011001_00110100_10001101_0;
      patterns[22839] = 25'b01011001_00110101_10001110_0;
      patterns[22840] = 25'b01011001_00110110_10001111_0;
      patterns[22841] = 25'b01011001_00110111_10010000_0;
      patterns[22842] = 25'b01011001_00111000_10010001_0;
      patterns[22843] = 25'b01011001_00111001_10010010_0;
      patterns[22844] = 25'b01011001_00111010_10010011_0;
      patterns[22845] = 25'b01011001_00111011_10010100_0;
      patterns[22846] = 25'b01011001_00111100_10010101_0;
      patterns[22847] = 25'b01011001_00111101_10010110_0;
      patterns[22848] = 25'b01011001_00111110_10010111_0;
      patterns[22849] = 25'b01011001_00111111_10011000_0;
      patterns[22850] = 25'b01011001_01000000_10011001_0;
      patterns[22851] = 25'b01011001_01000001_10011010_0;
      patterns[22852] = 25'b01011001_01000010_10011011_0;
      patterns[22853] = 25'b01011001_01000011_10011100_0;
      patterns[22854] = 25'b01011001_01000100_10011101_0;
      patterns[22855] = 25'b01011001_01000101_10011110_0;
      patterns[22856] = 25'b01011001_01000110_10011111_0;
      patterns[22857] = 25'b01011001_01000111_10100000_0;
      patterns[22858] = 25'b01011001_01001000_10100001_0;
      patterns[22859] = 25'b01011001_01001001_10100010_0;
      patterns[22860] = 25'b01011001_01001010_10100011_0;
      patterns[22861] = 25'b01011001_01001011_10100100_0;
      patterns[22862] = 25'b01011001_01001100_10100101_0;
      patterns[22863] = 25'b01011001_01001101_10100110_0;
      patterns[22864] = 25'b01011001_01001110_10100111_0;
      patterns[22865] = 25'b01011001_01001111_10101000_0;
      patterns[22866] = 25'b01011001_01010000_10101001_0;
      patterns[22867] = 25'b01011001_01010001_10101010_0;
      patterns[22868] = 25'b01011001_01010010_10101011_0;
      patterns[22869] = 25'b01011001_01010011_10101100_0;
      patterns[22870] = 25'b01011001_01010100_10101101_0;
      patterns[22871] = 25'b01011001_01010101_10101110_0;
      patterns[22872] = 25'b01011001_01010110_10101111_0;
      patterns[22873] = 25'b01011001_01010111_10110000_0;
      patterns[22874] = 25'b01011001_01011000_10110001_0;
      patterns[22875] = 25'b01011001_01011001_10110010_0;
      patterns[22876] = 25'b01011001_01011010_10110011_0;
      patterns[22877] = 25'b01011001_01011011_10110100_0;
      patterns[22878] = 25'b01011001_01011100_10110101_0;
      patterns[22879] = 25'b01011001_01011101_10110110_0;
      patterns[22880] = 25'b01011001_01011110_10110111_0;
      patterns[22881] = 25'b01011001_01011111_10111000_0;
      patterns[22882] = 25'b01011001_01100000_10111001_0;
      patterns[22883] = 25'b01011001_01100001_10111010_0;
      patterns[22884] = 25'b01011001_01100010_10111011_0;
      patterns[22885] = 25'b01011001_01100011_10111100_0;
      patterns[22886] = 25'b01011001_01100100_10111101_0;
      patterns[22887] = 25'b01011001_01100101_10111110_0;
      patterns[22888] = 25'b01011001_01100110_10111111_0;
      patterns[22889] = 25'b01011001_01100111_11000000_0;
      patterns[22890] = 25'b01011001_01101000_11000001_0;
      patterns[22891] = 25'b01011001_01101001_11000010_0;
      patterns[22892] = 25'b01011001_01101010_11000011_0;
      patterns[22893] = 25'b01011001_01101011_11000100_0;
      patterns[22894] = 25'b01011001_01101100_11000101_0;
      patterns[22895] = 25'b01011001_01101101_11000110_0;
      patterns[22896] = 25'b01011001_01101110_11000111_0;
      patterns[22897] = 25'b01011001_01101111_11001000_0;
      patterns[22898] = 25'b01011001_01110000_11001001_0;
      patterns[22899] = 25'b01011001_01110001_11001010_0;
      patterns[22900] = 25'b01011001_01110010_11001011_0;
      patterns[22901] = 25'b01011001_01110011_11001100_0;
      patterns[22902] = 25'b01011001_01110100_11001101_0;
      patterns[22903] = 25'b01011001_01110101_11001110_0;
      patterns[22904] = 25'b01011001_01110110_11001111_0;
      patterns[22905] = 25'b01011001_01110111_11010000_0;
      patterns[22906] = 25'b01011001_01111000_11010001_0;
      patterns[22907] = 25'b01011001_01111001_11010010_0;
      patterns[22908] = 25'b01011001_01111010_11010011_0;
      patterns[22909] = 25'b01011001_01111011_11010100_0;
      patterns[22910] = 25'b01011001_01111100_11010101_0;
      patterns[22911] = 25'b01011001_01111101_11010110_0;
      patterns[22912] = 25'b01011001_01111110_11010111_0;
      patterns[22913] = 25'b01011001_01111111_11011000_0;
      patterns[22914] = 25'b01011001_10000000_11011001_0;
      patterns[22915] = 25'b01011001_10000001_11011010_0;
      patterns[22916] = 25'b01011001_10000010_11011011_0;
      patterns[22917] = 25'b01011001_10000011_11011100_0;
      patterns[22918] = 25'b01011001_10000100_11011101_0;
      patterns[22919] = 25'b01011001_10000101_11011110_0;
      patterns[22920] = 25'b01011001_10000110_11011111_0;
      patterns[22921] = 25'b01011001_10000111_11100000_0;
      patterns[22922] = 25'b01011001_10001000_11100001_0;
      patterns[22923] = 25'b01011001_10001001_11100010_0;
      patterns[22924] = 25'b01011001_10001010_11100011_0;
      patterns[22925] = 25'b01011001_10001011_11100100_0;
      patterns[22926] = 25'b01011001_10001100_11100101_0;
      patterns[22927] = 25'b01011001_10001101_11100110_0;
      patterns[22928] = 25'b01011001_10001110_11100111_0;
      patterns[22929] = 25'b01011001_10001111_11101000_0;
      patterns[22930] = 25'b01011001_10010000_11101001_0;
      patterns[22931] = 25'b01011001_10010001_11101010_0;
      patterns[22932] = 25'b01011001_10010010_11101011_0;
      patterns[22933] = 25'b01011001_10010011_11101100_0;
      patterns[22934] = 25'b01011001_10010100_11101101_0;
      patterns[22935] = 25'b01011001_10010101_11101110_0;
      patterns[22936] = 25'b01011001_10010110_11101111_0;
      patterns[22937] = 25'b01011001_10010111_11110000_0;
      patterns[22938] = 25'b01011001_10011000_11110001_0;
      patterns[22939] = 25'b01011001_10011001_11110010_0;
      patterns[22940] = 25'b01011001_10011010_11110011_0;
      patterns[22941] = 25'b01011001_10011011_11110100_0;
      patterns[22942] = 25'b01011001_10011100_11110101_0;
      patterns[22943] = 25'b01011001_10011101_11110110_0;
      patterns[22944] = 25'b01011001_10011110_11110111_0;
      patterns[22945] = 25'b01011001_10011111_11111000_0;
      patterns[22946] = 25'b01011001_10100000_11111001_0;
      patterns[22947] = 25'b01011001_10100001_11111010_0;
      patterns[22948] = 25'b01011001_10100010_11111011_0;
      patterns[22949] = 25'b01011001_10100011_11111100_0;
      patterns[22950] = 25'b01011001_10100100_11111101_0;
      patterns[22951] = 25'b01011001_10100101_11111110_0;
      patterns[22952] = 25'b01011001_10100110_11111111_0;
      patterns[22953] = 25'b01011001_10100111_00000000_1;
      patterns[22954] = 25'b01011001_10101000_00000001_1;
      patterns[22955] = 25'b01011001_10101001_00000010_1;
      patterns[22956] = 25'b01011001_10101010_00000011_1;
      patterns[22957] = 25'b01011001_10101011_00000100_1;
      patterns[22958] = 25'b01011001_10101100_00000101_1;
      patterns[22959] = 25'b01011001_10101101_00000110_1;
      patterns[22960] = 25'b01011001_10101110_00000111_1;
      patterns[22961] = 25'b01011001_10101111_00001000_1;
      patterns[22962] = 25'b01011001_10110000_00001001_1;
      patterns[22963] = 25'b01011001_10110001_00001010_1;
      patterns[22964] = 25'b01011001_10110010_00001011_1;
      patterns[22965] = 25'b01011001_10110011_00001100_1;
      patterns[22966] = 25'b01011001_10110100_00001101_1;
      patterns[22967] = 25'b01011001_10110101_00001110_1;
      patterns[22968] = 25'b01011001_10110110_00001111_1;
      patterns[22969] = 25'b01011001_10110111_00010000_1;
      patterns[22970] = 25'b01011001_10111000_00010001_1;
      patterns[22971] = 25'b01011001_10111001_00010010_1;
      patterns[22972] = 25'b01011001_10111010_00010011_1;
      patterns[22973] = 25'b01011001_10111011_00010100_1;
      patterns[22974] = 25'b01011001_10111100_00010101_1;
      patterns[22975] = 25'b01011001_10111101_00010110_1;
      patterns[22976] = 25'b01011001_10111110_00010111_1;
      patterns[22977] = 25'b01011001_10111111_00011000_1;
      patterns[22978] = 25'b01011001_11000000_00011001_1;
      patterns[22979] = 25'b01011001_11000001_00011010_1;
      patterns[22980] = 25'b01011001_11000010_00011011_1;
      patterns[22981] = 25'b01011001_11000011_00011100_1;
      patterns[22982] = 25'b01011001_11000100_00011101_1;
      patterns[22983] = 25'b01011001_11000101_00011110_1;
      patterns[22984] = 25'b01011001_11000110_00011111_1;
      patterns[22985] = 25'b01011001_11000111_00100000_1;
      patterns[22986] = 25'b01011001_11001000_00100001_1;
      patterns[22987] = 25'b01011001_11001001_00100010_1;
      patterns[22988] = 25'b01011001_11001010_00100011_1;
      patterns[22989] = 25'b01011001_11001011_00100100_1;
      patterns[22990] = 25'b01011001_11001100_00100101_1;
      patterns[22991] = 25'b01011001_11001101_00100110_1;
      patterns[22992] = 25'b01011001_11001110_00100111_1;
      patterns[22993] = 25'b01011001_11001111_00101000_1;
      patterns[22994] = 25'b01011001_11010000_00101001_1;
      patterns[22995] = 25'b01011001_11010001_00101010_1;
      patterns[22996] = 25'b01011001_11010010_00101011_1;
      patterns[22997] = 25'b01011001_11010011_00101100_1;
      patterns[22998] = 25'b01011001_11010100_00101101_1;
      patterns[22999] = 25'b01011001_11010101_00101110_1;
      patterns[23000] = 25'b01011001_11010110_00101111_1;
      patterns[23001] = 25'b01011001_11010111_00110000_1;
      patterns[23002] = 25'b01011001_11011000_00110001_1;
      patterns[23003] = 25'b01011001_11011001_00110010_1;
      patterns[23004] = 25'b01011001_11011010_00110011_1;
      patterns[23005] = 25'b01011001_11011011_00110100_1;
      patterns[23006] = 25'b01011001_11011100_00110101_1;
      patterns[23007] = 25'b01011001_11011101_00110110_1;
      patterns[23008] = 25'b01011001_11011110_00110111_1;
      patterns[23009] = 25'b01011001_11011111_00111000_1;
      patterns[23010] = 25'b01011001_11100000_00111001_1;
      patterns[23011] = 25'b01011001_11100001_00111010_1;
      patterns[23012] = 25'b01011001_11100010_00111011_1;
      patterns[23013] = 25'b01011001_11100011_00111100_1;
      patterns[23014] = 25'b01011001_11100100_00111101_1;
      patterns[23015] = 25'b01011001_11100101_00111110_1;
      patterns[23016] = 25'b01011001_11100110_00111111_1;
      patterns[23017] = 25'b01011001_11100111_01000000_1;
      patterns[23018] = 25'b01011001_11101000_01000001_1;
      patterns[23019] = 25'b01011001_11101001_01000010_1;
      patterns[23020] = 25'b01011001_11101010_01000011_1;
      patterns[23021] = 25'b01011001_11101011_01000100_1;
      patterns[23022] = 25'b01011001_11101100_01000101_1;
      patterns[23023] = 25'b01011001_11101101_01000110_1;
      patterns[23024] = 25'b01011001_11101110_01000111_1;
      patterns[23025] = 25'b01011001_11101111_01001000_1;
      patterns[23026] = 25'b01011001_11110000_01001001_1;
      patterns[23027] = 25'b01011001_11110001_01001010_1;
      patterns[23028] = 25'b01011001_11110010_01001011_1;
      patterns[23029] = 25'b01011001_11110011_01001100_1;
      patterns[23030] = 25'b01011001_11110100_01001101_1;
      patterns[23031] = 25'b01011001_11110101_01001110_1;
      patterns[23032] = 25'b01011001_11110110_01001111_1;
      patterns[23033] = 25'b01011001_11110111_01010000_1;
      patterns[23034] = 25'b01011001_11111000_01010001_1;
      patterns[23035] = 25'b01011001_11111001_01010010_1;
      patterns[23036] = 25'b01011001_11111010_01010011_1;
      patterns[23037] = 25'b01011001_11111011_01010100_1;
      patterns[23038] = 25'b01011001_11111100_01010101_1;
      patterns[23039] = 25'b01011001_11111101_01010110_1;
      patterns[23040] = 25'b01011001_11111110_01010111_1;
      patterns[23041] = 25'b01011001_11111111_01011000_1;
      patterns[23042] = 25'b01011010_00000000_01011010_0;
      patterns[23043] = 25'b01011010_00000001_01011011_0;
      patterns[23044] = 25'b01011010_00000010_01011100_0;
      patterns[23045] = 25'b01011010_00000011_01011101_0;
      patterns[23046] = 25'b01011010_00000100_01011110_0;
      patterns[23047] = 25'b01011010_00000101_01011111_0;
      patterns[23048] = 25'b01011010_00000110_01100000_0;
      patterns[23049] = 25'b01011010_00000111_01100001_0;
      patterns[23050] = 25'b01011010_00001000_01100010_0;
      patterns[23051] = 25'b01011010_00001001_01100011_0;
      patterns[23052] = 25'b01011010_00001010_01100100_0;
      patterns[23053] = 25'b01011010_00001011_01100101_0;
      patterns[23054] = 25'b01011010_00001100_01100110_0;
      patterns[23055] = 25'b01011010_00001101_01100111_0;
      patterns[23056] = 25'b01011010_00001110_01101000_0;
      patterns[23057] = 25'b01011010_00001111_01101001_0;
      patterns[23058] = 25'b01011010_00010000_01101010_0;
      patterns[23059] = 25'b01011010_00010001_01101011_0;
      patterns[23060] = 25'b01011010_00010010_01101100_0;
      patterns[23061] = 25'b01011010_00010011_01101101_0;
      patterns[23062] = 25'b01011010_00010100_01101110_0;
      patterns[23063] = 25'b01011010_00010101_01101111_0;
      patterns[23064] = 25'b01011010_00010110_01110000_0;
      patterns[23065] = 25'b01011010_00010111_01110001_0;
      patterns[23066] = 25'b01011010_00011000_01110010_0;
      patterns[23067] = 25'b01011010_00011001_01110011_0;
      patterns[23068] = 25'b01011010_00011010_01110100_0;
      patterns[23069] = 25'b01011010_00011011_01110101_0;
      patterns[23070] = 25'b01011010_00011100_01110110_0;
      patterns[23071] = 25'b01011010_00011101_01110111_0;
      patterns[23072] = 25'b01011010_00011110_01111000_0;
      patterns[23073] = 25'b01011010_00011111_01111001_0;
      patterns[23074] = 25'b01011010_00100000_01111010_0;
      patterns[23075] = 25'b01011010_00100001_01111011_0;
      patterns[23076] = 25'b01011010_00100010_01111100_0;
      patterns[23077] = 25'b01011010_00100011_01111101_0;
      patterns[23078] = 25'b01011010_00100100_01111110_0;
      patterns[23079] = 25'b01011010_00100101_01111111_0;
      patterns[23080] = 25'b01011010_00100110_10000000_0;
      patterns[23081] = 25'b01011010_00100111_10000001_0;
      patterns[23082] = 25'b01011010_00101000_10000010_0;
      patterns[23083] = 25'b01011010_00101001_10000011_0;
      patterns[23084] = 25'b01011010_00101010_10000100_0;
      patterns[23085] = 25'b01011010_00101011_10000101_0;
      patterns[23086] = 25'b01011010_00101100_10000110_0;
      patterns[23087] = 25'b01011010_00101101_10000111_0;
      patterns[23088] = 25'b01011010_00101110_10001000_0;
      patterns[23089] = 25'b01011010_00101111_10001001_0;
      patterns[23090] = 25'b01011010_00110000_10001010_0;
      patterns[23091] = 25'b01011010_00110001_10001011_0;
      patterns[23092] = 25'b01011010_00110010_10001100_0;
      patterns[23093] = 25'b01011010_00110011_10001101_0;
      patterns[23094] = 25'b01011010_00110100_10001110_0;
      patterns[23095] = 25'b01011010_00110101_10001111_0;
      patterns[23096] = 25'b01011010_00110110_10010000_0;
      patterns[23097] = 25'b01011010_00110111_10010001_0;
      patterns[23098] = 25'b01011010_00111000_10010010_0;
      patterns[23099] = 25'b01011010_00111001_10010011_0;
      patterns[23100] = 25'b01011010_00111010_10010100_0;
      patterns[23101] = 25'b01011010_00111011_10010101_0;
      patterns[23102] = 25'b01011010_00111100_10010110_0;
      patterns[23103] = 25'b01011010_00111101_10010111_0;
      patterns[23104] = 25'b01011010_00111110_10011000_0;
      patterns[23105] = 25'b01011010_00111111_10011001_0;
      patterns[23106] = 25'b01011010_01000000_10011010_0;
      patterns[23107] = 25'b01011010_01000001_10011011_0;
      patterns[23108] = 25'b01011010_01000010_10011100_0;
      patterns[23109] = 25'b01011010_01000011_10011101_0;
      patterns[23110] = 25'b01011010_01000100_10011110_0;
      patterns[23111] = 25'b01011010_01000101_10011111_0;
      patterns[23112] = 25'b01011010_01000110_10100000_0;
      patterns[23113] = 25'b01011010_01000111_10100001_0;
      patterns[23114] = 25'b01011010_01001000_10100010_0;
      patterns[23115] = 25'b01011010_01001001_10100011_0;
      patterns[23116] = 25'b01011010_01001010_10100100_0;
      patterns[23117] = 25'b01011010_01001011_10100101_0;
      patterns[23118] = 25'b01011010_01001100_10100110_0;
      patterns[23119] = 25'b01011010_01001101_10100111_0;
      patterns[23120] = 25'b01011010_01001110_10101000_0;
      patterns[23121] = 25'b01011010_01001111_10101001_0;
      patterns[23122] = 25'b01011010_01010000_10101010_0;
      patterns[23123] = 25'b01011010_01010001_10101011_0;
      patterns[23124] = 25'b01011010_01010010_10101100_0;
      patterns[23125] = 25'b01011010_01010011_10101101_0;
      patterns[23126] = 25'b01011010_01010100_10101110_0;
      patterns[23127] = 25'b01011010_01010101_10101111_0;
      patterns[23128] = 25'b01011010_01010110_10110000_0;
      patterns[23129] = 25'b01011010_01010111_10110001_0;
      patterns[23130] = 25'b01011010_01011000_10110010_0;
      patterns[23131] = 25'b01011010_01011001_10110011_0;
      patterns[23132] = 25'b01011010_01011010_10110100_0;
      patterns[23133] = 25'b01011010_01011011_10110101_0;
      patterns[23134] = 25'b01011010_01011100_10110110_0;
      patterns[23135] = 25'b01011010_01011101_10110111_0;
      patterns[23136] = 25'b01011010_01011110_10111000_0;
      patterns[23137] = 25'b01011010_01011111_10111001_0;
      patterns[23138] = 25'b01011010_01100000_10111010_0;
      patterns[23139] = 25'b01011010_01100001_10111011_0;
      patterns[23140] = 25'b01011010_01100010_10111100_0;
      patterns[23141] = 25'b01011010_01100011_10111101_0;
      patterns[23142] = 25'b01011010_01100100_10111110_0;
      patterns[23143] = 25'b01011010_01100101_10111111_0;
      patterns[23144] = 25'b01011010_01100110_11000000_0;
      patterns[23145] = 25'b01011010_01100111_11000001_0;
      patterns[23146] = 25'b01011010_01101000_11000010_0;
      patterns[23147] = 25'b01011010_01101001_11000011_0;
      patterns[23148] = 25'b01011010_01101010_11000100_0;
      patterns[23149] = 25'b01011010_01101011_11000101_0;
      patterns[23150] = 25'b01011010_01101100_11000110_0;
      patterns[23151] = 25'b01011010_01101101_11000111_0;
      patterns[23152] = 25'b01011010_01101110_11001000_0;
      patterns[23153] = 25'b01011010_01101111_11001001_0;
      patterns[23154] = 25'b01011010_01110000_11001010_0;
      patterns[23155] = 25'b01011010_01110001_11001011_0;
      patterns[23156] = 25'b01011010_01110010_11001100_0;
      patterns[23157] = 25'b01011010_01110011_11001101_0;
      patterns[23158] = 25'b01011010_01110100_11001110_0;
      patterns[23159] = 25'b01011010_01110101_11001111_0;
      patterns[23160] = 25'b01011010_01110110_11010000_0;
      patterns[23161] = 25'b01011010_01110111_11010001_0;
      patterns[23162] = 25'b01011010_01111000_11010010_0;
      patterns[23163] = 25'b01011010_01111001_11010011_0;
      patterns[23164] = 25'b01011010_01111010_11010100_0;
      patterns[23165] = 25'b01011010_01111011_11010101_0;
      patterns[23166] = 25'b01011010_01111100_11010110_0;
      patterns[23167] = 25'b01011010_01111101_11010111_0;
      patterns[23168] = 25'b01011010_01111110_11011000_0;
      patterns[23169] = 25'b01011010_01111111_11011001_0;
      patterns[23170] = 25'b01011010_10000000_11011010_0;
      patterns[23171] = 25'b01011010_10000001_11011011_0;
      patterns[23172] = 25'b01011010_10000010_11011100_0;
      patterns[23173] = 25'b01011010_10000011_11011101_0;
      patterns[23174] = 25'b01011010_10000100_11011110_0;
      patterns[23175] = 25'b01011010_10000101_11011111_0;
      patterns[23176] = 25'b01011010_10000110_11100000_0;
      patterns[23177] = 25'b01011010_10000111_11100001_0;
      patterns[23178] = 25'b01011010_10001000_11100010_0;
      patterns[23179] = 25'b01011010_10001001_11100011_0;
      patterns[23180] = 25'b01011010_10001010_11100100_0;
      patterns[23181] = 25'b01011010_10001011_11100101_0;
      patterns[23182] = 25'b01011010_10001100_11100110_0;
      patterns[23183] = 25'b01011010_10001101_11100111_0;
      patterns[23184] = 25'b01011010_10001110_11101000_0;
      patterns[23185] = 25'b01011010_10001111_11101001_0;
      patterns[23186] = 25'b01011010_10010000_11101010_0;
      patterns[23187] = 25'b01011010_10010001_11101011_0;
      patterns[23188] = 25'b01011010_10010010_11101100_0;
      patterns[23189] = 25'b01011010_10010011_11101101_0;
      patterns[23190] = 25'b01011010_10010100_11101110_0;
      patterns[23191] = 25'b01011010_10010101_11101111_0;
      patterns[23192] = 25'b01011010_10010110_11110000_0;
      patterns[23193] = 25'b01011010_10010111_11110001_0;
      patterns[23194] = 25'b01011010_10011000_11110010_0;
      patterns[23195] = 25'b01011010_10011001_11110011_0;
      patterns[23196] = 25'b01011010_10011010_11110100_0;
      patterns[23197] = 25'b01011010_10011011_11110101_0;
      patterns[23198] = 25'b01011010_10011100_11110110_0;
      patterns[23199] = 25'b01011010_10011101_11110111_0;
      patterns[23200] = 25'b01011010_10011110_11111000_0;
      patterns[23201] = 25'b01011010_10011111_11111001_0;
      patterns[23202] = 25'b01011010_10100000_11111010_0;
      patterns[23203] = 25'b01011010_10100001_11111011_0;
      patterns[23204] = 25'b01011010_10100010_11111100_0;
      patterns[23205] = 25'b01011010_10100011_11111101_0;
      patterns[23206] = 25'b01011010_10100100_11111110_0;
      patterns[23207] = 25'b01011010_10100101_11111111_0;
      patterns[23208] = 25'b01011010_10100110_00000000_1;
      patterns[23209] = 25'b01011010_10100111_00000001_1;
      patterns[23210] = 25'b01011010_10101000_00000010_1;
      patterns[23211] = 25'b01011010_10101001_00000011_1;
      patterns[23212] = 25'b01011010_10101010_00000100_1;
      patterns[23213] = 25'b01011010_10101011_00000101_1;
      patterns[23214] = 25'b01011010_10101100_00000110_1;
      patterns[23215] = 25'b01011010_10101101_00000111_1;
      patterns[23216] = 25'b01011010_10101110_00001000_1;
      patterns[23217] = 25'b01011010_10101111_00001001_1;
      patterns[23218] = 25'b01011010_10110000_00001010_1;
      patterns[23219] = 25'b01011010_10110001_00001011_1;
      patterns[23220] = 25'b01011010_10110010_00001100_1;
      patterns[23221] = 25'b01011010_10110011_00001101_1;
      patterns[23222] = 25'b01011010_10110100_00001110_1;
      patterns[23223] = 25'b01011010_10110101_00001111_1;
      patterns[23224] = 25'b01011010_10110110_00010000_1;
      patterns[23225] = 25'b01011010_10110111_00010001_1;
      patterns[23226] = 25'b01011010_10111000_00010010_1;
      patterns[23227] = 25'b01011010_10111001_00010011_1;
      patterns[23228] = 25'b01011010_10111010_00010100_1;
      patterns[23229] = 25'b01011010_10111011_00010101_1;
      patterns[23230] = 25'b01011010_10111100_00010110_1;
      patterns[23231] = 25'b01011010_10111101_00010111_1;
      patterns[23232] = 25'b01011010_10111110_00011000_1;
      patterns[23233] = 25'b01011010_10111111_00011001_1;
      patterns[23234] = 25'b01011010_11000000_00011010_1;
      patterns[23235] = 25'b01011010_11000001_00011011_1;
      patterns[23236] = 25'b01011010_11000010_00011100_1;
      patterns[23237] = 25'b01011010_11000011_00011101_1;
      patterns[23238] = 25'b01011010_11000100_00011110_1;
      patterns[23239] = 25'b01011010_11000101_00011111_1;
      patterns[23240] = 25'b01011010_11000110_00100000_1;
      patterns[23241] = 25'b01011010_11000111_00100001_1;
      patterns[23242] = 25'b01011010_11001000_00100010_1;
      patterns[23243] = 25'b01011010_11001001_00100011_1;
      patterns[23244] = 25'b01011010_11001010_00100100_1;
      patterns[23245] = 25'b01011010_11001011_00100101_1;
      patterns[23246] = 25'b01011010_11001100_00100110_1;
      patterns[23247] = 25'b01011010_11001101_00100111_1;
      patterns[23248] = 25'b01011010_11001110_00101000_1;
      patterns[23249] = 25'b01011010_11001111_00101001_1;
      patterns[23250] = 25'b01011010_11010000_00101010_1;
      patterns[23251] = 25'b01011010_11010001_00101011_1;
      patterns[23252] = 25'b01011010_11010010_00101100_1;
      patterns[23253] = 25'b01011010_11010011_00101101_1;
      patterns[23254] = 25'b01011010_11010100_00101110_1;
      patterns[23255] = 25'b01011010_11010101_00101111_1;
      patterns[23256] = 25'b01011010_11010110_00110000_1;
      patterns[23257] = 25'b01011010_11010111_00110001_1;
      patterns[23258] = 25'b01011010_11011000_00110010_1;
      patterns[23259] = 25'b01011010_11011001_00110011_1;
      patterns[23260] = 25'b01011010_11011010_00110100_1;
      patterns[23261] = 25'b01011010_11011011_00110101_1;
      patterns[23262] = 25'b01011010_11011100_00110110_1;
      patterns[23263] = 25'b01011010_11011101_00110111_1;
      patterns[23264] = 25'b01011010_11011110_00111000_1;
      patterns[23265] = 25'b01011010_11011111_00111001_1;
      patterns[23266] = 25'b01011010_11100000_00111010_1;
      patterns[23267] = 25'b01011010_11100001_00111011_1;
      patterns[23268] = 25'b01011010_11100010_00111100_1;
      patterns[23269] = 25'b01011010_11100011_00111101_1;
      patterns[23270] = 25'b01011010_11100100_00111110_1;
      patterns[23271] = 25'b01011010_11100101_00111111_1;
      patterns[23272] = 25'b01011010_11100110_01000000_1;
      patterns[23273] = 25'b01011010_11100111_01000001_1;
      patterns[23274] = 25'b01011010_11101000_01000010_1;
      patterns[23275] = 25'b01011010_11101001_01000011_1;
      patterns[23276] = 25'b01011010_11101010_01000100_1;
      patterns[23277] = 25'b01011010_11101011_01000101_1;
      patterns[23278] = 25'b01011010_11101100_01000110_1;
      patterns[23279] = 25'b01011010_11101101_01000111_1;
      patterns[23280] = 25'b01011010_11101110_01001000_1;
      patterns[23281] = 25'b01011010_11101111_01001001_1;
      patterns[23282] = 25'b01011010_11110000_01001010_1;
      patterns[23283] = 25'b01011010_11110001_01001011_1;
      patterns[23284] = 25'b01011010_11110010_01001100_1;
      patterns[23285] = 25'b01011010_11110011_01001101_1;
      patterns[23286] = 25'b01011010_11110100_01001110_1;
      patterns[23287] = 25'b01011010_11110101_01001111_1;
      patterns[23288] = 25'b01011010_11110110_01010000_1;
      patterns[23289] = 25'b01011010_11110111_01010001_1;
      patterns[23290] = 25'b01011010_11111000_01010010_1;
      patterns[23291] = 25'b01011010_11111001_01010011_1;
      patterns[23292] = 25'b01011010_11111010_01010100_1;
      patterns[23293] = 25'b01011010_11111011_01010101_1;
      patterns[23294] = 25'b01011010_11111100_01010110_1;
      patterns[23295] = 25'b01011010_11111101_01010111_1;
      patterns[23296] = 25'b01011010_11111110_01011000_1;
      patterns[23297] = 25'b01011010_11111111_01011001_1;
      patterns[23298] = 25'b01011011_00000000_01011011_0;
      patterns[23299] = 25'b01011011_00000001_01011100_0;
      patterns[23300] = 25'b01011011_00000010_01011101_0;
      patterns[23301] = 25'b01011011_00000011_01011110_0;
      patterns[23302] = 25'b01011011_00000100_01011111_0;
      patterns[23303] = 25'b01011011_00000101_01100000_0;
      patterns[23304] = 25'b01011011_00000110_01100001_0;
      patterns[23305] = 25'b01011011_00000111_01100010_0;
      patterns[23306] = 25'b01011011_00001000_01100011_0;
      patterns[23307] = 25'b01011011_00001001_01100100_0;
      patterns[23308] = 25'b01011011_00001010_01100101_0;
      patterns[23309] = 25'b01011011_00001011_01100110_0;
      patterns[23310] = 25'b01011011_00001100_01100111_0;
      patterns[23311] = 25'b01011011_00001101_01101000_0;
      patterns[23312] = 25'b01011011_00001110_01101001_0;
      patterns[23313] = 25'b01011011_00001111_01101010_0;
      patterns[23314] = 25'b01011011_00010000_01101011_0;
      patterns[23315] = 25'b01011011_00010001_01101100_0;
      patterns[23316] = 25'b01011011_00010010_01101101_0;
      patterns[23317] = 25'b01011011_00010011_01101110_0;
      patterns[23318] = 25'b01011011_00010100_01101111_0;
      patterns[23319] = 25'b01011011_00010101_01110000_0;
      patterns[23320] = 25'b01011011_00010110_01110001_0;
      patterns[23321] = 25'b01011011_00010111_01110010_0;
      patterns[23322] = 25'b01011011_00011000_01110011_0;
      patterns[23323] = 25'b01011011_00011001_01110100_0;
      patterns[23324] = 25'b01011011_00011010_01110101_0;
      patterns[23325] = 25'b01011011_00011011_01110110_0;
      patterns[23326] = 25'b01011011_00011100_01110111_0;
      patterns[23327] = 25'b01011011_00011101_01111000_0;
      patterns[23328] = 25'b01011011_00011110_01111001_0;
      patterns[23329] = 25'b01011011_00011111_01111010_0;
      patterns[23330] = 25'b01011011_00100000_01111011_0;
      patterns[23331] = 25'b01011011_00100001_01111100_0;
      patterns[23332] = 25'b01011011_00100010_01111101_0;
      patterns[23333] = 25'b01011011_00100011_01111110_0;
      patterns[23334] = 25'b01011011_00100100_01111111_0;
      patterns[23335] = 25'b01011011_00100101_10000000_0;
      patterns[23336] = 25'b01011011_00100110_10000001_0;
      patterns[23337] = 25'b01011011_00100111_10000010_0;
      patterns[23338] = 25'b01011011_00101000_10000011_0;
      patterns[23339] = 25'b01011011_00101001_10000100_0;
      patterns[23340] = 25'b01011011_00101010_10000101_0;
      patterns[23341] = 25'b01011011_00101011_10000110_0;
      patterns[23342] = 25'b01011011_00101100_10000111_0;
      patterns[23343] = 25'b01011011_00101101_10001000_0;
      patterns[23344] = 25'b01011011_00101110_10001001_0;
      patterns[23345] = 25'b01011011_00101111_10001010_0;
      patterns[23346] = 25'b01011011_00110000_10001011_0;
      patterns[23347] = 25'b01011011_00110001_10001100_0;
      patterns[23348] = 25'b01011011_00110010_10001101_0;
      patterns[23349] = 25'b01011011_00110011_10001110_0;
      patterns[23350] = 25'b01011011_00110100_10001111_0;
      patterns[23351] = 25'b01011011_00110101_10010000_0;
      patterns[23352] = 25'b01011011_00110110_10010001_0;
      patterns[23353] = 25'b01011011_00110111_10010010_0;
      patterns[23354] = 25'b01011011_00111000_10010011_0;
      patterns[23355] = 25'b01011011_00111001_10010100_0;
      patterns[23356] = 25'b01011011_00111010_10010101_0;
      patterns[23357] = 25'b01011011_00111011_10010110_0;
      patterns[23358] = 25'b01011011_00111100_10010111_0;
      patterns[23359] = 25'b01011011_00111101_10011000_0;
      patterns[23360] = 25'b01011011_00111110_10011001_0;
      patterns[23361] = 25'b01011011_00111111_10011010_0;
      patterns[23362] = 25'b01011011_01000000_10011011_0;
      patterns[23363] = 25'b01011011_01000001_10011100_0;
      patterns[23364] = 25'b01011011_01000010_10011101_0;
      patterns[23365] = 25'b01011011_01000011_10011110_0;
      patterns[23366] = 25'b01011011_01000100_10011111_0;
      patterns[23367] = 25'b01011011_01000101_10100000_0;
      patterns[23368] = 25'b01011011_01000110_10100001_0;
      patterns[23369] = 25'b01011011_01000111_10100010_0;
      patterns[23370] = 25'b01011011_01001000_10100011_0;
      patterns[23371] = 25'b01011011_01001001_10100100_0;
      patterns[23372] = 25'b01011011_01001010_10100101_0;
      patterns[23373] = 25'b01011011_01001011_10100110_0;
      patterns[23374] = 25'b01011011_01001100_10100111_0;
      patterns[23375] = 25'b01011011_01001101_10101000_0;
      patterns[23376] = 25'b01011011_01001110_10101001_0;
      patterns[23377] = 25'b01011011_01001111_10101010_0;
      patterns[23378] = 25'b01011011_01010000_10101011_0;
      patterns[23379] = 25'b01011011_01010001_10101100_0;
      patterns[23380] = 25'b01011011_01010010_10101101_0;
      patterns[23381] = 25'b01011011_01010011_10101110_0;
      patterns[23382] = 25'b01011011_01010100_10101111_0;
      patterns[23383] = 25'b01011011_01010101_10110000_0;
      patterns[23384] = 25'b01011011_01010110_10110001_0;
      patterns[23385] = 25'b01011011_01010111_10110010_0;
      patterns[23386] = 25'b01011011_01011000_10110011_0;
      patterns[23387] = 25'b01011011_01011001_10110100_0;
      patterns[23388] = 25'b01011011_01011010_10110101_0;
      patterns[23389] = 25'b01011011_01011011_10110110_0;
      patterns[23390] = 25'b01011011_01011100_10110111_0;
      patterns[23391] = 25'b01011011_01011101_10111000_0;
      patterns[23392] = 25'b01011011_01011110_10111001_0;
      patterns[23393] = 25'b01011011_01011111_10111010_0;
      patterns[23394] = 25'b01011011_01100000_10111011_0;
      patterns[23395] = 25'b01011011_01100001_10111100_0;
      patterns[23396] = 25'b01011011_01100010_10111101_0;
      patterns[23397] = 25'b01011011_01100011_10111110_0;
      patterns[23398] = 25'b01011011_01100100_10111111_0;
      patterns[23399] = 25'b01011011_01100101_11000000_0;
      patterns[23400] = 25'b01011011_01100110_11000001_0;
      patterns[23401] = 25'b01011011_01100111_11000010_0;
      patterns[23402] = 25'b01011011_01101000_11000011_0;
      patterns[23403] = 25'b01011011_01101001_11000100_0;
      patterns[23404] = 25'b01011011_01101010_11000101_0;
      patterns[23405] = 25'b01011011_01101011_11000110_0;
      patterns[23406] = 25'b01011011_01101100_11000111_0;
      patterns[23407] = 25'b01011011_01101101_11001000_0;
      patterns[23408] = 25'b01011011_01101110_11001001_0;
      patterns[23409] = 25'b01011011_01101111_11001010_0;
      patterns[23410] = 25'b01011011_01110000_11001011_0;
      patterns[23411] = 25'b01011011_01110001_11001100_0;
      patterns[23412] = 25'b01011011_01110010_11001101_0;
      patterns[23413] = 25'b01011011_01110011_11001110_0;
      patterns[23414] = 25'b01011011_01110100_11001111_0;
      patterns[23415] = 25'b01011011_01110101_11010000_0;
      patterns[23416] = 25'b01011011_01110110_11010001_0;
      patterns[23417] = 25'b01011011_01110111_11010010_0;
      patterns[23418] = 25'b01011011_01111000_11010011_0;
      patterns[23419] = 25'b01011011_01111001_11010100_0;
      patterns[23420] = 25'b01011011_01111010_11010101_0;
      patterns[23421] = 25'b01011011_01111011_11010110_0;
      patterns[23422] = 25'b01011011_01111100_11010111_0;
      patterns[23423] = 25'b01011011_01111101_11011000_0;
      patterns[23424] = 25'b01011011_01111110_11011001_0;
      patterns[23425] = 25'b01011011_01111111_11011010_0;
      patterns[23426] = 25'b01011011_10000000_11011011_0;
      patterns[23427] = 25'b01011011_10000001_11011100_0;
      patterns[23428] = 25'b01011011_10000010_11011101_0;
      patterns[23429] = 25'b01011011_10000011_11011110_0;
      patterns[23430] = 25'b01011011_10000100_11011111_0;
      patterns[23431] = 25'b01011011_10000101_11100000_0;
      patterns[23432] = 25'b01011011_10000110_11100001_0;
      patterns[23433] = 25'b01011011_10000111_11100010_0;
      patterns[23434] = 25'b01011011_10001000_11100011_0;
      patterns[23435] = 25'b01011011_10001001_11100100_0;
      patterns[23436] = 25'b01011011_10001010_11100101_0;
      patterns[23437] = 25'b01011011_10001011_11100110_0;
      patterns[23438] = 25'b01011011_10001100_11100111_0;
      patterns[23439] = 25'b01011011_10001101_11101000_0;
      patterns[23440] = 25'b01011011_10001110_11101001_0;
      patterns[23441] = 25'b01011011_10001111_11101010_0;
      patterns[23442] = 25'b01011011_10010000_11101011_0;
      patterns[23443] = 25'b01011011_10010001_11101100_0;
      patterns[23444] = 25'b01011011_10010010_11101101_0;
      patterns[23445] = 25'b01011011_10010011_11101110_0;
      patterns[23446] = 25'b01011011_10010100_11101111_0;
      patterns[23447] = 25'b01011011_10010101_11110000_0;
      patterns[23448] = 25'b01011011_10010110_11110001_0;
      patterns[23449] = 25'b01011011_10010111_11110010_0;
      patterns[23450] = 25'b01011011_10011000_11110011_0;
      patterns[23451] = 25'b01011011_10011001_11110100_0;
      patterns[23452] = 25'b01011011_10011010_11110101_0;
      patterns[23453] = 25'b01011011_10011011_11110110_0;
      patterns[23454] = 25'b01011011_10011100_11110111_0;
      patterns[23455] = 25'b01011011_10011101_11111000_0;
      patterns[23456] = 25'b01011011_10011110_11111001_0;
      patterns[23457] = 25'b01011011_10011111_11111010_0;
      patterns[23458] = 25'b01011011_10100000_11111011_0;
      patterns[23459] = 25'b01011011_10100001_11111100_0;
      patterns[23460] = 25'b01011011_10100010_11111101_0;
      patterns[23461] = 25'b01011011_10100011_11111110_0;
      patterns[23462] = 25'b01011011_10100100_11111111_0;
      patterns[23463] = 25'b01011011_10100101_00000000_1;
      patterns[23464] = 25'b01011011_10100110_00000001_1;
      patterns[23465] = 25'b01011011_10100111_00000010_1;
      patterns[23466] = 25'b01011011_10101000_00000011_1;
      patterns[23467] = 25'b01011011_10101001_00000100_1;
      patterns[23468] = 25'b01011011_10101010_00000101_1;
      patterns[23469] = 25'b01011011_10101011_00000110_1;
      patterns[23470] = 25'b01011011_10101100_00000111_1;
      patterns[23471] = 25'b01011011_10101101_00001000_1;
      patterns[23472] = 25'b01011011_10101110_00001001_1;
      patterns[23473] = 25'b01011011_10101111_00001010_1;
      patterns[23474] = 25'b01011011_10110000_00001011_1;
      patterns[23475] = 25'b01011011_10110001_00001100_1;
      patterns[23476] = 25'b01011011_10110010_00001101_1;
      patterns[23477] = 25'b01011011_10110011_00001110_1;
      patterns[23478] = 25'b01011011_10110100_00001111_1;
      patterns[23479] = 25'b01011011_10110101_00010000_1;
      patterns[23480] = 25'b01011011_10110110_00010001_1;
      patterns[23481] = 25'b01011011_10110111_00010010_1;
      patterns[23482] = 25'b01011011_10111000_00010011_1;
      patterns[23483] = 25'b01011011_10111001_00010100_1;
      patterns[23484] = 25'b01011011_10111010_00010101_1;
      patterns[23485] = 25'b01011011_10111011_00010110_1;
      patterns[23486] = 25'b01011011_10111100_00010111_1;
      patterns[23487] = 25'b01011011_10111101_00011000_1;
      patterns[23488] = 25'b01011011_10111110_00011001_1;
      patterns[23489] = 25'b01011011_10111111_00011010_1;
      patterns[23490] = 25'b01011011_11000000_00011011_1;
      patterns[23491] = 25'b01011011_11000001_00011100_1;
      patterns[23492] = 25'b01011011_11000010_00011101_1;
      patterns[23493] = 25'b01011011_11000011_00011110_1;
      patterns[23494] = 25'b01011011_11000100_00011111_1;
      patterns[23495] = 25'b01011011_11000101_00100000_1;
      patterns[23496] = 25'b01011011_11000110_00100001_1;
      patterns[23497] = 25'b01011011_11000111_00100010_1;
      patterns[23498] = 25'b01011011_11001000_00100011_1;
      patterns[23499] = 25'b01011011_11001001_00100100_1;
      patterns[23500] = 25'b01011011_11001010_00100101_1;
      patterns[23501] = 25'b01011011_11001011_00100110_1;
      patterns[23502] = 25'b01011011_11001100_00100111_1;
      patterns[23503] = 25'b01011011_11001101_00101000_1;
      patterns[23504] = 25'b01011011_11001110_00101001_1;
      patterns[23505] = 25'b01011011_11001111_00101010_1;
      patterns[23506] = 25'b01011011_11010000_00101011_1;
      patterns[23507] = 25'b01011011_11010001_00101100_1;
      patterns[23508] = 25'b01011011_11010010_00101101_1;
      patterns[23509] = 25'b01011011_11010011_00101110_1;
      patterns[23510] = 25'b01011011_11010100_00101111_1;
      patterns[23511] = 25'b01011011_11010101_00110000_1;
      patterns[23512] = 25'b01011011_11010110_00110001_1;
      patterns[23513] = 25'b01011011_11010111_00110010_1;
      patterns[23514] = 25'b01011011_11011000_00110011_1;
      patterns[23515] = 25'b01011011_11011001_00110100_1;
      patterns[23516] = 25'b01011011_11011010_00110101_1;
      patterns[23517] = 25'b01011011_11011011_00110110_1;
      patterns[23518] = 25'b01011011_11011100_00110111_1;
      patterns[23519] = 25'b01011011_11011101_00111000_1;
      patterns[23520] = 25'b01011011_11011110_00111001_1;
      patterns[23521] = 25'b01011011_11011111_00111010_1;
      patterns[23522] = 25'b01011011_11100000_00111011_1;
      patterns[23523] = 25'b01011011_11100001_00111100_1;
      patterns[23524] = 25'b01011011_11100010_00111101_1;
      patterns[23525] = 25'b01011011_11100011_00111110_1;
      patterns[23526] = 25'b01011011_11100100_00111111_1;
      patterns[23527] = 25'b01011011_11100101_01000000_1;
      patterns[23528] = 25'b01011011_11100110_01000001_1;
      patterns[23529] = 25'b01011011_11100111_01000010_1;
      patterns[23530] = 25'b01011011_11101000_01000011_1;
      patterns[23531] = 25'b01011011_11101001_01000100_1;
      patterns[23532] = 25'b01011011_11101010_01000101_1;
      patterns[23533] = 25'b01011011_11101011_01000110_1;
      patterns[23534] = 25'b01011011_11101100_01000111_1;
      patterns[23535] = 25'b01011011_11101101_01001000_1;
      patterns[23536] = 25'b01011011_11101110_01001001_1;
      patterns[23537] = 25'b01011011_11101111_01001010_1;
      patterns[23538] = 25'b01011011_11110000_01001011_1;
      patterns[23539] = 25'b01011011_11110001_01001100_1;
      patterns[23540] = 25'b01011011_11110010_01001101_1;
      patterns[23541] = 25'b01011011_11110011_01001110_1;
      patterns[23542] = 25'b01011011_11110100_01001111_1;
      patterns[23543] = 25'b01011011_11110101_01010000_1;
      patterns[23544] = 25'b01011011_11110110_01010001_1;
      patterns[23545] = 25'b01011011_11110111_01010010_1;
      patterns[23546] = 25'b01011011_11111000_01010011_1;
      patterns[23547] = 25'b01011011_11111001_01010100_1;
      patterns[23548] = 25'b01011011_11111010_01010101_1;
      patterns[23549] = 25'b01011011_11111011_01010110_1;
      patterns[23550] = 25'b01011011_11111100_01010111_1;
      patterns[23551] = 25'b01011011_11111101_01011000_1;
      patterns[23552] = 25'b01011011_11111110_01011001_1;
      patterns[23553] = 25'b01011011_11111111_01011010_1;
      patterns[23554] = 25'b01011100_00000000_01011100_0;
      patterns[23555] = 25'b01011100_00000001_01011101_0;
      patterns[23556] = 25'b01011100_00000010_01011110_0;
      patterns[23557] = 25'b01011100_00000011_01011111_0;
      patterns[23558] = 25'b01011100_00000100_01100000_0;
      patterns[23559] = 25'b01011100_00000101_01100001_0;
      patterns[23560] = 25'b01011100_00000110_01100010_0;
      patterns[23561] = 25'b01011100_00000111_01100011_0;
      patterns[23562] = 25'b01011100_00001000_01100100_0;
      patterns[23563] = 25'b01011100_00001001_01100101_0;
      patterns[23564] = 25'b01011100_00001010_01100110_0;
      patterns[23565] = 25'b01011100_00001011_01100111_0;
      patterns[23566] = 25'b01011100_00001100_01101000_0;
      patterns[23567] = 25'b01011100_00001101_01101001_0;
      patterns[23568] = 25'b01011100_00001110_01101010_0;
      patterns[23569] = 25'b01011100_00001111_01101011_0;
      patterns[23570] = 25'b01011100_00010000_01101100_0;
      patterns[23571] = 25'b01011100_00010001_01101101_0;
      patterns[23572] = 25'b01011100_00010010_01101110_0;
      patterns[23573] = 25'b01011100_00010011_01101111_0;
      patterns[23574] = 25'b01011100_00010100_01110000_0;
      patterns[23575] = 25'b01011100_00010101_01110001_0;
      patterns[23576] = 25'b01011100_00010110_01110010_0;
      patterns[23577] = 25'b01011100_00010111_01110011_0;
      patterns[23578] = 25'b01011100_00011000_01110100_0;
      patterns[23579] = 25'b01011100_00011001_01110101_0;
      patterns[23580] = 25'b01011100_00011010_01110110_0;
      patterns[23581] = 25'b01011100_00011011_01110111_0;
      patterns[23582] = 25'b01011100_00011100_01111000_0;
      patterns[23583] = 25'b01011100_00011101_01111001_0;
      patterns[23584] = 25'b01011100_00011110_01111010_0;
      patterns[23585] = 25'b01011100_00011111_01111011_0;
      patterns[23586] = 25'b01011100_00100000_01111100_0;
      patterns[23587] = 25'b01011100_00100001_01111101_0;
      patterns[23588] = 25'b01011100_00100010_01111110_0;
      patterns[23589] = 25'b01011100_00100011_01111111_0;
      patterns[23590] = 25'b01011100_00100100_10000000_0;
      patterns[23591] = 25'b01011100_00100101_10000001_0;
      patterns[23592] = 25'b01011100_00100110_10000010_0;
      patterns[23593] = 25'b01011100_00100111_10000011_0;
      patterns[23594] = 25'b01011100_00101000_10000100_0;
      patterns[23595] = 25'b01011100_00101001_10000101_0;
      patterns[23596] = 25'b01011100_00101010_10000110_0;
      patterns[23597] = 25'b01011100_00101011_10000111_0;
      patterns[23598] = 25'b01011100_00101100_10001000_0;
      patterns[23599] = 25'b01011100_00101101_10001001_0;
      patterns[23600] = 25'b01011100_00101110_10001010_0;
      patterns[23601] = 25'b01011100_00101111_10001011_0;
      patterns[23602] = 25'b01011100_00110000_10001100_0;
      patterns[23603] = 25'b01011100_00110001_10001101_0;
      patterns[23604] = 25'b01011100_00110010_10001110_0;
      patterns[23605] = 25'b01011100_00110011_10001111_0;
      patterns[23606] = 25'b01011100_00110100_10010000_0;
      patterns[23607] = 25'b01011100_00110101_10010001_0;
      patterns[23608] = 25'b01011100_00110110_10010010_0;
      patterns[23609] = 25'b01011100_00110111_10010011_0;
      patterns[23610] = 25'b01011100_00111000_10010100_0;
      patterns[23611] = 25'b01011100_00111001_10010101_0;
      patterns[23612] = 25'b01011100_00111010_10010110_0;
      patterns[23613] = 25'b01011100_00111011_10010111_0;
      patterns[23614] = 25'b01011100_00111100_10011000_0;
      patterns[23615] = 25'b01011100_00111101_10011001_0;
      patterns[23616] = 25'b01011100_00111110_10011010_0;
      patterns[23617] = 25'b01011100_00111111_10011011_0;
      patterns[23618] = 25'b01011100_01000000_10011100_0;
      patterns[23619] = 25'b01011100_01000001_10011101_0;
      patterns[23620] = 25'b01011100_01000010_10011110_0;
      patterns[23621] = 25'b01011100_01000011_10011111_0;
      patterns[23622] = 25'b01011100_01000100_10100000_0;
      patterns[23623] = 25'b01011100_01000101_10100001_0;
      patterns[23624] = 25'b01011100_01000110_10100010_0;
      patterns[23625] = 25'b01011100_01000111_10100011_0;
      patterns[23626] = 25'b01011100_01001000_10100100_0;
      patterns[23627] = 25'b01011100_01001001_10100101_0;
      patterns[23628] = 25'b01011100_01001010_10100110_0;
      patterns[23629] = 25'b01011100_01001011_10100111_0;
      patterns[23630] = 25'b01011100_01001100_10101000_0;
      patterns[23631] = 25'b01011100_01001101_10101001_0;
      patterns[23632] = 25'b01011100_01001110_10101010_0;
      patterns[23633] = 25'b01011100_01001111_10101011_0;
      patterns[23634] = 25'b01011100_01010000_10101100_0;
      patterns[23635] = 25'b01011100_01010001_10101101_0;
      patterns[23636] = 25'b01011100_01010010_10101110_0;
      patterns[23637] = 25'b01011100_01010011_10101111_0;
      patterns[23638] = 25'b01011100_01010100_10110000_0;
      patterns[23639] = 25'b01011100_01010101_10110001_0;
      patterns[23640] = 25'b01011100_01010110_10110010_0;
      patterns[23641] = 25'b01011100_01010111_10110011_0;
      patterns[23642] = 25'b01011100_01011000_10110100_0;
      patterns[23643] = 25'b01011100_01011001_10110101_0;
      patterns[23644] = 25'b01011100_01011010_10110110_0;
      patterns[23645] = 25'b01011100_01011011_10110111_0;
      patterns[23646] = 25'b01011100_01011100_10111000_0;
      patterns[23647] = 25'b01011100_01011101_10111001_0;
      patterns[23648] = 25'b01011100_01011110_10111010_0;
      patterns[23649] = 25'b01011100_01011111_10111011_0;
      patterns[23650] = 25'b01011100_01100000_10111100_0;
      patterns[23651] = 25'b01011100_01100001_10111101_0;
      patterns[23652] = 25'b01011100_01100010_10111110_0;
      patterns[23653] = 25'b01011100_01100011_10111111_0;
      patterns[23654] = 25'b01011100_01100100_11000000_0;
      patterns[23655] = 25'b01011100_01100101_11000001_0;
      patterns[23656] = 25'b01011100_01100110_11000010_0;
      patterns[23657] = 25'b01011100_01100111_11000011_0;
      patterns[23658] = 25'b01011100_01101000_11000100_0;
      patterns[23659] = 25'b01011100_01101001_11000101_0;
      patterns[23660] = 25'b01011100_01101010_11000110_0;
      patterns[23661] = 25'b01011100_01101011_11000111_0;
      patterns[23662] = 25'b01011100_01101100_11001000_0;
      patterns[23663] = 25'b01011100_01101101_11001001_0;
      patterns[23664] = 25'b01011100_01101110_11001010_0;
      patterns[23665] = 25'b01011100_01101111_11001011_0;
      patterns[23666] = 25'b01011100_01110000_11001100_0;
      patterns[23667] = 25'b01011100_01110001_11001101_0;
      patterns[23668] = 25'b01011100_01110010_11001110_0;
      patterns[23669] = 25'b01011100_01110011_11001111_0;
      patterns[23670] = 25'b01011100_01110100_11010000_0;
      patterns[23671] = 25'b01011100_01110101_11010001_0;
      patterns[23672] = 25'b01011100_01110110_11010010_0;
      patterns[23673] = 25'b01011100_01110111_11010011_0;
      patterns[23674] = 25'b01011100_01111000_11010100_0;
      patterns[23675] = 25'b01011100_01111001_11010101_0;
      patterns[23676] = 25'b01011100_01111010_11010110_0;
      patterns[23677] = 25'b01011100_01111011_11010111_0;
      patterns[23678] = 25'b01011100_01111100_11011000_0;
      patterns[23679] = 25'b01011100_01111101_11011001_0;
      patterns[23680] = 25'b01011100_01111110_11011010_0;
      patterns[23681] = 25'b01011100_01111111_11011011_0;
      patterns[23682] = 25'b01011100_10000000_11011100_0;
      patterns[23683] = 25'b01011100_10000001_11011101_0;
      patterns[23684] = 25'b01011100_10000010_11011110_0;
      patterns[23685] = 25'b01011100_10000011_11011111_0;
      patterns[23686] = 25'b01011100_10000100_11100000_0;
      patterns[23687] = 25'b01011100_10000101_11100001_0;
      patterns[23688] = 25'b01011100_10000110_11100010_0;
      patterns[23689] = 25'b01011100_10000111_11100011_0;
      patterns[23690] = 25'b01011100_10001000_11100100_0;
      patterns[23691] = 25'b01011100_10001001_11100101_0;
      patterns[23692] = 25'b01011100_10001010_11100110_0;
      patterns[23693] = 25'b01011100_10001011_11100111_0;
      patterns[23694] = 25'b01011100_10001100_11101000_0;
      patterns[23695] = 25'b01011100_10001101_11101001_0;
      patterns[23696] = 25'b01011100_10001110_11101010_0;
      patterns[23697] = 25'b01011100_10001111_11101011_0;
      patterns[23698] = 25'b01011100_10010000_11101100_0;
      patterns[23699] = 25'b01011100_10010001_11101101_0;
      patterns[23700] = 25'b01011100_10010010_11101110_0;
      patterns[23701] = 25'b01011100_10010011_11101111_0;
      patterns[23702] = 25'b01011100_10010100_11110000_0;
      patterns[23703] = 25'b01011100_10010101_11110001_0;
      patterns[23704] = 25'b01011100_10010110_11110010_0;
      patterns[23705] = 25'b01011100_10010111_11110011_0;
      patterns[23706] = 25'b01011100_10011000_11110100_0;
      patterns[23707] = 25'b01011100_10011001_11110101_0;
      patterns[23708] = 25'b01011100_10011010_11110110_0;
      patterns[23709] = 25'b01011100_10011011_11110111_0;
      patterns[23710] = 25'b01011100_10011100_11111000_0;
      patterns[23711] = 25'b01011100_10011101_11111001_0;
      patterns[23712] = 25'b01011100_10011110_11111010_0;
      patterns[23713] = 25'b01011100_10011111_11111011_0;
      patterns[23714] = 25'b01011100_10100000_11111100_0;
      patterns[23715] = 25'b01011100_10100001_11111101_0;
      patterns[23716] = 25'b01011100_10100010_11111110_0;
      patterns[23717] = 25'b01011100_10100011_11111111_0;
      patterns[23718] = 25'b01011100_10100100_00000000_1;
      patterns[23719] = 25'b01011100_10100101_00000001_1;
      patterns[23720] = 25'b01011100_10100110_00000010_1;
      patterns[23721] = 25'b01011100_10100111_00000011_1;
      patterns[23722] = 25'b01011100_10101000_00000100_1;
      patterns[23723] = 25'b01011100_10101001_00000101_1;
      patterns[23724] = 25'b01011100_10101010_00000110_1;
      patterns[23725] = 25'b01011100_10101011_00000111_1;
      patterns[23726] = 25'b01011100_10101100_00001000_1;
      patterns[23727] = 25'b01011100_10101101_00001001_1;
      patterns[23728] = 25'b01011100_10101110_00001010_1;
      patterns[23729] = 25'b01011100_10101111_00001011_1;
      patterns[23730] = 25'b01011100_10110000_00001100_1;
      patterns[23731] = 25'b01011100_10110001_00001101_1;
      patterns[23732] = 25'b01011100_10110010_00001110_1;
      patterns[23733] = 25'b01011100_10110011_00001111_1;
      patterns[23734] = 25'b01011100_10110100_00010000_1;
      patterns[23735] = 25'b01011100_10110101_00010001_1;
      patterns[23736] = 25'b01011100_10110110_00010010_1;
      patterns[23737] = 25'b01011100_10110111_00010011_1;
      patterns[23738] = 25'b01011100_10111000_00010100_1;
      patterns[23739] = 25'b01011100_10111001_00010101_1;
      patterns[23740] = 25'b01011100_10111010_00010110_1;
      patterns[23741] = 25'b01011100_10111011_00010111_1;
      patterns[23742] = 25'b01011100_10111100_00011000_1;
      patterns[23743] = 25'b01011100_10111101_00011001_1;
      patterns[23744] = 25'b01011100_10111110_00011010_1;
      patterns[23745] = 25'b01011100_10111111_00011011_1;
      patterns[23746] = 25'b01011100_11000000_00011100_1;
      patterns[23747] = 25'b01011100_11000001_00011101_1;
      patterns[23748] = 25'b01011100_11000010_00011110_1;
      patterns[23749] = 25'b01011100_11000011_00011111_1;
      patterns[23750] = 25'b01011100_11000100_00100000_1;
      patterns[23751] = 25'b01011100_11000101_00100001_1;
      patterns[23752] = 25'b01011100_11000110_00100010_1;
      patterns[23753] = 25'b01011100_11000111_00100011_1;
      patterns[23754] = 25'b01011100_11001000_00100100_1;
      patterns[23755] = 25'b01011100_11001001_00100101_1;
      patterns[23756] = 25'b01011100_11001010_00100110_1;
      patterns[23757] = 25'b01011100_11001011_00100111_1;
      patterns[23758] = 25'b01011100_11001100_00101000_1;
      patterns[23759] = 25'b01011100_11001101_00101001_1;
      patterns[23760] = 25'b01011100_11001110_00101010_1;
      patterns[23761] = 25'b01011100_11001111_00101011_1;
      patterns[23762] = 25'b01011100_11010000_00101100_1;
      patterns[23763] = 25'b01011100_11010001_00101101_1;
      patterns[23764] = 25'b01011100_11010010_00101110_1;
      patterns[23765] = 25'b01011100_11010011_00101111_1;
      patterns[23766] = 25'b01011100_11010100_00110000_1;
      patterns[23767] = 25'b01011100_11010101_00110001_1;
      patterns[23768] = 25'b01011100_11010110_00110010_1;
      patterns[23769] = 25'b01011100_11010111_00110011_1;
      patterns[23770] = 25'b01011100_11011000_00110100_1;
      patterns[23771] = 25'b01011100_11011001_00110101_1;
      patterns[23772] = 25'b01011100_11011010_00110110_1;
      patterns[23773] = 25'b01011100_11011011_00110111_1;
      patterns[23774] = 25'b01011100_11011100_00111000_1;
      patterns[23775] = 25'b01011100_11011101_00111001_1;
      patterns[23776] = 25'b01011100_11011110_00111010_1;
      patterns[23777] = 25'b01011100_11011111_00111011_1;
      patterns[23778] = 25'b01011100_11100000_00111100_1;
      patterns[23779] = 25'b01011100_11100001_00111101_1;
      patterns[23780] = 25'b01011100_11100010_00111110_1;
      patterns[23781] = 25'b01011100_11100011_00111111_1;
      patterns[23782] = 25'b01011100_11100100_01000000_1;
      patterns[23783] = 25'b01011100_11100101_01000001_1;
      patterns[23784] = 25'b01011100_11100110_01000010_1;
      patterns[23785] = 25'b01011100_11100111_01000011_1;
      patterns[23786] = 25'b01011100_11101000_01000100_1;
      patterns[23787] = 25'b01011100_11101001_01000101_1;
      patterns[23788] = 25'b01011100_11101010_01000110_1;
      patterns[23789] = 25'b01011100_11101011_01000111_1;
      patterns[23790] = 25'b01011100_11101100_01001000_1;
      patterns[23791] = 25'b01011100_11101101_01001001_1;
      patterns[23792] = 25'b01011100_11101110_01001010_1;
      patterns[23793] = 25'b01011100_11101111_01001011_1;
      patterns[23794] = 25'b01011100_11110000_01001100_1;
      patterns[23795] = 25'b01011100_11110001_01001101_1;
      patterns[23796] = 25'b01011100_11110010_01001110_1;
      patterns[23797] = 25'b01011100_11110011_01001111_1;
      patterns[23798] = 25'b01011100_11110100_01010000_1;
      patterns[23799] = 25'b01011100_11110101_01010001_1;
      patterns[23800] = 25'b01011100_11110110_01010010_1;
      patterns[23801] = 25'b01011100_11110111_01010011_1;
      patterns[23802] = 25'b01011100_11111000_01010100_1;
      patterns[23803] = 25'b01011100_11111001_01010101_1;
      patterns[23804] = 25'b01011100_11111010_01010110_1;
      patterns[23805] = 25'b01011100_11111011_01010111_1;
      patterns[23806] = 25'b01011100_11111100_01011000_1;
      patterns[23807] = 25'b01011100_11111101_01011001_1;
      patterns[23808] = 25'b01011100_11111110_01011010_1;
      patterns[23809] = 25'b01011100_11111111_01011011_1;
      patterns[23810] = 25'b01011101_00000000_01011101_0;
      patterns[23811] = 25'b01011101_00000001_01011110_0;
      patterns[23812] = 25'b01011101_00000010_01011111_0;
      patterns[23813] = 25'b01011101_00000011_01100000_0;
      patterns[23814] = 25'b01011101_00000100_01100001_0;
      patterns[23815] = 25'b01011101_00000101_01100010_0;
      patterns[23816] = 25'b01011101_00000110_01100011_0;
      patterns[23817] = 25'b01011101_00000111_01100100_0;
      patterns[23818] = 25'b01011101_00001000_01100101_0;
      patterns[23819] = 25'b01011101_00001001_01100110_0;
      patterns[23820] = 25'b01011101_00001010_01100111_0;
      patterns[23821] = 25'b01011101_00001011_01101000_0;
      patterns[23822] = 25'b01011101_00001100_01101001_0;
      patterns[23823] = 25'b01011101_00001101_01101010_0;
      patterns[23824] = 25'b01011101_00001110_01101011_0;
      patterns[23825] = 25'b01011101_00001111_01101100_0;
      patterns[23826] = 25'b01011101_00010000_01101101_0;
      patterns[23827] = 25'b01011101_00010001_01101110_0;
      patterns[23828] = 25'b01011101_00010010_01101111_0;
      patterns[23829] = 25'b01011101_00010011_01110000_0;
      patterns[23830] = 25'b01011101_00010100_01110001_0;
      patterns[23831] = 25'b01011101_00010101_01110010_0;
      patterns[23832] = 25'b01011101_00010110_01110011_0;
      patterns[23833] = 25'b01011101_00010111_01110100_0;
      patterns[23834] = 25'b01011101_00011000_01110101_0;
      patterns[23835] = 25'b01011101_00011001_01110110_0;
      patterns[23836] = 25'b01011101_00011010_01110111_0;
      patterns[23837] = 25'b01011101_00011011_01111000_0;
      patterns[23838] = 25'b01011101_00011100_01111001_0;
      patterns[23839] = 25'b01011101_00011101_01111010_0;
      patterns[23840] = 25'b01011101_00011110_01111011_0;
      patterns[23841] = 25'b01011101_00011111_01111100_0;
      patterns[23842] = 25'b01011101_00100000_01111101_0;
      patterns[23843] = 25'b01011101_00100001_01111110_0;
      patterns[23844] = 25'b01011101_00100010_01111111_0;
      patterns[23845] = 25'b01011101_00100011_10000000_0;
      patterns[23846] = 25'b01011101_00100100_10000001_0;
      patterns[23847] = 25'b01011101_00100101_10000010_0;
      patterns[23848] = 25'b01011101_00100110_10000011_0;
      patterns[23849] = 25'b01011101_00100111_10000100_0;
      patterns[23850] = 25'b01011101_00101000_10000101_0;
      patterns[23851] = 25'b01011101_00101001_10000110_0;
      patterns[23852] = 25'b01011101_00101010_10000111_0;
      patterns[23853] = 25'b01011101_00101011_10001000_0;
      patterns[23854] = 25'b01011101_00101100_10001001_0;
      patterns[23855] = 25'b01011101_00101101_10001010_0;
      patterns[23856] = 25'b01011101_00101110_10001011_0;
      patterns[23857] = 25'b01011101_00101111_10001100_0;
      patterns[23858] = 25'b01011101_00110000_10001101_0;
      patterns[23859] = 25'b01011101_00110001_10001110_0;
      patterns[23860] = 25'b01011101_00110010_10001111_0;
      patterns[23861] = 25'b01011101_00110011_10010000_0;
      patterns[23862] = 25'b01011101_00110100_10010001_0;
      patterns[23863] = 25'b01011101_00110101_10010010_0;
      patterns[23864] = 25'b01011101_00110110_10010011_0;
      patterns[23865] = 25'b01011101_00110111_10010100_0;
      patterns[23866] = 25'b01011101_00111000_10010101_0;
      patterns[23867] = 25'b01011101_00111001_10010110_0;
      patterns[23868] = 25'b01011101_00111010_10010111_0;
      patterns[23869] = 25'b01011101_00111011_10011000_0;
      patterns[23870] = 25'b01011101_00111100_10011001_0;
      patterns[23871] = 25'b01011101_00111101_10011010_0;
      patterns[23872] = 25'b01011101_00111110_10011011_0;
      patterns[23873] = 25'b01011101_00111111_10011100_0;
      patterns[23874] = 25'b01011101_01000000_10011101_0;
      patterns[23875] = 25'b01011101_01000001_10011110_0;
      patterns[23876] = 25'b01011101_01000010_10011111_0;
      patterns[23877] = 25'b01011101_01000011_10100000_0;
      patterns[23878] = 25'b01011101_01000100_10100001_0;
      patterns[23879] = 25'b01011101_01000101_10100010_0;
      patterns[23880] = 25'b01011101_01000110_10100011_0;
      patterns[23881] = 25'b01011101_01000111_10100100_0;
      patterns[23882] = 25'b01011101_01001000_10100101_0;
      patterns[23883] = 25'b01011101_01001001_10100110_0;
      patterns[23884] = 25'b01011101_01001010_10100111_0;
      patterns[23885] = 25'b01011101_01001011_10101000_0;
      patterns[23886] = 25'b01011101_01001100_10101001_0;
      patterns[23887] = 25'b01011101_01001101_10101010_0;
      patterns[23888] = 25'b01011101_01001110_10101011_0;
      patterns[23889] = 25'b01011101_01001111_10101100_0;
      patterns[23890] = 25'b01011101_01010000_10101101_0;
      patterns[23891] = 25'b01011101_01010001_10101110_0;
      patterns[23892] = 25'b01011101_01010010_10101111_0;
      patterns[23893] = 25'b01011101_01010011_10110000_0;
      patterns[23894] = 25'b01011101_01010100_10110001_0;
      patterns[23895] = 25'b01011101_01010101_10110010_0;
      patterns[23896] = 25'b01011101_01010110_10110011_0;
      patterns[23897] = 25'b01011101_01010111_10110100_0;
      patterns[23898] = 25'b01011101_01011000_10110101_0;
      patterns[23899] = 25'b01011101_01011001_10110110_0;
      patterns[23900] = 25'b01011101_01011010_10110111_0;
      patterns[23901] = 25'b01011101_01011011_10111000_0;
      patterns[23902] = 25'b01011101_01011100_10111001_0;
      patterns[23903] = 25'b01011101_01011101_10111010_0;
      patterns[23904] = 25'b01011101_01011110_10111011_0;
      patterns[23905] = 25'b01011101_01011111_10111100_0;
      patterns[23906] = 25'b01011101_01100000_10111101_0;
      patterns[23907] = 25'b01011101_01100001_10111110_0;
      patterns[23908] = 25'b01011101_01100010_10111111_0;
      patterns[23909] = 25'b01011101_01100011_11000000_0;
      patterns[23910] = 25'b01011101_01100100_11000001_0;
      patterns[23911] = 25'b01011101_01100101_11000010_0;
      patterns[23912] = 25'b01011101_01100110_11000011_0;
      patterns[23913] = 25'b01011101_01100111_11000100_0;
      patterns[23914] = 25'b01011101_01101000_11000101_0;
      patterns[23915] = 25'b01011101_01101001_11000110_0;
      patterns[23916] = 25'b01011101_01101010_11000111_0;
      patterns[23917] = 25'b01011101_01101011_11001000_0;
      patterns[23918] = 25'b01011101_01101100_11001001_0;
      patterns[23919] = 25'b01011101_01101101_11001010_0;
      patterns[23920] = 25'b01011101_01101110_11001011_0;
      patterns[23921] = 25'b01011101_01101111_11001100_0;
      patterns[23922] = 25'b01011101_01110000_11001101_0;
      patterns[23923] = 25'b01011101_01110001_11001110_0;
      patterns[23924] = 25'b01011101_01110010_11001111_0;
      patterns[23925] = 25'b01011101_01110011_11010000_0;
      patterns[23926] = 25'b01011101_01110100_11010001_0;
      patterns[23927] = 25'b01011101_01110101_11010010_0;
      patterns[23928] = 25'b01011101_01110110_11010011_0;
      patterns[23929] = 25'b01011101_01110111_11010100_0;
      patterns[23930] = 25'b01011101_01111000_11010101_0;
      patterns[23931] = 25'b01011101_01111001_11010110_0;
      patterns[23932] = 25'b01011101_01111010_11010111_0;
      patterns[23933] = 25'b01011101_01111011_11011000_0;
      patterns[23934] = 25'b01011101_01111100_11011001_0;
      patterns[23935] = 25'b01011101_01111101_11011010_0;
      patterns[23936] = 25'b01011101_01111110_11011011_0;
      patterns[23937] = 25'b01011101_01111111_11011100_0;
      patterns[23938] = 25'b01011101_10000000_11011101_0;
      patterns[23939] = 25'b01011101_10000001_11011110_0;
      patterns[23940] = 25'b01011101_10000010_11011111_0;
      patterns[23941] = 25'b01011101_10000011_11100000_0;
      patterns[23942] = 25'b01011101_10000100_11100001_0;
      patterns[23943] = 25'b01011101_10000101_11100010_0;
      patterns[23944] = 25'b01011101_10000110_11100011_0;
      patterns[23945] = 25'b01011101_10000111_11100100_0;
      patterns[23946] = 25'b01011101_10001000_11100101_0;
      patterns[23947] = 25'b01011101_10001001_11100110_0;
      patterns[23948] = 25'b01011101_10001010_11100111_0;
      patterns[23949] = 25'b01011101_10001011_11101000_0;
      patterns[23950] = 25'b01011101_10001100_11101001_0;
      patterns[23951] = 25'b01011101_10001101_11101010_0;
      patterns[23952] = 25'b01011101_10001110_11101011_0;
      patterns[23953] = 25'b01011101_10001111_11101100_0;
      patterns[23954] = 25'b01011101_10010000_11101101_0;
      patterns[23955] = 25'b01011101_10010001_11101110_0;
      patterns[23956] = 25'b01011101_10010010_11101111_0;
      patterns[23957] = 25'b01011101_10010011_11110000_0;
      patterns[23958] = 25'b01011101_10010100_11110001_0;
      patterns[23959] = 25'b01011101_10010101_11110010_0;
      patterns[23960] = 25'b01011101_10010110_11110011_0;
      patterns[23961] = 25'b01011101_10010111_11110100_0;
      patterns[23962] = 25'b01011101_10011000_11110101_0;
      patterns[23963] = 25'b01011101_10011001_11110110_0;
      patterns[23964] = 25'b01011101_10011010_11110111_0;
      patterns[23965] = 25'b01011101_10011011_11111000_0;
      patterns[23966] = 25'b01011101_10011100_11111001_0;
      patterns[23967] = 25'b01011101_10011101_11111010_0;
      patterns[23968] = 25'b01011101_10011110_11111011_0;
      patterns[23969] = 25'b01011101_10011111_11111100_0;
      patterns[23970] = 25'b01011101_10100000_11111101_0;
      patterns[23971] = 25'b01011101_10100001_11111110_0;
      patterns[23972] = 25'b01011101_10100010_11111111_0;
      patterns[23973] = 25'b01011101_10100011_00000000_1;
      patterns[23974] = 25'b01011101_10100100_00000001_1;
      patterns[23975] = 25'b01011101_10100101_00000010_1;
      patterns[23976] = 25'b01011101_10100110_00000011_1;
      patterns[23977] = 25'b01011101_10100111_00000100_1;
      patterns[23978] = 25'b01011101_10101000_00000101_1;
      patterns[23979] = 25'b01011101_10101001_00000110_1;
      patterns[23980] = 25'b01011101_10101010_00000111_1;
      patterns[23981] = 25'b01011101_10101011_00001000_1;
      patterns[23982] = 25'b01011101_10101100_00001001_1;
      patterns[23983] = 25'b01011101_10101101_00001010_1;
      patterns[23984] = 25'b01011101_10101110_00001011_1;
      patterns[23985] = 25'b01011101_10101111_00001100_1;
      patterns[23986] = 25'b01011101_10110000_00001101_1;
      patterns[23987] = 25'b01011101_10110001_00001110_1;
      patterns[23988] = 25'b01011101_10110010_00001111_1;
      patterns[23989] = 25'b01011101_10110011_00010000_1;
      patterns[23990] = 25'b01011101_10110100_00010001_1;
      patterns[23991] = 25'b01011101_10110101_00010010_1;
      patterns[23992] = 25'b01011101_10110110_00010011_1;
      patterns[23993] = 25'b01011101_10110111_00010100_1;
      patterns[23994] = 25'b01011101_10111000_00010101_1;
      patterns[23995] = 25'b01011101_10111001_00010110_1;
      patterns[23996] = 25'b01011101_10111010_00010111_1;
      patterns[23997] = 25'b01011101_10111011_00011000_1;
      patterns[23998] = 25'b01011101_10111100_00011001_1;
      patterns[23999] = 25'b01011101_10111101_00011010_1;
      patterns[24000] = 25'b01011101_10111110_00011011_1;
      patterns[24001] = 25'b01011101_10111111_00011100_1;
      patterns[24002] = 25'b01011101_11000000_00011101_1;
      patterns[24003] = 25'b01011101_11000001_00011110_1;
      patterns[24004] = 25'b01011101_11000010_00011111_1;
      patterns[24005] = 25'b01011101_11000011_00100000_1;
      patterns[24006] = 25'b01011101_11000100_00100001_1;
      patterns[24007] = 25'b01011101_11000101_00100010_1;
      patterns[24008] = 25'b01011101_11000110_00100011_1;
      patterns[24009] = 25'b01011101_11000111_00100100_1;
      patterns[24010] = 25'b01011101_11001000_00100101_1;
      patterns[24011] = 25'b01011101_11001001_00100110_1;
      patterns[24012] = 25'b01011101_11001010_00100111_1;
      patterns[24013] = 25'b01011101_11001011_00101000_1;
      patterns[24014] = 25'b01011101_11001100_00101001_1;
      patterns[24015] = 25'b01011101_11001101_00101010_1;
      patterns[24016] = 25'b01011101_11001110_00101011_1;
      patterns[24017] = 25'b01011101_11001111_00101100_1;
      patterns[24018] = 25'b01011101_11010000_00101101_1;
      patterns[24019] = 25'b01011101_11010001_00101110_1;
      patterns[24020] = 25'b01011101_11010010_00101111_1;
      patterns[24021] = 25'b01011101_11010011_00110000_1;
      patterns[24022] = 25'b01011101_11010100_00110001_1;
      patterns[24023] = 25'b01011101_11010101_00110010_1;
      patterns[24024] = 25'b01011101_11010110_00110011_1;
      patterns[24025] = 25'b01011101_11010111_00110100_1;
      patterns[24026] = 25'b01011101_11011000_00110101_1;
      patterns[24027] = 25'b01011101_11011001_00110110_1;
      patterns[24028] = 25'b01011101_11011010_00110111_1;
      patterns[24029] = 25'b01011101_11011011_00111000_1;
      patterns[24030] = 25'b01011101_11011100_00111001_1;
      patterns[24031] = 25'b01011101_11011101_00111010_1;
      patterns[24032] = 25'b01011101_11011110_00111011_1;
      patterns[24033] = 25'b01011101_11011111_00111100_1;
      patterns[24034] = 25'b01011101_11100000_00111101_1;
      patterns[24035] = 25'b01011101_11100001_00111110_1;
      patterns[24036] = 25'b01011101_11100010_00111111_1;
      patterns[24037] = 25'b01011101_11100011_01000000_1;
      patterns[24038] = 25'b01011101_11100100_01000001_1;
      patterns[24039] = 25'b01011101_11100101_01000010_1;
      patterns[24040] = 25'b01011101_11100110_01000011_1;
      patterns[24041] = 25'b01011101_11100111_01000100_1;
      patterns[24042] = 25'b01011101_11101000_01000101_1;
      patterns[24043] = 25'b01011101_11101001_01000110_1;
      patterns[24044] = 25'b01011101_11101010_01000111_1;
      patterns[24045] = 25'b01011101_11101011_01001000_1;
      patterns[24046] = 25'b01011101_11101100_01001001_1;
      patterns[24047] = 25'b01011101_11101101_01001010_1;
      patterns[24048] = 25'b01011101_11101110_01001011_1;
      patterns[24049] = 25'b01011101_11101111_01001100_1;
      patterns[24050] = 25'b01011101_11110000_01001101_1;
      patterns[24051] = 25'b01011101_11110001_01001110_1;
      patterns[24052] = 25'b01011101_11110010_01001111_1;
      patterns[24053] = 25'b01011101_11110011_01010000_1;
      patterns[24054] = 25'b01011101_11110100_01010001_1;
      patterns[24055] = 25'b01011101_11110101_01010010_1;
      patterns[24056] = 25'b01011101_11110110_01010011_1;
      patterns[24057] = 25'b01011101_11110111_01010100_1;
      patterns[24058] = 25'b01011101_11111000_01010101_1;
      patterns[24059] = 25'b01011101_11111001_01010110_1;
      patterns[24060] = 25'b01011101_11111010_01010111_1;
      patterns[24061] = 25'b01011101_11111011_01011000_1;
      patterns[24062] = 25'b01011101_11111100_01011001_1;
      patterns[24063] = 25'b01011101_11111101_01011010_1;
      patterns[24064] = 25'b01011101_11111110_01011011_1;
      patterns[24065] = 25'b01011101_11111111_01011100_1;
      patterns[24066] = 25'b01011110_00000000_01011110_0;
      patterns[24067] = 25'b01011110_00000001_01011111_0;
      patterns[24068] = 25'b01011110_00000010_01100000_0;
      patterns[24069] = 25'b01011110_00000011_01100001_0;
      patterns[24070] = 25'b01011110_00000100_01100010_0;
      patterns[24071] = 25'b01011110_00000101_01100011_0;
      patterns[24072] = 25'b01011110_00000110_01100100_0;
      patterns[24073] = 25'b01011110_00000111_01100101_0;
      patterns[24074] = 25'b01011110_00001000_01100110_0;
      patterns[24075] = 25'b01011110_00001001_01100111_0;
      patterns[24076] = 25'b01011110_00001010_01101000_0;
      patterns[24077] = 25'b01011110_00001011_01101001_0;
      patterns[24078] = 25'b01011110_00001100_01101010_0;
      patterns[24079] = 25'b01011110_00001101_01101011_0;
      patterns[24080] = 25'b01011110_00001110_01101100_0;
      patterns[24081] = 25'b01011110_00001111_01101101_0;
      patterns[24082] = 25'b01011110_00010000_01101110_0;
      patterns[24083] = 25'b01011110_00010001_01101111_0;
      patterns[24084] = 25'b01011110_00010010_01110000_0;
      patterns[24085] = 25'b01011110_00010011_01110001_0;
      patterns[24086] = 25'b01011110_00010100_01110010_0;
      patterns[24087] = 25'b01011110_00010101_01110011_0;
      patterns[24088] = 25'b01011110_00010110_01110100_0;
      patterns[24089] = 25'b01011110_00010111_01110101_0;
      patterns[24090] = 25'b01011110_00011000_01110110_0;
      patterns[24091] = 25'b01011110_00011001_01110111_0;
      patterns[24092] = 25'b01011110_00011010_01111000_0;
      patterns[24093] = 25'b01011110_00011011_01111001_0;
      patterns[24094] = 25'b01011110_00011100_01111010_0;
      patterns[24095] = 25'b01011110_00011101_01111011_0;
      patterns[24096] = 25'b01011110_00011110_01111100_0;
      patterns[24097] = 25'b01011110_00011111_01111101_0;
      patterns[24098] = 25'b01011110_00100000_01111110_0;
      patterns[24099] = 25'b01011110_00100001_01111111_0;
      patterns[24100] = 25'b01011110_00100010_10000000_0;
      patterns[24101] = 25'b01011110_00100011_10000001_0;
      patterns[24102] = 25'b01011110_00100100_10000010_0;
      patterns[24103] = 25'b01011110_00100101_10000011_0;
      patterns[24104] = 25'b01011110_00100110_10000100_0;
      patterns[24105] = 25'b01011110_00100111_10000101_0;
      patterns[24106] = 25'b01011110_00101000_10000110_0;
      patterns[24107] = 25'b01011110_00101001_10000111_0;
      patterns[24108] = 25'b01011110_00101010_10001000_0;
      patterns[24109] = 25'b01011110_00101011_10001001_0;
      patterns[24110] = 25'b01011110_00101100_10001010_0;
      patterns[24111] = 25'b01011110_00101101_10001011_0;
      patterns[24112] = 25'b01011110_00101110_10001100_0;
      patterns[24113] = 25'b01011110_00101111_10001101_0;
      patterns[24114] = 25'b01011110_00110000_10001110_0;
      patterns[24115] = 25'b01011110_00110001_10001111_0;
      patterns[24116] = 25'b01011110_00110010_10010000_0;
      patterns[24117] = 25'b01011110_00110011_10010001_0;
      patterns[24118] = 25'b01011110_00110100_10010010_0;
      patterns[24119] = 25'b01011110_00110101_10010011_0;
      patterns[24120] = 25'b01011110_00110110_10010100_0;
      patterns[24121] = 25'b01011110_00110111_10010101_0;
      patterns[24122] = 25'b01011110_00111000_10010110_0;
      patterns[24123] = 25'b01011110_00111001_10010111_0;
      patterns[24124] = 25'b01011110_00111010_10011000_0;
      patterns[24125] = 25'b01011110_00111011_10011001_0;
      patterns[24126] = 25'b01011110_00111100_10011010_0;
      patterns[24127] = 25'b01011110_00111101_10011011_0;
      patterns[24128] = 25'b01011110_00111110_10011100_0;
      patterns[24129] = 25'b01011110_00111111_10011101_0;
      patterns[24130] = 25'b01011110_01000000_10011110_0;
      patterns[24131] = 25'b01011110_01000001_10011111_0;
      patterns[24132] = 25'b01011110_01000010_10100000_0;
      patterns[24133] = 25'b01011110_01000011_10100001_0;
      patterns[24134] = 25'b01011110_01000100_10100010_0;
      patterns[24135] = 25'b01011110_01000101_10100011_0;
      patterns[24136] = 25'b01011110_01000110_10100100_0;
      patterns[24137] = 25'b01011110_01000111_10100101_0;
      patterns[24138] = 25'b01011110_01001000_10100110_0;
      patterns[24139] = 25'b01011110_01001001_10100111_0;
      patterns[24140] = 25'b01011110_01001010_10101000_0;
      patterns[24141] = 25'b01011110_01001011_10101001_0;
      patterns[24142] = 25'b01011110_01001100_10101010_0;
      patterns[24143] = 25'b01011110_01001101_10101011_0;
      patterns[24144] = 25'b01011110_01001110_10101100_0;
      patterns[24145] = 25'b01011110_01001111_10101101_0;
      patterns[24146] = 25'b01011110_01010000_10101110_0;
      patterns[24147] = 25'b01011110_01010001_10101111_0;
      patterns[24148] = 25'b01011110_01010010_10110000_0;
      patterns[24149] = 25'b01011110_01010011_10110001_0;
      patterns[24150] = 25'b01011110_01010100_10110010_0;
      patterns[24151] = 25'b01011110_01010101_10110011_0;
      patterns[24152] = 25'b01011110_01010110_10110100_0;
      patterns[24153] = 25'b01011110_01010111_10110101_0;
      patterns[24154] = 25'b01011110_01011000_10110110_0;
      patterns[24155] = 25'b01011110_01011001_10110111_0;
      patterns[24156] = 25'b01011110_01011010_10111000_0;
      patterns[24157] = 25'b01011110_01011011_10111001_0;
      patterns[24158] = 25'b01011110_01011100_10111010_0;
      patterns[24159] = 25'b01011110_01011101_10111011_0;
      patterns[24160] = 25'b01011110_01011110_10111100_0;
      patterns[24161] = 25'b01011110_01011111_10111101_0;
      patterns[24162] = 25'b01011110_01100000_10111110_0;
      patterns[24163] = 25'b01011110_01100001_10111111_0;
      patterns[24164] = 25'b01011110_01100010_11000000_0;
      patterns[24165] = 25'b01011110_01100011_11000001_0;
      patterns[24166] = 25'b01011110_01100100_11000010_0;
      patterns[24167] = 25'b01011110_01100101_11000011_0;
      patterns[24168] = 25'b01011110_01100110_11000100_0;
      patterns[24169] = 25'b01011110_01100111_11000101_0;
      patterns[24170] = 25'b01011110_01101000_11000110_0;
      patterns[24171] = 25'b01011110_01101001_11000111_0;
      patterns[24172] = 25'b01011110_01101010_11001000_0;
      patterns[24173] = 25'b01011110_01101011_11001001_0;
      patterns[24174] = 25'b01011110_01101100_11001010_0;
      patterns[24175] = 25'b01011110_01101101_11001011_0;
      patterns[24176] = 25'b01011110_01101110_11001100_0;
      patterns[24177] = 25'b01011110_01101111_11001101_0;
      patterns[24178] = 25'b01011110_01110000_11001110_0;
      patterns[24179] = 25'b01011110_01110001_11001111_0;
      patterns[24180] = 25'b01011110_01110010_11010000_0;
      patterns[24181] = 25'b01011110_01110011_11010001_0;
      patterns[24182] = 25'b01011110_01110100_11010010_0;
      patterns[24183] = 25'b01011110_01110101_11010011_0;
      patterns[24184] = 25'b01011110_01110110_11010100_0;
      patterns[24185] = 25'b01011110_01110111_11010101_0;
      patterns[24186] = 25'b01011110_01111000_11010110_0;
      patterns[24187] = 25'b01011110_01111001_11010111_0;
      patterns[24188] = 25'b01011110_01111010_11011000_0;
      patterns[24189] = 25'b01011110_01111011_11011001_0;
      patterns[24190] = 25'b01011110_01111100_11011010_0;
      patterns[24191] = 25'b01011110_01111101_11011011_0;
      patterns[24192] = 25'b01011110_01111110_11011100_0;
      patterns[24193] = 25'b01011110_01111111_11011101_0;
      patterns[24194] = 25'b01011110_10000000_11011110_0;
      patterns[24195] = 25'b01011110_10000001_11011111_0;
      patterns[24196] = 25'b01011110_10000010_11100000_0;
      patterns[24197] = 25'b01011110_10000011_11100001_0;
      patterns[24198] = 25'b01011110_10000100_11100010_0;
      patterns[24199] = 25'b01011110_10000101_11100011_0;
      patterns[24200] = 25'b01011110_10000110_11100100_0;
      patterns[24201] = 25'b01011110_10000111_11100101_0;
      patterns[24202] = 25'b01011110_10001000_11100110_0;
      patterns[24203] = 25'b01011110_10001001_11100111_0;
      patterns[24204] = 25'b01011110_10001010_11101000_0;
      patterns[24205] = 25'b01011110_10001011_11101001_0;
      patterns[24206] = 25'b01011110_10001100_11101010_0;
      patterns[24207] = 25'b01011110_10001101_11101011_0;
      patterns[24208] = 25'b01011110_10001110_11101100_0;
      patterns[24209] = 25'b01011110_10001111_11101101_0;
      patterns[24210] = 25'b01011110_10010000_11101110_0;
      patterns[24211] = 25'b01011110_10010001_11101111_0;
      patterns[24212] = 25'b01011110_10010010_11110000_0;
      patterns[24213] = 25'b01011110_10010011_11110001_0;
      patterns[24214] = 25'b01011110_10010100_11110010_0;
      patterns[24215] = 25'b01011110_10010101_11110011_0;
      patterns[24216] = 25'b01011110_10010110_11110100_0;
      patterns[24217] = 25'b01011110_10010111_11110101_0;
      patterns[24218] = 25'b01011110_10011000_11110110_0;
      patterns[24219] = 25'b01011110_10011001_11110111_0;
      patterns[24220] = 25'b01011110_10011010_11111000_0;
      patterns[24221] = 25'b01011110_10011011_11111001_0;
      patterns[24222] = 25'b01011110_10011100_11111010_0;
      patterns[24223] = 25'b01011110_10011101_11111011_0;
      patterns[24224] = 25'b01011110_10011110_11111100_0;
      patterns[24225] = 25'b01011110_10011111_11111101_0;
      patterns[24226] = 25'b01011110_10100000_11111110_0;
      patterns[24227] = 25'b01011110_10100001_11111111_0;
      patterns[24228] = 25'b01011110_10100010_00000000_1;
      patterns[24229] = 25'b01011110_10100011_00000001_1;
      patterns[24230] = 25'b01011110_10100100_00000010_1;
      patterns[24231] = 25'b01011110_10100101_00000011_1;
      patterns[24232] = 25'b01011110_10100110_00000100_1;
      patterns[24233] = 25'b01011110_10100111_00000101_1;
      patterns[24234] = 25'b01011110_10101000_00000110_1;
      patterns[24235] = 25'b01011110_10101001_00000111_1;
      patterns[24236] = 25'b01011110_10101010_00001000_1;
      patterns[24237] = 25'b01011110_10101011_00001001_1;
      patterns[24238] = 25'b01011110_10101100_00001010_1;
      patterns[24239] = 25'b01011110_10101101_00001011_1;
      patterns[24240] = 25'b01011110_10101110_00001100_1;
      patterns[24241] = 25'b01011110_10101111_00001101_1;
      patterns[24242] = 25'b01011110_10110000_00001110_1;
      patterns[24243] = 25'b01011110_10110001_00001111_1;
      patterns[24244] = 25'b01011110_10110010_00010000_1;
      patterns[24245] = 25'b01011110_10110011_00010001_1;
      patterns[24246] = 25'b01011110_10110100_00010010_1;
      patterns[24247] = 25'b01011110_10110101_00010011_1;
      patterns[24248] = 25'b01011110_10110110_00010100_1;
      patterns[24249] = 25'b01011110_10110111_00010101_1;
      patterns[24250] = 25'b01011110_10111000_00010110_1;
      patterns[24251] = 25'b01011110_10111001_00010111_1;
      patterns[24252] = 25'b01011110_10111010_00011000_1;
      patterns[24253] = 25'b01011110_10111011_00011001_1;
      patterns[24254] = 25'b01011110_10111100_00011010_1;
      patterns[24255] = 25'b01011110_10111101_00011011_1;
      patterns[24256] = 25'b01011110_10111110_00011100_1;
      patterns[24257] = 25'b01011110_10111111_00011101_1;
      patterns[24258] = 25'b01011110_11000000_00011110_1;
      patterns[24259] = 25'b01011110_11000001_00011111_1;
      patterns[24260] = 25'b01011110_11000010_00100000_1;
      patterns[24261] = 25'b01011110_11000011_00100001_1;
      patterns[24262] = 25'b01011110_11000100_00100010_1;
      patterns[24263] = 25'b01011110_11000101_00100011_1;
      patterns[24264] = 25'b01011110_11000110_00100100_1;
      patterns[24265] = 25'b01011110_11000111_00100101_1;
      patterns[24266] = 25'b01011110_11001000_00100110_1;
      patterns[24267] = 25'b01011110_11001001_00100111_1;
      patterns[24268] = 25'b01011110_11001010_00101000_1;
      patterns[24269] = 25'b01011110_11001011_00101001_1;
      patterns[24270] = 25'b01011110_11001100_00101010_1;
      patterns[24271] = 25'b01011110_11001101_00101011_1;
      patterns[24272] = 25'b01011110_11001110_00101100_1;
      patterns[24273] = 25'b01011110_11001111_00101101_1;
      patterns[24274] = 25'b01011110_11010000_00101110_1;
      patterns[24275] = 25'b01011110_11010001_00101111_1;
      patterns[24276] = 25'b01011110_11010010_00110000_1;
      patterns[24277] = 25'b01011110_11010011_00110001_1;
      patterns[24278] = 25'b01011110_11010100_00110010_1;
      patterns[24279] = 25'b01011110_11010101_00110011_1;
      patterns[24280] = 25'b01011110_11010110_00110100_1;
      patterns[24281] = 25'b01011110_11010111_00110101_1;
      patterns[24282] = 25'b01011110_11011000_00110110_1;
      patterns[24283] = 25'b01011110_11011001_00110111_1;
      patterns[24284] = 25'b01011110_11011010_00111000_1;
      patterns[24285] = 25'b01011110_11011011_00111001_1;
      patterns[24286] = 25'b01011110_11011100_00111010_1;
      patterns[24287] = 25'b01011110_11011101_00111011_1;
      patterns[24288] = 25'b01011110_11011110_00111100_1;
      patterns[24289] = 25'b01011110_11011111_00111101_1;
      patterns[24290] = 25'b01011110_11100000_00111110_1;
      patterns[24291] = 25'b01011110_11100001_00111111_1;
      patterns[24292] = 25'b01011110_11100010_01000000_1;
      patterns[24293] = 25'b01011110_11100011_01000001_1;
      patterns[24294] = 25'b01011110_11100100_01000010_1;
      patterns[24295] = 25'b01011110_11100101_01000011_1;
      patterns[24296] = 25'b01011110_11100110_01000100_1;
      patterns[24297] = 25'b01011110_11100111_01000101_1;
      patterns[24298] = 25'b01011110_11101000_01000110_1;
      patterns[24299] = 25'b01011110_11101001_01000111_1;
      patterns[24300] = 25'b01011110_11101010_01001000_1;
      patterns[24301] = 25'b01011110_11101011_01001001_1;
      patterns[24302] = 25'b01011110_11101100_01001010_1;
      patterns[24303] = 25'b01011110_11101101_01001011_1;
      patterns[24304] = 25'b01011110_11101110_01001100_1;
      patterns[24305] = 25'b01011110_11101111_01001101_1;
      patterns[24306] = 25'b01011110_11110000_01001110_1;
      patterns[24307] = 25'b01011110_11110001_01001111_1;
      patterns[24308] = 25'b01011110_11110010_01010000_1;
      patterns[24309] = 25'b01011110_11110011_01010001_1;
      patterns[24310] = 25'b01011110_11110100_01010010_1;
      patterns[24311] = 25'b01011110_11110101_01010011_1;
      patterns[24312] = 25'b01011110_11110110_01010100_1;
      patterns[24313] = 25'b01011110_11110111_01010101_1;
      patterns[24314] = 25'b01011110_11111000_01010110_1;
      patterns[24315] = 25'b01011110_11111001_01010111_1;
      patterns[24316] = 25'b01011110_11111010_01011000_1;
      patterns[24317] = 25'b01011110_11111011_01011001_1;
      patterns[24318] = 25'b01011110_11111100_01011010_1;
      patterns[24319] = 25'b01011110_11111101_01011011_1;
      patterns[24320] = 25'b01011110_11111110_01011100_1;
      patterns[24321] = 25'b01011110_11111111_01011101_1;
      patterns[24322] = 25'b01011111_00000000_01011111_0;
      patterns[24323] = 25'b01011111_00000001_01100000_0;
      patterns[24324] = 25'b01011111_00000010_01100001_0;
      patterns[24325] = 25'b01011111_00000011_01100010_0;
      patterns[24326] = 25'b01011111_00000100_01100011_0;
      patterns[24327] = 25'b01011111_00000101_01100100_0;
      patterns[24328] = 25'b01011111_00000110_01100101_0;
      patterns[24329] = 25'b01011111_00000111_01100110_0;
      patterns[24330] = 25'b01011111_00001000_01100111_0;
      patterns[24331] = 25'b01011111_00001001_01101000_0;
      patterns[24332] = 25'b01011111_00001010_01101001_0;
      patterns[24333] = 25'b01011111_00001011_01101010_0;
      patterns[24334] = 25'b01011111_00001100_01101011_0;
      patterns[24335] = 25'b01011111_00001101_01101100_0;
      patterns[24336] = 25'b01011111_00001110_01101101_0;
      patterns[24337] = 25'b01011111_00001111_01101110_0;
      patterns[24338] = 25'b01011111_00010000_01101111_0;
      patterns[24339] = 25'b01011111_00010001_01110000_0;
      patterns[24340] = 25'b01011111_00010010_01110001_0;
      patterns[24341] = 25'b01011111_00010011_01110010_0;
      patterns[24342] = 25'b01011111_00010100_01110011_0;
      patterns[24343] = 25'b01011111_00010101_01110100_0;
      patterns[24344] = 25'b01011111_00010110_01110101_0;
      patterns[24345] = 25'b01011111_00010111_01110110_0;
      patterns[24346] = 25'b01011111_00011000_01110111_0;
      patterns[24347] = 25'b01011111_00011001_01111000_0;
      patterns[24348] = 25'b01011111_00011010_01111001_0;
      patterns[24349] = 25'b01011111_00011011_01111010_0;
      patterns[24350] = 25'b01011111_00011100_01111011_0;
      patterns[24351] = 25'b01011111_00011101_01111100_0;
      patterns[24352] = 25'b01011111_00011110_01111101_0;
      patterns[24353] = 25'b01011111_00011111_01111110_0;
      patterns[24354] = 25'b01011111_00100000_01111111_0;
      patterns[24355] = 25'b01011111_00100001_10000000_0;
      patterns[24356] = 25'b01011111_00100010_10000001_0;
      patterns[24357] = 25'b01011111_00100011_10000010_0;
      patterns[24358] = 25'b01011111_00100100_10000011_0;
      patterns[24359] = 25'b01011111_00100101_10000100_0;
      patterns[24360] = 25'b01011111_00100110_10000101_0;
      patterns[24361] = 25'b01011111_00100111_10000110_0;
      patterns[24362] = 25'b01011111_00101000_10000111_0;
      patterns[24363] = 25'b01011111_00101001_10001000_0;
      patterns[24364] = 25'b01011111_00101010_10001001_0;
      patterns[24365] = 25'b01011111_00101011_10001010_0;
      patterns[24366] = 25'b01011111_00101100_10001011_0;
      patterns[24367] = 25'b01011111_00101101_10001100_0;
      patterns[24368] = 25'b01011111_00101110_10001101_0;
      patterns[24369] = 25'b01011111_00101111_10001110_0;
      patterns[24370] = 25'b01011111_00110000_10001111_0;
      patterns[24371] = 25'b01011111_00110001_10010000_0;
      patterns[24372] = 25'b01011111_00110010_10010001_0;
      patterns[24373] = 25'b01011111_00110011_10010010_0;
      patterns[24374] = 25'b01011111_00110100_10010011_0;
      patterns[24375] = 25'b01011111_00110101_10010100_0;
      patterns[24376] = 25'b01011111_00110110_10010101_0;
      patterns[24377] = 25'b01011111_00110111_10010110_0;
      patterns[24378] = 25'b01011111_00111000_10010111_0;
      patterns[24379] = 25'b01011111_00111001_10011000_0;
      patterns[24380] = 25'b01011111_00111010_10011001_0;
      patterns[24381] = 25'b01011111_00111011_10011010_0;
      patterns[24382] = 25'b01011111_00111100_10011011_0;
      patterns[24383] = 25'b01011111_00111101_10011100_0;
      patterns[24384] = 25'b01011111_00111110_10011101_0;
      patterns[24385] = 25'b01011111_00111111_10011110_0;
      patterns[24386] = 25'b01011111_01000000_10011111_0;
      patterns[24387] = 25'b01011111_01000001_10100000_0;
      patterns[24388] = 25'b01011111_01000010_10100001_0;
      patterns[24389] = 25'b01011111_01000011_10100010_0;
      patterns[24390] = 25'b01011111_01000100_10100011_0;
      patterns[24391] = 25'b01011111_01000101_10100100_0;
      patterns[24392] = 25'b01011111_01000110_10100101_0;
      patterns[24393] = 25'b01011111_01000111_10100110_0;
      patterns[24394] = 25'b01011111_01001000_10100111_0;
      patterns[24395] = 25'b01011111_01001001_10101000_0;
      patterns[24396] = 25'b01011111_01001010_10101001_0;
      patterns[24397] = 25'b01011111_01001011_10101010_0;
      patterns[24398] = 25'b01011111_01001100_10101011_0;
      patterns[24399] = 25'b01011111_01001101_10101100_0;
      patterns[24400] = 25'b01011111_01001110_10101101_0;
      patterns[24401] = 25'b01011111_01001111_10101110_0;
      patterns[24402] = 25'b01011111_01010000_10101111_0;
      patterns[24403] = 25'b01011111_01010001_10110000_0;
      patterns[24404] = 25'b01011111_01010010_10110001_0;
      patterns[24405] = 25'b01011111_01010011_10110010_0;
      patterns[24406] = 25'b01011111_01010100_10110011_0;
      patterns[24407] = 25'b01011111_01010101_10110100_0;
      patterns[24408] = 25'b01011111_01010110_10110101_0;
      patterns[24409] = 25'b01011111_01010111_10110110_0;
      patterns[24410] = 25'b01011111_01011000_10110111_0;
      patterns[24411] = 25'b01011111_01011001_10111000_0;
      patterns[24412] = 25'b01011111_01011010_10111001_0;
      patterns[24413] = 25'b01011111_01011011_10111010_0;
      patterns[24414] = 25'b01011111_01011100_10111011_0;
      patterns[24415] = 25'b01011111_01011101_10111100_0;
      patterns[24416] = 25'b01011111_01011110_10111101_0;
      patterns[24417] = 25'b01011111_01011111_10111110_0;
      patterns[24418] = 25'b01011111_01100000_10111111_0;
      patterns[24419] = 25'b01011111_01100001_11000000_0;
      patterns[24420] = 25'b01011111_01100010_11000001_0;
      patterns[24421] = 25'b01011111_01100011_11000010_0;
      patterns[24422] = 25'b01011111_01100100_11000011_0;
      patterns[24423] = 25'b01011111_01100101_11000100_0;
      patterns[24424] = 25'b01011111_01100110_11000101_0;
      patterns[24425] = 25'b01011111_01100111_11000110_0;
      patterns[24426] = 25'b01011111_01101000_11000111_0;
      patterns[24427] = 25'b01011111_01101001_11001000_0;
      patterns[24428] = 25'b01011111_01101010_11001001_0;
      patterns[24429] = 25'b01011111_01101011_11001010_0;
      patterns[24430] = 25'b01011111_01101100_11001011_0;
      patterns[24431] = 25'b01011111_01101101_11001100_0;
      patterns[24432] = 25'b01011111_01101110_11001101_0;
      patterns[24433] = 25'b01011111_01101111_11001110_0;
      patterns[24434] = 25'b01011111_01110000_11001111_0;
      patterns[24435] = 25'b01011111_01110001_11010000_0;
      patterns[24436] = 25'b01011111_01110010_11010001_0;
      patterns[24437] = 25'b01011111_01110011_11010010_0;
      patterns[24438] = 25'b01011111_01110100_11010011_0;
      patterns[24439] = 25'b01011111_01110101_11010100_0;
      patterns[24440] = 25'b01011111_01110110_11010101_0;
      patterns[24441] = 25'b01011111_01110111_11010110_0;
      patterns[24442] = 25'b01011111_01111000_11010111_0;
      patterns[24443] = 25'b01011111_01111001_11011000_0;
      patterns[24444] = 25'b01011111_01111010_11011001_0;
      patterns[24445] = 25'b01011111_01111011_11011010_0;
      patterns[24446] = 25'b01011111_01111100_11011011_0;
      patterns[24447] = 25'b01011111_01111101_11011100_0;
      patterns[24448] = 25'b01011111_01111110_11011101_0;
      patterns[24449] = 25'b01011111_01111111_11011110_0;
      patterns[24450] = 25'b01011111_10000000_11011111_0;
      patterns[24451] = 25'b01011111_10000001_11100000_0;
      patterns[24452] = 25'b01011111_10000010_11100001_0;
      patterns[24453] = 25'b01011111_10000011_11100010_0;
      patterns[24454] = 25'b01011111_10000100_11100011_0;
      patterns[24455] = 25'b01011111_10000101_11100100_0;
      patterns[24456] = 25'b01011111_10000110_11100101_0;
      patterns[24457] = 25'b01011111_10000111_11100110_0;
      patterns[24458] = 25'b01011111_10001000_11100111_0;
      patterns[24459] = 25'b01011111_10001001_11101000_0;
      patterns[24460] = 25'b01011111_10001010_11101001_0;
      patterns[24461] = 25'b01011111_10001011_11101010_0;
      patterns[24462] = 25'b01011111_10001100_11101011_0;
      patterns[24463] = 25'b01011111_10001101_11101100_0;
      patterns[24464] = 25'b01011111_10001110_11101101_0;
      patterns[24465] = 25'b01011111_10001111_11101110_0;
      patterns[24466] = 25'b01011111_10010000_11101111_0;
      patterns[24467] = 25'b01011111_10010001_11110000_0;
      patterns[24468] = 25'b01011111_10010010_11110001_0;
      patterns[24469] = 25'b01011111_10010011_11110010_0;
      patterns[24470] = 25'b01011111_10010100_11110011_0;
      patterns[24471] = 25'b01011111_10010101_11110100_0;
      patterns[24472] = 25'b01011111_10010110_11110101_0;
      patterns[24473] = 25'b01011111_10010111_11110110_0;
      patterns[24474] = 25'b01011111_10011000_11110111_0;
      patterns[24475] = 25'b01011111_10011001_11111000_0;
      patterns[24476] = 25'b01011111_10011010_11111001_0;
      patterns[24477] = 25'b01011111_10011011_11111010_0;
      patterns[24478] = 25'b01011111_10011100_11111011_0;
      patterns[24479] = 25'b01011111_10011101_11111100_0;
      patterns[24480] = 25'b01011111_10011110_11111101_0;
      patterns[24481] = 25'b01011111_10011111_11111110_0;
      patterns[24482] = 25'b01011111_10100000_11111111_0;
      patterns[24483] = 25'b01011111_10100001_00000000_1;
      patterns[24484] = 25'b01011111_10100010_00000001_1;
      patterns[24485] = 25'b01011111_10100011_00000010_1;
      patterns[24486] = 25'b01011111_10100100_00000011_1;
      patterns[24487] = 25'b01011111_10100101_00000100_1;
      patterns[24488] = 25'b01011111_10100110_00000101_1;
      patterns[24489] = 25'b01011111_10100111_00000110_1;
      patterns[24490] = 25'b01011111_10101000_00000111_1;
      patterns[24491] = 25'b01011111_10101001_00001000_1;
      patterns[24492] = 25'b01011111_10101010_00001001_1;
      patterns[24493] = 25'b01011111_10101011_00001010_1;
      patterns[24494] = 25'b01011111_10101100_00001011_1;
      patterns[24495] = 25'b01011111_10101101_00001100_1;
      patterns[24496] = 25'b01011111_10101110_00001101_1;
      patterns[24497] = 25'b01011111_10101111_00001110_1;
      patterns[24498] = 25'b01011111_10110000_00001111_1;
      patterns[24499] = 25'b01011111_10110001_00010000_1;
      patterns[24500] = 25'b01011111_10110010_00010001_1;
      patterns[24501] = 25'b01011111_10110011_00010010_1;
      patterns[24502] = 25'b01011111_10110100_00010011_1;
      patterns[24503] = 25'b01011111_10110101_00010100_1;
      patterns[24504] = 25'b01011111_10110110_00010101_1;
      patterns[24505] = 25'b01011111_10110111_00010110_1;
      patterns[24506] = 25'b01011111_10111000_00010111_1;
      patterns[24507] = 25'b01011111_10111001_00011000_1;
      patterns[24508] = 25'b01011111_10111010_00011001_1;
      patterns[24509] = 25'b01011111_10111011_00011010_1;
      patterns[24510] = 25'b01011111_10111100_00011011_1;
      patterns[24511] = 25'b01011111_10111101_00011100_1;
      patterns[24512] = 25'b01011111_10111110_00011101_1;
      patterns[24513] = 25'b01011111_10111111_00011110_1;
      patterns[24514] = 25'b01011111_11000000_00011111_1;
      patterns[24515] = 25'b01011111_11000001_00100000_1;
      patterns[24516] = 25'b01011111_11000010_00100001_1;
      patterns[24517] = 25'b01011111_11000011_00100010_1;
      patterns[24518] = 25'b01011111_11000100_00100011_1;
      patterns[24519] = 25'b01011111_11000101_00100100_1;
      patterns[24520] = 25'b01011111_11000110_00100101_1;
      patterns[24521] = 25'b01011111_11000111_00100110_1;
      patterns[24522] = 25'b01011111_11001000_00100111_1;
      patterns[24523] = 25'b01011111_11001001_00101000_1;
      patterns[24524] = 25'b01011111_11001010_00101001_1;
      patterns[24525] = 25'b01011111_11001011_00101010_1;
      patterns[24526] = 25'b01011111_11001100_00101011_1;
      patterns[24527] = 25'b01011111_11001101_00101100_1;
      patterns[24528] = 25'b01011111_11001110_00101101_1;
      patterns[24529] = 25'b01011111_11001111_00101110_1;
      patterns[24530] = 25'b01011111_11010000_00101111_1;
      patterns[24531] = 25'b01011111_11010001_00110000_1;
      patterns[24532] = 25'b01011111_11010010_00110001_1;
      patterns[24533] = 25'b01011111_11010011_00110010_1;
      patterns[24534] = 25'b01011111_11010100_00110011_1;
      patterns[24535] = 25'b01011111_11010101_00110100_1;
      patterns[24536] = 25'b01011111_11010110_00110101_1;
      patterns[24537] = 25'b01011111_11010111_00110110_1;
      patterns[24538] = 25'b01011111_11011000_00110111_1;
      patterns[24539] = 25'b01011111_11011001_00111000_1;
      patterns[24540] = 25'b01011111_11011010_00111001_1;
      patterns[24541] = 25'b01011111_11011011_00111010_1;
      patterns[24542] = 25'b01011111_11011100_00111011_1;
      patterns[24543] = 25'b01011111_11011101_00111100_1;
      patterns[24544] = 25'b01011111_11011110_00111101_1;
      patterns[24545] = 25'b01011111_11011111_00111110_1;
      patterns[24546] = 25'b01011111_11100000_00111111_1;
      patterns[24547] = 25'b01011111_11100001_01000000_1;
      patterns[24548] = 25'b01011111_11100010_01000001_1;
      patterns[24549] = 25'b01011111_11100011_01000010_1;
      patterns[24550] = 25'b01011111_11100100_01000011_1;
      patterns[24551] = 25'b01011111_11100101_01000100_1;
      patterns[24552] = 25'b01011111_11100110_01000101_1;
      patterns[24553] = 25'b01011111_11100111_01000110_1;
      patterns[24554] = 25'b01011111_11101000_01000111_1;
      patterns[24555] = 25'b01011111_11101001_01001000_1;
      patterns[24556] = 25'b01011111_11101010_01001001_1;
      patterns[24557] = 25'b01011111_11101011_01001010_1;
      patterns[24558] = 25'b01011111_11101100_01001011_1;
      patterns[24559] = 25'b01011111_11101101_01001100_1;
      patterns[24560] = 25'b01011111_11101110_01001101_1;
      patterns[24561] = 25'b01011111_11101111_01001110_1;
      patterns[24562] = 25'b01011111_11110000_01001111_1;
      patterns[24563] = 25'b01011111_11110001_01010000_1;
      patterns[24564] = 25'b01011111_11110010_01010001_1;
      patterns[24565] = 25'b01011111_11110011_01010010_1;
      patterns[24566] = 25'b01011111_11110100_01010011_1;
      patterns[24567] = 25'b01011111_11110101_01010100_1;
      patterns[24568] = 25'b01011111_11110110_01010101_1;
      patterns[24569] = 25'b01011111_11110111_01010110_1;
      patterns[24570] = 25'b01011111_11111000_01010111_1;
      patterns[24571] = 25'b01011111_11111001_01011000_1;
      patterns[24572] = 25'b01011111_11111010_01011001_1;
      patterns[24573] = 25'b01011111_11111011_01011010_1;
      patterns[24574] = 25'b01011111_11111100_01011011_1;
      patterns[24575] = 25'b01011111_11111101_01011100_1;
      patterns[24576] = 25'b01011111_11111110_01011101_1;
      patterns[24577] = 25'b01011111_11111111_01011110_1;
      patterns[24578] = 25'b01100000_00000000_01100000_0;
      patterns[24579] = 25'b01100000_00000001_01100001_0;
      patterns[24580] = 25'b01100000_00000010_01100010_0;
      patterns[24581] = 25'b01100000_00000011_01100011_0;
      patterns[24582] = 25'b01100000_00000100_01100100_0;
      patterns[24583] = 25'b01100000_00000101_01100101_0;
      patterns[24584] = 25'b01100000_00000110_01100110_0;
      patterns[24585] = 25'b01100000_00000111_01100111_0;
      patterns[24586] = 25'b01100000_00001000_01101000_0;
      patterns[24587] = 25'b01100000_00001001_01101001_0;
      patterns[24588] = 25'b01100000_00001010_01101010_0;
      patterns[24589] = 25'b01100000_00001011_01101011_0;
      patterns[24590] = 25'b01100000_00001100_01101100_0;
      patterns[24591] = 25'b01100000_00001101_01101101_0;
      patterns[24592] = 25'b01100000_00001110_01101110_0;
      patterns[24593] = 25'b01100000_00001111_01101111_0;
      patterns[24594] = 25'b01100000_00010000_01110000_0;
      patterns[24595] = 25'b01100000_00010001_01110001_0;
      patterns[24596] = 25'b01100000_00010010_01110010_0;
      patterns[24597] = 25'b01100000_00010011_01110011_0;
      patterns[24598] = 25'b01100000_00010100_01110100_0;
      patterns[24599] = 25'b01100000_00010101_01110101_0;
      patterns[24600] = 25'b01100000_00010110_01110110_0;
      patterns[24601] = 25'b01100000_00010111_01110111_0;
      patterns[24602] = 25'b01100000_00011000_01111000_0;
      patterns[24603] = 25'b01100000_00011001_01111001_0;
      patterns[24604] = 25'b01100000_00011010_01111010_0;
      patterns[24605] = 25'b01100000_00011011_01111011_0;
      patterns[24606] = 25'b01100000_00011100_01111100_0;
      patterns[24607] = 25'b01100000_00011101_01111101_0;
      patterns[24608] = 25'b01100000_00011110_01111110_0;
      patterns[24609] = 25'b01100000_00011111_01111111_0;
      patterns[24610] = 25'b01100000_00100000_10000000_0;
      patterns[24611] = 25'b01100000_00100001_10000001_0;
      patterns[24612] = 25'b01100000_00100010_10000010_0;
      patterns[24613] = 25'b01100000_00100011_10000011_0;
      patterns[24614] = 25'b01100000_00100100_10000100_0;
      patterns[24615] = 25'b01100000_00100101_10000101_0;
      patterns[24616] = 25'b01100000_00100110_10000110_0;
      patterns[24617] = 25'b01100000_00100111_10000111_0;
      patterns[24618] = 25'b01100000_00101000_10001000_0;
      patterns[24619] = 25'b01100000_00101001_10001001_0;
      patterns[24620] = 25'b01100000_00101010_10001010_0;
      patterns[24621] = 25'b01100000_00101011_10001011_0;
      patterns[24622] = 25'b01100000_00101100_10001100_0;
      patterns[24623] = 25'b01100000_00101101_10001101_0;
      patterns[24624] = 25'b01100000_00101110_10001110_0;
      patterns[24625] = 25'b01100000_00101111_10001111_0;
      patterns[24626] = 25'b01100000_00110000_10010000_0;
      patterns[24627] = 25'b01100000_00110001_10010001_0;
      patterns[24628] = 25'b01100000_00110010_10010010_0;
      patterns[24629] = 25'b01100000_00110011_10010011_0;
      patterns[24630] = 25'b01100000_00110100_10010100_0;
      patterns[24631] = 25'b01100000_00110101_10010101_0;
      patterns[24632] = 25'b01100000_00110110_10010110_0;
      patterns[24633] = 25'b01100000_00110111_10010111_0;
      patterns[24634] = 25'b01100000_00111000_10011000_0;
      patterns[24635] = 25'b01100000_00111001_10011001_0;
      patterns[24636] = 25'b01100000_00111010_10011010_0;
      patterns[24637] = 25'b01100000_00111011_10011011_0;
      patterns[24638] = 25'b01100000_00111100_10011100_0;
      patterns[24639] = 25'b01100000_00111101_10011101_0;
      patterns[24640] = 25'b01100000_00111110_10011110_0;
      patterns[24641] = 25'b01100000_00111111_10011111_0;
      patterns[24642] = 25'b01100000_01000000_10100000_0;
      patterns[24643] = 25'b01100000_01000001_10100001_0;
      patterns[24644] = 25'b01100000_01000010_10100010_0;
      patterns[24645] = 25'b01100000_01000011_10100011_0;
      patterns[24646] = 25'b01100000_01000100_10100100_0;
      patterns[24647] = 25'b01100000_01000101_10100101_0;
      patterns[24648] = 25'b01100000_01000110_10100110_0;
      patterns[24649] = 25'b01100000_01000111_10100111_0;
      patterns[24650] = 25'b01100000_01001000_10101000_0;
      patterns[24651] = 25'b01100000_01001001_10101001_0;
      patterns[24652] = 25'b01100000_01001010_10101010_0;
      patterns[24653] = 25'b01100000_01001011_10101011_0;
      patterns[24654] = 25'b01100000_01001100_10101100_0;
      patterns[24655] = 25'b01100000_01001101_10101101_0;
      patterns[24656] = 25'b01100000_01001110_10101110_0;
      patterns[24657] = 25'b01100000_01001111_10101111_0;
      patterns[24658] = 25'b01100000_01010000_10110000_0;
      patterns[24659] = 25'b01100000_01010001_10110001_0;
      patterns[24660] = 25'b01100000_01010010_10110010_0;
      patterns[24661] = 25'b01100000_01010011_10110011_0;
      patterns[24662] = 25'b01100000_01010100_10110100_0;
      patterns[24663] = 25'b01100000_01010101_10110101_0;
      patterns[24664] = 25'b01100000_01010110_10110110_0;
      patterns[24665] = 25'b01100000_01010111_10110111_0;
      patterns[24666] = 25'b01100000_01011000_10111000_0;
      patterns[24667] = 25'b01100000_01011001_10111001_0;
      patterns[24668] = 25'b01100000_01011010_10111010_0;
      patterns[24669] = 25'b01100000_01011011_10111011_0;
      patterns[24670] = 25'b01100000_01011100_10111100_0;
      patterns[24671] = 25'b01100000_01011101_10111101_0;
      patterns[24672] = 25'b01100000_01011110_10111110_0;
      patterns[24673] = 25'b01100000_01011111_10111111_0;
      patterns[24674] = 25'b01100000_01100000_11000000_0;
      patterns[24675] = 25'b01100000_01100001_11000001_0;
      patterns[24676] = 25'b01100000_01100010_11000010_0;
      patterns[24677] = 25'b01100000_01100011_11000011_0;
      patterns[24678] = 25'b01100000_01100100_11000100_0;
      patterns[24679] = 25'b01100000_01100101_11000101_0;
      patterns[24680] = 25'b01100000_01100110_11000110_0;
      patterns[24681] = 25'b01100000_01100111_11000111_0;
      patterns[24682] = 25'b01100000_01101000_11001000_0;
      patterns[24683] = 25'b01100000_01101001_11001001_0;
      patterns[24684] = 25'b01100000_01101010_11001010_0;
      patterns[24685] = 25'b01100000_01101011_11001011_0;
      patterns[24686] = 25'b01100000_01101100_11001100_0;
      patterns[24687] = 25'b01100000_01101101_11001101_0;
      patterns[24688] = 25'b01100000_01101110_11001110_0;
      patterns[24689] = 25'b01100000_01101111_11001111_0;
      patterns[24690] = 25'b01100000_01110000_11010000_0;
      patterns[24691] = 25'b01100000_01110001_11010001_0;
      patterns[24692] = 25'b01100000_01110010_11010010_0;
      patterns[24693] = 25'b01100000_01110011_11010011_0;
      patterns[24694] = 25'b01100000_01110100_11010100_0;
      patterns[24695] = 25'b01100000_01110101_11010101_0;
      patterns[24696] = 25'b01100000_01110110_11010110_0;
      patterns[24697] = 25'b01100000_01110111_11010111_0;
      patterns[24698] = 25'b01100000_01111000_11011000_0;
      patterns[24699] = 25'b01100000_01111001_11011001_0;
      patterns[24700] = 25'b01100000_01111010_11011010_0;
      patterns[24701] = 25'b01100000_01111011_11011011_0;
      patterns[24702] = 25'b01100000_01111100_11011100_0;
      patterns[24703] = 25'b01100000_01111101_11011101_0;
      patterns[24704] = 25'b01100000_01111110_11011110_0;
      patterns[24705] = 25'b01100000_01111111_11011111_0;
      patterns[24706] = 25'b01100000_10000000_11100000_0;
      patterns[24707] = 25'b01100000_10000001_11100001_0;
      patterns[24708] = 25'b01100000_10000010_11100010_0;
      patterns[24709] = 25'b01100000_10000011_11100011_0;
      patterns[24710] = 25'b01100000_10000100_11100100_0;
      patterns[24711] = 25'b01100000_10000101_11100101_0;
      patterns[24712] = 25'b01100000_10000110_11100110_0;
      patterns[24713] = 25'b01100000_10000111_11100111_0;
      patterns[24714] = 25'b01100000_10001000_11101000_0;
      patterns[24715] = 25'b01100000_10001001_11101001_0;
      patterns[24716] = 25'b01100000_10001010_11101010_0;
      patterns[24717] = 25'b01100000_10001011_11101011_0;
      patterns[24718] = 25'b01100000_10001100_11101100_0;
      patterns[24719] = 25'b01100000_10001101_11101101_0;
      patterns[24720] = 25'b01100000_10001110_11101110_0;
      patterns[24721] = 25'b01100000_10001111_11101111_0;
      patterns[24722] = 25'b01100000_10010000_11110000_0;
      patterns[24723] = 25'b01100000_10010001_11110001_0;
      patterns[24724] = 25'b01100000_10010010_11110010_0;
      patterns[24725] = 25'b01100000_10010011_11110011_0;
      patterns[24726] = 25'b01100000_10010100_11110100_0;
      patterns[24727] = 25'b01100000_10010101_11110101_0;
      patterns[24728] = 25'b01100000_10010110_11110110_0;
      patterns[24729] = 25'b01100000_10010111_11110111_0;
      patterns[24730] = 25'b01100000_10011000_11111000_0;
      patterns[24731] = 25'b01100000_10011001_11111001_0;
      patterns[24732] = 25'b01100000_10011010_11111010_0;
      patterns[24733] = 25'b01100000_10011011_11111011_0;
      patterns[24734] = 25'b01100000_10011100_11111100_0;
      patterns[24735] = 25'b01100000_10011101_11111101_0;
      patterns[24736] = 25'b01100000_10011110_11111110_0;
      patterns[24737] = 25'b01100000_10011111_11111111_0;
      patterns[24738] = 25'b01100000_10100000_00000000_1;
      patterns[24739] = 25'b01100000_10100001_00000001_1;
      patterns[24740] = 25'b01100000_10100010_00000010_1;
      patterns[24741] = 25'b01100000_10100011_00000011_1;
      patterns[24742] = 25'b01100000_10100100_00000100_1;
      patterns[24743] = 25'b01100000_10100101_00000101_1;
      patterns[24744] = 25'b01100000_10100110_00000110_1;
      patterns[24745] = 25'b01100000_10100111_00000111_1;
      patterns[24746] = 25'b01100000_10101000_00001000_1;
      patterns[24747] = 25'b01100000_10101001_00001001_1;
      patterns[24748] = 25'b01100000_10101010_00001010_1;
      patterns[24749] = 25'b01100000_10101011_00001011_1;
      patterns[24750] = 25'b01100000_10101100_00001100_1;
      patterns[24751] = 25'b01100000_10101101_00001101_1;
      patterns[24752] = 25'b01100000_10101110_00001110_1;
      patterns[24753] = 25'b01100000_10101111_00001111_1;
      patterns[24754] = 25'b01100000_10110000_00010000_1;
      patterns[24755] = 25'b01100000_10110001_00010001_1;
      patterns[24756] = 25'b01100000_10110010_00010010_1;
      patterns[24757] = 25'b01100000_10110011_00010011_1;
      patterns[24758] = 25'b01100000_10110100_00010100_1;
      patterns[24759] = 25'b01100000_10110101_00010101_1;
      patterns[24760] = 25'b01100000_10110110_00010110_1;
      patterns[24761] = 25'b01100000_10110111_00010111_1;
      patterns[24762] = 25'b01100000_10111000_00011000_1;
      patterns[24763] = 25'b01100000_10111001_00011001_1;
      patterns[24764] = 25'b01100000_10111010_00011010_1;
      patterns[24765] = 25'b01100000_10111011_00011011_1;
      patterns[24766] = 25'b01100000_10111100_00011100_1;
      patterns[24767] = 25'b01100000_10111101_00011101_1;
      patterns[24768] = 25'b01100000_10111110_00011110_1;
      patterns[24769] = 25'b01100000_10111111_00011111_1;
      patterns[24770] = 25'b01100000_11000000_00100000_1;
      patterns[24771] = 25'b01100000_11000001_00100001_1;
      patterns[24772] = 25'b01100000_11000010_00100010_1;
      patterns[24773] = 25'b01100000_11000011_00100011_1;
      patterns[24774] = 25'b01100000_11000100_00100100_1;
      patterns[24775] = 25'b01100000_11000101_00100101_1;
      patterns[24776] = 25'b01100000_11000110_00100110_1;
      patterns[24777] = 25'b01100000_11000111_00100111_1;
      patterns[24778] = 25'b01100000_11001000_00101000_1;
      patterns[24779] = 25'b01100000_11001001_00101001_1;
      patterns[24780] = 25'b01100000_11001010_00101010_1;
      patterns[24781] = 25'b01100000_11001011_00101011_1;
      patterns[24782] = 25'b01100000_11001100_00101100_1;
      patterns[24783] = 25'b01100000_11001101_00101101_1;
      patterns[24784] = 25'b01100000_11001110_00101110_1;
      patterns[24785] = 25'b01100000_11001111_00101111_1;
      patterns[24786] = 25'b01100000_11010000_00110000_1;
      patterns[24787] = 25'b01100000_11010001_00110001_1;
      patterns[24788] = 25'b01100000_11010010_00110010_1;
      patterns[24789] = 25'b01100000_11010011_00110011_1;
      patterns[24790] = 25'b01100000_11010100_00110100_1;
      patterns[24791] = 25'b01100000_11010101_00110101_1;
      patterns[24792] = 25'b01100000_11010110_00110110_1;
      patterns[24793] = 25'b01100000_11010111_00110111_1;
      patterns[24794] = 25'b01100000_11011000_00111000_1;
      patterns[24795] = 25'b01100000_11011001_00111001_1;
      patterns[24796] = 25'b01100000_11011010_00111010_1;
      patterns[24797] = 25'b01100000_11011011_00111011_1;
      patterns[24798] = 25'b01100000_11011100_00111100_1;
      patterns[24799] = 25'b01100000_11011101_00111101_1;
      patterns[24800] = 25'b01100000_11011110_00111110_1;
      patterns[24801] = 25'b01100000_11011111_00111111_1;
      patterns[24802] = 25'b01100000_11100000_01000000_1;
      patterns[24803] = 25'b01100000_11100001_01000001_1;
      patterns[24804] = 25'b01100000_11100010_01000010_1;
      patterns[24805] = 25'b01100000_11100011_01000011_1;
      patterns[24806] = 25'b01100000_11100100_01000100_1;
      patterns[24807] = 25'b01100000_11100101_01000101_1;
      patterns[24808] = 25'b01100000_11100110_01000110_1;
      patterns[24809] = 25'b01100000_11100111_01000111_1;
      patterns[24810] = 25'b01100000_11101000_01001000_1;
      patterns[24811] = 25'b01100000_11101001_01001001_1;
      patterns[24812] = 25'b01100000_11101010_01001010_1;
      patterns[24813] = 25'b01100000_11101011_01001011_1;
      patterns[24814] = 25'b01100000_11101100_01001100_1;
      patterns[24815] = 25'b01100000_11101101_01001101_1;
      patterns[24816] = 25'b01100000_11101110_01001110_1;
      patterns[24817] = 25'b01100000_11101111_01001111_1;
      patterns[24818] = 25'b01100000_11110000_01010000_1;
      patterns[24819] = 25'b01100000_11110001_01010001_1;
      patterns[24820] = 25'b01100000_11110010_01010010_1;
      patterns[24821] = 25'b01100000_11110011_01010011_1;
      patterns[24822] = 25'b01100000_11110100_01010100_1;
      patterns[24823] = 25'b01100000_11110101_01010101_1;
      patterns[24824] = 25'b01100000_11110110_01010110_1;
      patterns[24825] = 25'b01100000_11110111_01010111_1;
      patterns[24826] = 25'b01100000_11111000_01011000_1;
      patterns[24827] = 25'b01100000_11111001_01011001_1;
      patterns[24828] = 25'b01100000_11111010_01011010_1;
      patterns[24829] = 25'b01100000_11111011_01011011_1;
      patterns[24830] = 25'b01100000_11111100_01011100_1;
      patterns[24831] = 25'b01100000_11111101_01011101_1;
      patterns[24832] = 25'b01100000_11111110_01011110_1;
      patterns[24833] = 25'b01100000_11111111_01011111_1;
      patterns[24834] = 25'b01100001_00000000_01100001_0;
      patterns[24835] = 25'b01100001_00000001_01100010_0;
      patterns[24836] = 25'b01100001_00000010_01100011_0;
      patterns[24837] = 25'b01100001_00000011_01100100_0;
      patterns[24838] = 25'b01100001_00000100_01100101_0;
      patterns[24839] = 25'b01100001_00000101_01100110_0;
      patterns[24840] = 25'b01100001_00000110_01100111_0;
      patterns[24841] = 25'b01100001_00000111_01101000_0;
      patterns[24842] = 25'b01100001_00001000_01101001_0;
      patterns[24843] = 25'b01100001_00001001_01101010_0;
      patterns[24844] = 25'b01100001_00001010_01101011_0;
      patterns[24845] = 25'b01100001_00001011_01101100_0;
      patterns[24846] = 25'b01100001_00001100_01101101_0;
      patterns[24847] = 25'b01100001_00001101_01101110_0;
      patterns[24848] = 25'b01100001_00001110_01101111_0;
      patterns[24849] = 25'b01100001_00001111_01110000_0;
      patterns[24850] = 25'b01100001_00010000_01110001_0;
      patterns[24851] = 25'b01100001_00010001_01110010_0;
      patterns[24852] = 25'b01100001_00010010_01110011_0;
      patterns[24853] = 25'b01100001_00010011_01110100_0;
      patterns[24854] = 25'b01100001_00010100_01110101_0;
      patterns[24855] = 25'b01100001_00010101_01110110_0;
      patterns[24856] = 25'b01100001_00010110_01110111_0;
      patterns[24857] = 25'b01100001_00010111_01111000_0;
      patterns[24858] = 25'b01100001_00011000_01111001_0;
      patterns[24859] = 25'b01100001_00011001_01111010_0;
      patterns[24860] = 25'b01100001_00011010_01111011_0;
      patterns[24861] = 25'b01100001_00011011_01111100_0;
      patterns[24862] = 25'b01100001_00011100_01111101_0;
      patterns[24863] = 25'b01100001_00011101_01111110_0;
      patterns[24864] = 25'b01100001_00011110_01111111_0;
      patterns[24865] = 25'b01100001_00011111_10000000_0;
      patterns[24866] = 25'b01100001_00100000_10000001_0;
      patterns[24867] = 25'b01100001_00100001_10000010_0;
      patterns[24868] = 25'b01100001_00100010_10000011_0;
      patterns[24869] = 25'b01100001_00100011_10000100_0;
      patterns[24870] = 25'b01100001_00100100_10000101_0;
      patterns[24871] = 25'b01100001_00100101_10000110_0;
      patterns[24872] = 25'b01100001_00100110_10000111_0;
      patterns[24873] = 25'b01100001_00100111_10001000_0;
      patterns[24874] = 25'b01100001_00101000_10001001_0;
      patterns[24875] = 25'b01100001_00101001_10001010_0;
      patterns[24876] = 25'b01100001_00101010_10001011_0;
      patterns[24877] = 25'b01100001_00101011_10001100_0;
      patterns[24878] = 25'b01100001_00101100_10001101_0;
      patterns[24879] = 25'b01100001_00101101_10001110_0;
      patterns[24880] = 25'b01100001_00101110_10001111_0;
      patterns[24881] = 25'b01100001_00101111_10010000_0;
      patterns[24882] = 25'b01100001_00110000_10010001_0;
      patterns[24883] = 25'b01100001_00110001_10010010_0;
      patterns[24884] = 25'b01100001_00110010_10010011_0;
      patterns[24885] = 25'b01100001_00110011_10010100_0;
      patterns[24886] = 25'b01100001_00110100_10010101_0;
      patterns[24887] = 25'b01100001_00110101_10010110_0;
      patterns[24888] = 25'b01100001_00110110_10010111_0;
      patterns[24889] = 25'b01100001_00110111_10011000_0;
      patterns[24890] = 25'b01100001_00111000_10011001_0;
      patterns[24891] = 25'b01100001_00111001_10011010_0;
      patterns[24892] = 25'b01100001_00111010_10011011_0;
      patterns[24893] = 25'b01100001_00111011_10011100_0;
      patterns[24894] = 25'b01100001_00111100_10011101_0;
      patterns[24895] = 25'b01100001_00111101_10011110_0;
      patterns[24896] = 25'b01100001_00111110_10011111_0;
      patterns[24897] = 25'b01100001_00111111_10100000_0;
      patterns[24898] = 25'b01100001_01000000_10100001_0;
      patterns[24899] = 25'b01100001_01000001_10100010_0;
      patterns[24900] = 25'b01100001_01000010_10100011_0;
      patterns[24901] = 25'b01100001_01000011_10100100_0;
      patterns[24902] = 25'b01100001_01000100_10100101_0;
      patterns[24903] = 25'b01100001_01000101_10100110_0;
      patterns[24904] = 25'b01100001_01000110_10100111_0;
      patterns[24905] = 25'b01100001_01000111_10101000_0;
      patterns[24906] = 25'b01100001_01001000_10101001_0;
      patterns[24907] = 25'b01100001_01001001_10101010_0;
      patterns[24908] = 25'b01100001_01001010_10101011_0;
      patterns[24909] = 25'b01100001_01001011_10101100_0;
      patterns[24910] = 25'b01100001_01001100_10101101_0;
      patterns[24911] = 25'b01100001_01001101_10101110_0;
      patterns[24912] = 25'b01100001_01001110_10101111_0;
      patterns[24913] = 25'b01100001_01001111_10110000_0;
      patterns[24914] = 25'b01100001_01010000_10110001_0;
      patterns[24915] = 25'b01100001_01010001_10110010_0;
      patterns[24916] = 25'b01100001_01010010_10110011_0;
      patterns[24917] = 25'b01100001_01010011_10110100_0;
      patterns[24918] = 25'b01100001_01010100_10110101_0;
      patterns[24919] = 25'b01100001_01010101_10110110_0;
      patterns[24920] = 25'b01100001_01010110_10110111_0;
      patterns[24921] = 25'b01100001_01010111_10111000_0;
      patterns[24922] = 25'b01100001_01011000_10111001_0;
      patterns[24923] = 25'b01100001_01011001_10111010_0;
      patterns[24924] = 25'b01100001_01011010_10111011_0;
      patterns[24925] = 25'b01100001_01011011_10111100_0;
      patterns[24926] = 25'b01100001_01011100_10111101_0;
      patterns[24927] = 25'b01100001_01011101_10111110_0;
      patterns[24928] = 25'b01100001_01011110_10111111_0;
      patterns[24929] = 25'b01100001_01011111_11000000_0;
      patterns[24930] = 25'b01100001_01100000_11000001_0;
      patterns[24931] = 25'b01100001_01100001_11000010_0;
      patterns[24932] = 25'b01100001_01100010_11000011_0;
      patterns[24933] = 25'b01100001_01100011_11000100_0;
      patterns[24934] = 25'b01100001_01100100_11000101_0;
      patterns[24935] = 25'b01100001_01100101_11000110_0;
      patterns[24936] = 25'b01100001_01100110_11000111_0;
      patterns[24937] = 25'b01100001_01100111_11001000_0;
      patterns[24938] = 25'b01100001_01101000_11001001_0;
      patterns[24939] = 25'b01100001_01101001_11001010_0;
      patterns[24940] = 25'b01100001_01101010_11001011_0;
      patterns[24941] = 25'b01100001_01101011_11001100_0;
      patterns[24942] = 25'b01100001_01101100_11001101_0;
      patterns[24943] = 25'b01100001_01101101_11001110_0;
      patterns[24944] = 25'b01100001_01101110_11001111_0;
      patterns[24945] = 25'b01100001_01101111_11010000_0;
      patterns[24946] = 25'b01100001_01110000_11010001_0;
      patterns[24947] = 25'b01100001_01110001_11010010_0;
      patterns[24948] = 25'b01100001_01110010_11010011_0;
      patterns[24949] = 25'b01100001_01110011_11010100_0;
      patterns[24950] = 25'b01100001_01110100_11010101_0;
      patterns[24951] = 25'b01100001_01110101_11010110_0;
      patterns[24952] = 25'b01100001_01110110_11010111_0;
      patterns[24953] = 25'b01100001_01110111_11011000_0;
      patterns[24954] = 25'b01100001_01111000_11011001_0;
      patterns[24955] = 25'b01100001_01111001_11011010_0;
      patterns[24956] = 25'b01100001_01111010_11011011_0;
      patterns[24957] = 25'b01100001_01111011_11011100_0;
      patterns[24958] = 25'b01100001_01111100_11011101_0;
      patterns[24959] = 25'b01100001_01111101_11011110_0;
      patterns[24960] = 25'b01100001_01111110_11011111_0;
      patterns[24961] = 25'b01100001_01111111_11100000_0;
      patterns[24962] = 25'b01100001_10000000_11100001_0;
      patterns[24963] = 25'b01100001_10000001_11100010_0;
      patterns[24964] = 25'b01100001_10000010_11100011_0;
      patterns[24965] = 25'b01100001_10000011_11100100_0;
      patterns[24966] = 25'b01100001_10000100_11100101_0;
      patterns[24967] = 25'b01100001_10000101_11100110_0;
      patterns[24968] = 25'b01100001_10000110_11100111_0;
      patterns[24969] = 25'b01100001_10000111_11101000_0;
      patterns[24970] = 25'b01100001_10001000_11101001_0;
      patterns[24971] = 25'b01100001_10001001_11101010_0;
      patterns[24972] = 25'b01100001_10001010_11101011_0;
      patterns[24973] = 25'b01100001_10001011_11101100_0;
      patterns[24974] = 25'b01100001_10001100_11101101_0;
      patterns[24975] = 25'b01100001_10001101_11101110_0;
      patterns[24976] = 25'b01100001_10001110_11101111_0;
      patterns[24977] = 25'b01100001_10001111_11110000_0;
      patterns[24978] = 25'b01100001_10010000_11110001_0;
      patterns[24979] = 25'b01100001_10010001_11110010_0;
      patterns[24980] = 25'b01100001_10010010_11110011_0;
      patterns[24981] = 25'b01100001_10010011_11110100_0;
      patterns[24982] = 25'b01100001_10010100_11110101_0;
      patterns[24983] = 25'b01100001_10010101_11110110_0;
      patterns[24984] = 25'b01100001_10010110_11110111_0;
      patterns[24985] = 25'b01100001_10010111_11111000_0;
      patterns[24986] = 25'b01100001_10011000_11111001_0;
      patterns[24987] = 25'b01100001_10011001_11111010_0;
      patterns[24988] = 25'b01100001_10011010_11111011_0;
      patterns[24989] = 25'b01100001_10011011_11111100_0;
      patterns[24990] = 25'b01100001_10011100_11111101_0;
      patterns[24991] = 25'b01100001_10011101_11111110_0;
      patterns[24992] = 25'b01100001_10011110_11111111_0;
      patterns[24993] = 25'b01100001_10011111_00000000_1;
      patterns[24994] = 25'b01100001_10100000_00000001_1;
      patterns[24995] = 25'b01100001_10100001_00000010_1;
      patterns[24996] = 25'b01100001_10100010_00000011_1;
      patterns[24997] = 25'b01100001_10100011_00000100_1;
      patterns[24998] = 25'b01100001_10100100_00000101_1;
      patterns[24999] = 25'b01100001_10100101_00000110_1;
      patterns[25000] = 25'b01100001_10100110_00000111_1;
      patterns[25001] = 25'b01100001_10100111_00001000_1;
      patterns[25002] = 25'b01100001_10101000_00001001_1;
      patterns[25003] = 25'b01100001_10101001_00001010_1;
      patterns[25004] = 25'b01100001_10101010_00001011_1;
      patterns[25005] = 25'b01100001_10101011_00001100_1;
      patterns[25006] = 25'b01100001_10101100_00001101_1;
      patterns[25007] = 25'b01100001_10101101_00001110_1;
      patterns[25008] = 25'b01100001_10101110_00001111_1;
      patterns[25009] = 25'b01100001_10101111_00010000_1;
      patterns[25010] = 25'b01100001_10110000_00010001_1;
      patterns[25011] = 25'b01100001_10110001_00010010_1;
      patterns[25012] = 25'b01100001_10110010_00010011_1;
      patterns[25013] = 25'b01100001_10110011_00010100_1;
      patterns[25014] = 25'b01100001_10110100_00010101_1;
      patterns[25015] = 25'b01100001_10110101_00010110_1;
      patterns[25016] = 25'b01100001_10110110_00010111_1;
      patterns[25017] = 25'b01100001_10110111_00011000_1;
      patterns[25018] = 25'b01100001_10111000_00011001_1;
      patterns[25019] = 25'b01100001_10111001_00011010_1;
      patterns[25020] = 25'b01100001_10111010_00011011_1;
      patterns[25021] = 25'b01100001_10111011_00011100_1;
      patterns[25022] = 25'b01100001_10111100_00011101_1;
      patterns[25023] = 25'b01100001_10111101_00011110_1;
      patterns[25024] = 25'b01100001_10111110_00011111_1;
      patterns[25025] = 25'b01100001_10111111_00100000_1;
      patterns[25026] = 25'b01100001_11000000_00100001_1;
      patterns[25027] = 25'b01100001_11000001_00100010_1;
      patterns[25028] = 25'b01100001_11000010_00100011_1;
      patterns[25029] = 25'b01100001_11000011_00100100_1;
      patterns[25030] = 25'b01100001_11000100_00100101_1;
      patterns[25031] = 25'b01100001_11000101_00100110_1;
      patterns[25032] = 25'b01100001_11000110_00100111_1;
      patterns[25033] = 25'b01100001_11000111_00101000_1;
      patterns[25034] = 25'b01100001_11001000_00101001_1;
      patterns[25035] = 25'b01100001_11001001_00101010_1;
      patterns[25036] = 25'b01100001_11001010_00101011_1;
      patterns[25037] = 25'b01100001_11001011_00101100_1;
      patterns[25038] = 25'b01100001_11001100_00101101_1;
      patterns[25039] = 25'b01100001_11001101_00101110_1;
      patterns[25040] = 25'b01100001_11001110_00101111_1;
      patterns[25041] = 25'b01100001_11001111_00110000_1;
      patterns[25042] = 25'b01100001_11010000_00110001_1;
      patterns[25043] = 25'b01100001_11010001_00110010_1;
      patterns[25044] = 25'b01100001_11010010_00110011_1;
      patterns[25045] = 25'b01100001_11010011_00110100_1;
      patterns[25046] = 25'b01100001_11010100_00110101_1;
      patterns[25047] = 25'b01100001_11010101_00110110_1;
      patterns[25048] = 25'b01100001_11010110_00110111_1;
      patterns[25049] = 25'b01100001_11010111_00111000_1;
      patterns[25050] = 25'b01100001_11011000_00111001_1;
      patterns[25051] = 25'b01100001_11011001_00111010_1;
      patterns[25052] = 25'b01100001_11011010_00111011_1;
      patterns[25053] = 25'b01100001_11011011_00111100_1;
      patterns[25054] = 25'b01100001_11011100_00111101_1;
      patterns[25055] = 25'b01100001_11011101_00111110_1;
      patterns[25056] = 25'b01100001_11011110_00111111_1;
      patterns[25057] = 25'b01100001_11011111_01000000_1;
      patterns[25058] = 25'b01100001_11100000_01000001_1;
      patterns[25059] = 25'b01100001_11100001_01000010_1;
      patterns[25060] = 25'b01100001_11100010_01000011_1;
      patterns[25061] = 25'b01100001_11100011_01000100_1;
      patterns[25062] = 25'b01100001_11100100_01000101_1;
      patterns[25063] = 25'b01100001_11100101_01000110_1;
      patterns[25064] = 25'b01100001_11100110_01000111_1;
      patterns[25065] = 25'b01100001_11100111_01001000_1;
      patterns[25066] = 25'b01100001_11101000_01001001_1;
      patterns[25067] = 25'b01100001_11101001_01001010_1;
      patterns[25068] = 25'b01100001_11101010_01001011_1;
      patterns[25069] = 25'b01100001_11101011_01001100_1;
      patterns[25070] = 25'b01100001_11101100_01001101_1;
      patterns[25071] = 25'b01100001_11101101_01001110_1;
      patterns[25072] = 25'b01100001_11101110_01001111_1;
      patterns[25073] = 25'b01100001_11101111_01010000_1;
      patterns[25074] = 25'b01100001_11110000_01010001_1;
      patterns[25075] = 25'b01100001_11110001_01010010_1;
      patterns[25076] = 25'b01100001_11110010_01010011_1;
      patterns[25077] = 25'b01100001_11110011_01010100_1;
      patterns[25078] = 25'b01100001_11110100_01010101_1;
      patterns[25079] = 25'b01100001_11110101_01010110_1;
      patterns[25080] = 25'b01100001_11110110_01010111_1;
      patterns[25081] = 25'b01100001_11110111_01011000_1;
      patterns[25082] = 25'b01100001_11111000_01011001_1;
      patterns[25083] = 25'b01100001_11111001_01011010_1;
      patterns[25084] = 25'b01100001_11111010_01011011_1;
      patterns[25085] = 25'b01100001_11111011_01011100_1;
      patterns[25086] = 25'b01100001_11111100_01011101_1;
      patterns[25087] = 25'b01100001_11111101_01011110_1;
      patterns[25088] = 25'b01100001_11111110_01011111_1;
      patterns[25089] = 25'b01100001_11111111_01100000_1;
      patterns[25090] = 25'b01100010_00000000_01100010_0;
      patterns[25091] = 25'b01100010_00000001_01100011_0;
      patterns[25092] = 25'b01100010_00000010_01100100_0;
      patterns[25093] = 25'b01100010_00000011_01100101_0;
      patterns[25094] = 25'b01100010_00000100_01100110_0;
      patterns[25095] = 25'b01100010_00000101_01100111_0;
      patterns[25096] = 25'b01100010_00000110_01101000_0;
      patterns[25097] = 25'b01100010_00000111_01101001_0;
      patterns[25098] = 25'b01100010_00001000_01101010_0;
      patterns[25099] = 25'b01100010_00001001_01101011_0;
      patterns[25100] = 25'b01100010_00001010_01101100_0;
      patterns[25101] = 25'b01100010_00001011_01101101_0;
      patterns[25102] = 25'b01100010_00001100_01101110_0;
      patterns[25103] = 25'b01100010_00001101_01101111_0;
      patterns[25104] = 25'b01100010_00001110_01110000_0;
      patterns[25105] = 25'b01100010_00001111_01110001_0;
      patterns[25106] = 25'b01100010_00010000_01110010_0;
      patterns[25107] = 25'b01100010_00010001_01110011_0;
      patterns[25108] = 25'b01100010_00010010_01110100_0;
      patterns[25109] = 25'b01100010_00010011_01110101_0;
      patterns[25110] = 25'b01100010_00010100_01110110_0;
      patterns[25111] = 25'b01100010_00010101_01110111_0;
      patterns[25112] = 25'b01100010_00010110_01111000_0;
      patterns[25113] = 25'b01100010_00010111_01111001_0;
      patterns[25114] = 25'b01100010_00011000_01111010_0;
      patterns[25115] = 25'b01100010_00011001_01111011_0;
      patterns[25116] = 25'b01100010_00011010_01111100_0;
      patterns[25117] = 25'b01100010_00011011_01111101_0;
      patterns[25118] = 25'b01100010_00011100_01111110_0;
      patterns[25119] = 25'b01100010_00011101_01111111_0;
      patterns[25120] = 25'b01100010_00011110_10000000_0;
      patterns[25121] = 25'b01100010_00011111_10000001_0;
      patterns[25122] = 25'b01100010_00100000_10000010_0;
      patterns[25123] = 25'b01100010_00100001_10000011_0;
      patterns[25124] = 25'b01100010_00100010_10000100_0;
      patterns[25125] = 25'b01100010_00100011_10000101_0;
      patterns[25126] = 25'b01100010_00100100_10000110_0;
      patterns[25127] = 25'b01100010_00100101_10000111_0;
      patterns[25128] = 25'b01100010_00100110_10001000_0;
      patterns[25129] = 25'b01100010_00100111_10001001_0;
      patterns[25130] = 25'b01100010_00101000_10001010_0;
      patterns[25131] = 25'b01100010_00101001_10001011_0;
      patterns[25132] = 25'b01100010_00101010_10001100_0;
      patterns[25133] = 25'b01100010_00101011_10001101_0;
      patterns[25134] = 25'b01100010_00101100_10001110_0;
      patterns[25135] = 25'b01100010_00101101_10001111_0;
      patterns[25136] = 25'b01100010_00101110_10010000_0;
      patterns[25137] = 25'b01100010_00101111_10010001_0;
      patterns[25138] = 25'b01100010_00110000_10010010_0;
      patterns[25139] = 25'b01100010_00110001_10010011_0;
      patterns[25140] = 25'b01100010_00110010_10010100_0;
      patterns[25141] = 25'b01100010_00110011_10010101_0;
      patterns[25142] = 25'b01100010_00110100_10010110_0;
      patterns[25143] = 25'b01100010_00110101_10010111_0;
      patterns[25144] = 25'b01100010_00110110_10011000_0;
      patterns[25145] = 25'b01100010_00110111_10011001_0;
      patterns[25146] = 25'b01100010_00111000_10011010_0;
      patterns[25147] = 25'b01100010_00111001_10011011_0;
      patterns[25148] = 25'b01100010_00111010_10011100_0;
      patterns[25149] = 25'b01100010_00111011_10011101_0;
      patterns[25150] = 25'b01100010_00111100_10011110_0;
      patterns[25151] = 25'b01100010_00111101_10011111_0;
      patterns[25152] = 25'b01100010_00111110_10100000_0;
      patterns[25153] = 25'b01100010_00111111_10100001_0;
      patterns[25154] = 25'b01100010_01000000_10100010_0;
      patterns[25155] = 25'b01100010_01000001_10100011_0;
      patterns[25156] = 25'b01100010_01000010_10100100_0;
      patterns[25157] = 25'b01100010_01000011_10100101_0;
      patterns[25158] = 25'b01100010_01000100_10100110_0;
      patterns[25159] = 25'b01100010_01000101_10100111_0;
      patterns[25160] = 25'b01100010_01000110_10101000_0;
      patterns[25161] = 25'b01100010_01000111_10101001_0;
      patterns[25162] = 25'b01100010_01001000_10101010_0;
      patterns[25163] = 25'b01100010_01001001_10101011_0;
      patterns[25164] = 25'b01100010_01001010_10101100_0;
      patterns[25165] = 25'b01100010_01001011_10101101_0;
      patterns[25166] = 25'b01100010_01001100_10101110_0;
      patterns[25167] = 25'b01100010_01001101_10101111_0;
      patterns[25168] = 25'b01100010_01001110_10110000_0;
      patterns[25169] = 25'b01100010_01001111_10110001_0;
      patterns[25170] = 25'b01100010_01010000_10110010_0;
      patterns[25171] = 25'b01100010_01010001_10110011_0;
      patterns[25172] = 25'b01100010_01010010_10110100_0;
      patterns[25173] = 25'b01100010_01010011_10110101_0;
      patterns[25174] = 25'b01100010_01010100_10110110_0;
      patterns[25175] = 25'b01100010_01010101_10110111_0;
      patterns[25176] = 25'b01100010_01010110_10111000_0;
      patterns[25177] = 25'b01100010_01010111_10111001_0;
      patterns[25178] = 25'b01100010_01011000_10111010_0;
      patterns[25179] = 25'b01100010_01011001_10111011_0;
      patterns[25180] = 25'b01100010_01011010_10111100_0;
      patterns[25181] = 25'b01100010_01011011_10111101_0;
      patterns[25182] = 25'b01100010_01011100_10111110_0;
      patterns[25183] = 25'b01100010_01011101_10111111_0;
      patterns[25184] = 25'b01100010_01011110_11000000_0;
      patterns[25185] = 25'b01100010_01011111_11000001_0;
      patterns[25186] = 25'b01100010_01100000_11000010_0;
      patterns[25187] = 25'b01100010_01100001_11000011_0;
      patterns[25188] = 25'b01100010_01100010_11000100_0;
      patterns[25189] = 25'b01100010_01100011_11000101_0;
      patterns[25190] = 25'b01100010_01100100_11000110_0;
      patterns[25191] = 25'b01100010_01100101_11000111_0;
      patterns[25192] = 25'b01100010_01100110_11001000_0;
      patterns[25193] = 25'b01100010_01100111_11001001_0;
      patterns[25194] = 25'b01100010_01101000_11001010_0;
      patterns[25195] = 25'b01100010_01101001_11001011_0;
      patterns[25196] = 25'b01100010_01101010_11001100_0;
      patterns[25197] = 25'b01100010_01101011_11001101_0;
      patterns[25198] = 25'b01100010_01101100_11001110_0;
      patterns[25199] = 25'b01100010_01101101_11001111_0;
      patterns[25200] = 25'b01100010_01101110_11010000_0;
      patterns[25201] = 25'b01100010_01101111_11010001_0;
      patterns[25202] = 25'b01100010_01110000_11010010_0;
      patterns[25203] = 25'b01100010_01110001_11010011_0;
      patterns[25204] = 25'b01100010_01110010_11010100_0;
      patterns[25205] = 25'b01100010_01110011_11010101_0;
      patterns[25206] = 25'b01100010_01110100_11010110_0;
      patterns[25207] = 25'b01100010_01110101_11010111_0;
      patterns[25208] = 25'b01100010_01110110_11011000_0;
      patterns[25209] = 25'b01100010_01110111_11011001_0;
      patterns[25210] = 25'b01100010_01111000_11011010_0;
      patterns[25211] = 25'b01100010_01111001_11011011_0;
      patterns[25212] = 25'b01100010_01111010_11011100_0;
      patterns[25213] = 25'b01100010_01111011_11011101_0;
      patterns[25214] = 25'b01100010_01111100_11011110_0;
      patterns[25215] = 25'b01100010_01111101_11011111_0;
      patterns[25216] = 25'b01100010_01111110_11100000_0;
      patterns[25217] = 25'b01100010_01111111_11100001_0;
      patterns[25218] = 25'b01100010_10000000_11100010_0;
      patterns[25219] = 25'b01100010_10000001_11100011_0;
      patterns[25220] = 25'b01100010_10000010_11100100_0;
      patterns[25221] = 25'b01100010_10000011_11100101_0;
      patterns[25222] = 25'b01100010_10000100_11100110_0;
      patterns[25223] = 25'b01100010_10000101_11100111_0;
      patterns[25224] = 25'b01100010_10000110_11101000_0;
      patterns[25225] = 25'b01100010_10000111_11101001_0;
      patterns[25226] = 25'b01100010_10001000_11101010_0;
      patterns[25227] = 25'b01100010_10001001_11101011_0;
      patterns[25228] = 25'b01100010_10001010_11101100_0;
      patterns[25229] = 25'b01100010_10001011_11101101_0;
      patterns[25230] = 25'b01100010_10001100_11101110_0;
      patterns[25231] = 25'b01100010_10001101_11101111_0;
      patterns[25232] = 25'b01100010_10001110_11110000_0;
      patterns[25233] = 25'b01100010_10001111_11110001_0;
      patterns[25234] = 25'b01100010_10010000_11110010_0;
      patterns[25235] = 25'b01100010_10010001_11110011_0;
      patterns[25236] = 25'b01100010_10010010_11110100_0;
      patterns[25237] = 25'b01100010_10010011_11110101_0;
      patterns[25238] = 25'b01100010_10010100_11110110_0;
      patterns[25239] = 25'b01100010_10010101_11110111_0;
      patterns[25240] = 25'b01100010_10010110_11111000_0;
      patterns[25241] = 25'b01100010_10010111_11111001_0;
      patterns[25242] = 25'b01100010_10011000_11111010_0;
      patterns[25243] = 25'b01100010_10011001_11111011_0;
      patterns[25244] = 25'b01100010_10011010_11111100_0;
      patterns[25245] = 25'b01100010_10011011_11111101_0;
      patterns[25246] = 25'b01100010_10011100_11111110_0;
      patterns[25247] = 25'b01100010_10011101_11111111_0;
      patterns[25248] = 25'b01100010_10011110_00000000_1;
      patterns[25249] = 25'b01100010_10011111_00000001_1;
      patterns[25250] = 25'b01100010_10100000_00000010_1;
      patterns[25251] = 25'b01100010_10100001_00000011_1;
      patterns[25252] = 25'b01100010_10100010_00000100_1;
      patterns[25253] = 25'b01100010_10100011_00000101_1;
      patterns[25254] = 25'b01100010_10100100_00000110_1;
      patterns[25255] = 25'b01100010_10100101_00000111_1;
      patterns[25256] = 25'b01100010_10100110_00001000_1;
      patterns[25257] = 25'b01100010_10100111_00001001_1;
      patterns[25258] = 25'b01100010_10101000_00001010_1;
      patterns[25259] = 25'b01100010_10101001_00001011_1;
      patterns[25260] = 25'b01100010_10101010_00001100_1;
      patterns[25261] = 25'b01100010_10101011_00001101_1;
      patterns[25262] = 25'b01100010_10101100_00001110_1;
      patterns[25263] = 25'b01100010_10101101_00001111_1;
      patterns[25264] = 25'b01100010_10101110_00010000_1;
      patterns[25265] = 25'b01100010_10101111_00010001_1;
      patterns[25266] = 25'b01100010_10110000_00010010_1;
      patterns[25267] = 25'b01100010_10110001_00010011_1;
      patterns[25268] = 25'b01100010_10110010_00010100_1;
      patterns[25269] = 25'b01100010_10110011_00010101_1;
      patterns[25270] = 25'b01100010_10110100_00010110_1;
      patterns[25271] = 25'b01100010_10110101_00010111_1;
      patterns[25272] = 25'b01100010_10110110_00011000_1;
      patterns[25273] = 25'b01100010_10110111_00011001_1;
      patterns[25274] = 25'b01100010_10111000_00011010_1;
      patterns[25275] = 25'b01100010_10111001_00011011_1;
      patterns[25276] = 25'b01100010_10111010_00011100_1;
      patterns[25277] = 25'b01100010_10111011_00011101_1;
      patterns[25278] = 25'b01100010_10111100_00011110_1;
      patterns[25279] = 25'b01100010_10111101_00011111_1;
      patterns[25280] = 25'b01100010_10111110_00100000_1;
      patterns[25281] = 25'b01100010_10111111_00100001_1;
      patterns[25282] = 25'b01100010_11000000_00100010_1;
      patterns[25283] = 25'b01100010_11000001_00100011_1;
      patterns[25284] = 25'b01100010_11000010_00100100_1;
      patterns[25285] = 25'b01100010_11000011_00100101_1;
      patterns[25286] = 25'b01100010_11000100_00100110_1;
      patterns[25287] = 25'b01100010_11000101_00100111_1;
      patterns[25288] = 25'b01100010_11000110_00101000_1;
      patterns[25289] = 25'b01100010_11000111_00101001_1;
      patterns[25290] = 25'b01100010_11001000_00101010_1;
      patterns[25291] = 25'b01100010_11001001_00101011_1;
      patterns[25292] = 25'b01100010_11001010_00101100_1;
      patterns[25293] = 25'b01100010_11001011_00101101_1;
      patterns[25294] = 25'b01100010_11001100_00101110_1;
      patterns[25295] = 25'b01100010_11001101_00101111_1;
      patterns[25296] = 25'b01100010_11001110_00110000_1;
      patterns[25297] = 25'b01100010_11001111_00110001_1;
      patterns[25298] = 25'b01100010_11010000_00110010_1;
      patterns[25299] = 25'b01100010_11010001_00110011_1;
      patterns[25300] = 25'b01100010_11010010_00110100_1;
      patterns[25301] = 25'b01100010_11010011_00110101_1;
      patterns[25302] = 25'b01100010_11010100_00110110_1;
      patterns[25303] = 25'b01100010_11010101_00110111_1;
      patterns[25304] = 25'b01100010_11010110_00111000_1;
      patterns[25305] = 25'b01100010_11010111_00111001_1;
      patterns[25306] = 25'b01100010_11011000_00111010_1;
      patterns[25307] = 25'b01100010_11011001_00111011_1;
      patterns[25308] = 25'b01100010_11011010_00111100_1;
      patterns[25309] = 25'b01100010_11011011_00111101_1;
      patterns[25310] = 25'b01100010_11011100_00111110_1;
      patterns[25311] = 25'b01100010_11011101_00111111_1;
      patterns[25312] = 25'b01100010_11011110_01000000_1;
      patterns[25313] = 25'b01100010_11011111_01000001_1;
      patterns[25314] = 25'b01100010_11100000_01000010_1;
      patterns[25315] = 25'b01100010_11100001_01000011_1;
      patterns[25316] = 25'b01100010_11100010_01000100_1;
      patterns[25317] = 25'b01100010_11100011_01000101_1;
      patterns[25318] = 25'b01100010_11100100_01000110_1;
      patterns[25319] = 25'b01100010_11100101_01000111_1;
      patterns[25320] = 25'b01100010_11100110_01001000_1;
      patterns[25321] = 25'b01100010_11100111_01001001_1;
      patterns[25322] = 25'b01100010_11101000_01001010_1;
      patterns[25323] = 25'b01100010_11101001_01001011_1;
      patterns[25324] = 25'b01100010_11101010_01001100_1;
      patterns[25325] = 25'b01100010_11101011_01001101_1;
      patterns[25326] = 25'b01100010_11101100_01001110_1;
      patterns[25327] = 25'b01100010_11101101_01001111_1;
      patterns[25328] = 25'b01100010_11101110_01010000_1;
      patterns[25329] = 25'b01100010_11101111_01010001_1;
      patterns[25330] = 25'b01100010_11110000_01010010_1;
      patterns[25331] = 25'b01100010_11110001_01010011_1;
      patterns[25332] = 25'b01100010_11110010_01010100_1;
      patterns[25333] = 25'b01100010_11110011_01010101_1;
      patterns[25334] = 25'b01100010_11110100_01010110_1;
      patterns[25335] = 25'b01100010_11110101_01010111_1;
      patterns[25336] = 25'b01100010_11110110_01011000_1;
      patterns[25337] = 25'b01100010_11110111_01011001_1;
      patterns[25338] = 25'b01100010_11111000_01011010_1;
      patterns[25339] = 25'b01100010_11111001_01011011_1;
      patterns[25340] = 25'b01100010_11111010_01011100_1;
      patterns[25341] = 25'b01100010_11111011_01011101_1;
      patterns[25342] = 25'b01100010_11111100_01011110_1;
      patterns[25343] = 25'b01100010_11111101_01011111_1;
      patterns[25344] = 25'b01100010_11111110_01100000_1;
      patterns[25345] = 25'b01100010_11111111_01100001_1;
      patterns[25346] = 25'b01100011_00000000_01100011_0;
      patterns[25347] = 25'b01100011_00000001_01100100_0;
      patterns[25348] = 25'b01100011_00000010_01100101_0;
      patterns[25349] = 25'b01100011_00000011_01100110_0;
      patterns[25350] = 25'b01100011_00000100_01100111_0;
      patterns[25351] = 25'b01100011_00000101_01101000_0;
      patterns[25352] = 25'b01100011_00000110_01101001_0;
      patterns[25353] = 25'b01100011_00000111_01101010_0;
      patterns[25354] = 25'b01100011_00001000_01101011_0;
      patterns[25355] = 25'b01100011_00001001_01101100_0;
      patterns[25356] = 25'b01100011_00001010_01101101_0;
      patterns[25357] = 25'b01100011_00001011_01101110_0;
      patterns[25358] = 25'b01100011_00001100_01101111_0;
      patterns[25359] = 25'b01100011_00001101_01110000_0;
      patterns[25360] = 25'b01100011_00001110_01110001_0;
      patterns[25361] = 25'b01100011_00001111_01110010_0;
      patterns[25362] = 25'b01100011_00010000_01110011_0;
      patterns[25363] = 25'b01100011_00010001_01110100_0;
      patterns[25364] = 25'b01100011_00010010_01110101_0;
      patterns[25365] = 25'b01100011_00010011_01110110_0;
      patterns[25366] = 25'b01100011_00010100_01110111_0;
      patterns[25367] = 25'b01100011_00010101_01111000_0;
      patterns[25368] = 25'b01100011_00010110_01111001_0;
      patterns[25369] = 25'b01100011_00010111_01111010_0;
      patterns[25370] = 25'b01100011_00011000_01111011_0;
      patterns[25371] = 25'b01100011_00011001_01111100_0;
      patterns[25372] = 25'b01100011_00011010_01111101_0;
      patterns[25373] = 25'b01100011_00011011_01111110_0;
      patterns[25374] = 25'b01100011_00011100_01111111_0;
      patterns[25375] = 25'b01100011_00011101_10000000_0;
      patterns[25376] = 25'b01100011_00011110_10000001_0;
      patterns[25377] = 25'b01100011_00011111_10000010_0;
      patterns[25378] = 25'b01100011_00100000_10000011_0;
      patterns[25379] = 25'b01100011_00100001_10000100_0;
      patterns[25380] = 25'b01100011_00100010_10000101_0;
      patterns[25381] = 25'b01100011_00100011_10000110_0;
      patterns[25382] = 25'b01100011_00100100_10000111_0;
      patterns[25383] = 25'b01100011_00100101_10001000_0;
      patterns[25384] = 25'b01100011_00100110_10001001_0;
      patterns[25385] = 25'b01100011_00100111_10001010_0;
      patterns[25386] = 25'b01100011_00101000_10001011_0;
      patterns[25387] = 25'b01100011_00101001_10001100_0;
      patterns[25388] = 25'b01100011_00101010_10001101_0;
      patterns[25389] = 25'b01100011_00101011_10001110_0;
      patterns[25390] = 25'b01100011_00101100_10001111_0;
      patterns[25391] = 25'b01100011_00101101_10010000_0;
      patterns[25392] = 25'b01100011_00101110_10010001_0;
      patterns[25393] = 25'b01100011_00101111_10010010_0;
      patterns[25394] = 25'b01100011_00110000_10010011_0;
      patterns[25395] = 25'b01100011_00110001_10010100_0;
      patterns[25396] = 25'b01100011_00110010_10010101_0;
      patterns[25397] = 25'b01100011_00110011_10010110_0;
      patterns[25398] = 25'b01100011_00110100_10010111_0;
      patterns[25399] = 25'b01100011_00110101_10011000_0;
      patterns[25400] = 25'b01100011_00110110_10011001_0;
      patterns[25401] = 25'b01100011_00110111_10011010_0;
      patterns[25402] = 25'b01100011_00111000_10011011_0;
      patterns[25403] = 25'b01100011_00111001_10011100_0;
      patterns[25404] = 25'b01100011_00111010_10011101_0;
      patterns[25405] = 25'b01100011_00111011_10011110_0;
      patterns[25406] = 25'b01100011_00111100_10011111_0;
      patterns[25407] = 25'b01100011_00111101_10100000_0;
      patterns[25408] = 25'b01100011_00111110_10100001_0;
      patterns[25409] = 25'b01100011_00111111_10100010_0;
      patterns[25410] = 25'b01100011_01000000_10100011_0;
      patterns[25411] = 25'b01100011_01000001_10100100_0;
      patterns[25412] = 25'b01100011_01000010_10100101_0;
      patterns[25413] = 25'b01100011_01000011_10100110_0;
      patterns[25414] = 25'b01100011_01000100_10100111_0;
      patterns[25415] = 25'b01100011_01000101_10101000_0;
      patterns[25416] = 25'b01100011_01000110_10101001_0;
      patterns[25417] = 25'b01100011_01000111_10101010_0;
      patterns[25418] = 25'b01100011_01001000_10101011_0;
      patterns[25419] = 25'b01100011_01001001_10101100_0;
      patterns[25420] = 25'b01100011_01001010_10101101_0;
      patterns[25421] = 25'b01100011_01001011_10101110_0;
      patterns[25422] = 25'b01100011_01001100_10101111_0;
      patterns[25423] = 25'b01100011_01001101_10110000_0;
      patterns[25424] = 25'b01100011_01001110_10110001_0;
      patterns[25425] = 25'b01100011_01001111_10110010_0;
      patterns[25426] = 25'b01100011_01010000_10110011_0;
      patterns[25427] = 25'b01100011_01010001_10110100_0;
      patterns[25428] = 25'b01100011_01010010_10110101_0;
      patterns[25429] = 25'b01100011_01010011_10110110_0;
      patterns[25430] = 25'b01100011_01010100_10110111_0;
      patterns[25431] = 25'b01100011_01010101_10111000_0;
      patterns[25432] = 25'b01100011_01010110_10111001_0;
      patterns[25433] = 25'b01100011_01010111_10111010_0;
      patterns[25434] = 25'b01100011_01011000_10111011_0;
      patterns[25435] = 25'b01100011_01011001_10111100_0;
      patterns[25436] = 25'b01100011_01011010_10111101_0;
      patterns[25437] = 25'b01100011_01011011_10111110_0;
      patterns[25438] = 25'b01100011_01011100_10111111_0;
      patterns[25439] = 25'b01100011_01011101_11000000_0;
      patterns[25440] = 25'b01100011_01011110_11000001_0;
      patterns[25441] = 25'b01100011_01011111_11000010_0;
      patterns[25442] = 25'b01100011_01100000_11000011_0;
      patterns[25443] = 25'b01100011_01100001_11000100_0;
      patterns[25444] = 25'b01100011_01100010_11000101_0;
      patterns[25445] = 25'b01100011_01100011_11000110_0;
      patterns[25446] = 25'b01100011_01100100_11000111_0;
      patterns[25447] = 25'b01100011_01100101_11001000_0;
      patterns[25448] = 25'b01100011_01100110_11001001_0;
      patterns[25449] = 25'b01100011_01100111_11001010_0;
      patterns[25450] = 25'b01100011_01101000_11001011_0;
      patterns[25451] = 25'b01100011_01101001_11001100_0;
      patterns[25452] = 25'b01100011_01101010_11001101_0;
      patterns[25453] = 25'b01100011_01101011_11001110_0;
      patterns[25454] = 25'b01100011_01101100_11001111_0;
      patterns[25455] = 25'b01100011_01101101_11010000_0;
      patterns[25456] = 25'b01100011_01101110_11010001_0;
      patterns[25457] = 25'b01100011_01101111_11010010_0;
      patterns[25458] = 25'b01100011_01110000_11010011_0;
      patterns[25459] = 25'b01100011_01110001_11010100_0;
      patterns[25460] = 25'b01100011_01110010_11010101_0;
      patterns[25461] = 25'b01100011_01110011_11010110_0;
      patterns[25462] = 25'b01100011_01110100_11010111_0;
      patterns[25463] = 25'b01100011_01110101_11011000_0;
      patterns[25464] = 25'b01100011_01110110_11011001_0;
      patterns[25465] = 25'b01100011_01110111_11011010_0;
      patterns[25466] = 25'b01100011_01111000_11011011_0;
      patterns[25467] = 25'b01100011_01111001_11011100_0;
      patterns[25468] = 25'b01100011_01111010_11011101_0;
      patterns[25469] = 25'b01100011_01111011_11011110_0;
      patterns[25470] = 25'b01100011_01111100_11011111_0;
      patterns[25471] = 25'b01100011_01111101_11100000_0;
      patterns[25472] = 25'b01100011_01111110_11100001_0;
      patterns[25473] = 25'b01100011_01111111_11100010_0;
      patterns[25474] = 25'b01100011_10000000_11100011_0;
      patterns[25475] = 25'b01100011_10000001_11100100_0;
      patterns[25476] = 25'b01100011_10000010_11100101_0;
      patterns[25477] = 25'b01100011_10000011_11100110_0;
      patterns[25478] = 25'b01100011_10000100_11100111_0;
      patterns[25479] = 25'b01100011_10000101_11101000_0;
      patterns[25480] = 25'b01100011_10000110_11101001_0;
      patterns[25481] = 25'b01100011_10000111_11101010_0;
      patterns[25482] = 25'b01100011_10001000_11101011_0;
      patterns[25483] = 25'b01100011_10001001_11101100_0;
      patterns[25484] = 25'b01100011_10001010_11101101_0;
      patterns[25485] = 25'b01100011_10001011_11101110_0;
      patterns[25486] = 25'b01100011_10001100_11101111_0;
      patterns[25487] = 25'b01100011_10001101_11110000_0;
      patterns[25488] = 25'b01100011_10001110_11110001_0;
      patterns[25489] = 25'b01100011_10001111_11110010_0;
      patterns[25490] = 25'b01100011_10010000_11110011_0;
      patterns[25491] = 25'b01100011_10010001_11110100_0;
      patterns[25492] = 25'b01100011_10010010_11110101_0;
      patterns[25493] = 25'b01100011_10010011_11110110_0;
      patterns[25494] = 25'b01100011_10010100_11110111_0;
      patterns[25495] = 25'b01100011_10010101_11111000_0;
      patterns[25496] = 25'b01100011_10010110_11111001_0;
      patterns[25497] = 25'b01100011_10010111_11111010_0;
      patterns[25498] = 25'b01100011_10011000_11111011_0;
      patterns[25499] = 25'b01100011_10011001_11111100_0;
      patterns[25500] = 25'b01100011_10011010_11111101_0;
      patterns[25501] = 25'b01100011_10011011_11111110_0;
      patterns[25502] = 25'b01100011_10011100_11111111_0;
      patterns[25503] = 25'b01100011_10011101_00000000_1;
      patterns[25504] = 25'b01100011_10011110_00000001_1;
      patterns[25505] = 25'b01100011_10011111_00000010_1;
      patterns[25506] = 25'b01100011_10100000_00000011_1;
      patterns[25507] = 25'b01100011_10100001_00000100_1;
      patterns[25508] = 25'b01100011_10100010_00000101_1;
      patterns[25509] = 25'b01100011_10100011_00000110_1;
      patterns[25510] = 25'b01100011_10100100_00000111_1;
      patterns[25511] = 25'b01100011_10100101_00001000_1;
      patterns[25512] = 25'b01100011_10100110_00001001_1;
      patterns[25513] = 25'b01100011_10100111_00001010_1;
      patterns[25514] = 25'b01100011_10101000_00001011_1;
      patterns[25515] = 25'b01100011_10101001_00001100_1;
      patterns[25516] = 25'b01100011_10101010_00001101_1;
      patterns[25517] = 25'b01100011_10101011_00001110_1;
      patterns[25518] = 25'b01100011_10101100_00001111_1;
      patterns[25519] = 25'b01100011_10101101_00010000_1;
      patterns[25520] = 25'b01100011_10101110_00010001_1;
      patterns[25521] = 25'b01100011_10101111_00010010_1;
      patterns[25522] = 25'b01100011_10110000_00010011_1;
      patterns[25523] = 25'b01100011_10110001_00010100_1;
      patterns[25524] = 25'b01100011_10110010_00010101_1;
      patterns[25525] = 25'b01100011_10110011_00010110_1;
      patterns[25526] = 25'b01100011_10110100_00010111_1;
      patterns[25527] = 25'b01100011_10110101_00011000_1;
      patterns[25528] = 25'b01100011_10110110_00011001_1;
      patterns[25529] = 25'b01100011_10110111_00011010_1;
      patterns[25530] = 25'b01100011_10111000_00011011_1;
      patterns[25531] = 25'b01100011_10111001_00011100_1;
      patterns[25532] = 25'b01100011_10111010_00011101_1;
      patterns[25533] = 25'b01100011_10111011_00011110_1;
      patterns[25534] = 25'b01100011_10111100_00011111_1;
      patterns[25535] = 25'b01100011_10111101_00100000_1;
      patterns[25536] = 25'b01100011_10111110_00100001_1;
      patterns[25537] = 25'b01100011_10111111_00100010_1;
      patterns[25538] = 25'b01100011_11000000_00100011_1;
      patterns[25539] = 25'b01100011_11000001_00100100_1;
      patterns[25540] = 25'b01100011_11000010_00100101_1;
      patterns[25541] = 25'b01100011_11000011_00100110_1;
      patterns[25542] = 25'b01100011_11000100_00100111_1;
      patterns[25543] = 25'b01100011_11000101_00101000_1;
      patterns[25544] = 25'b01100011_11000110_00101001_1;
      patterns[25545] = 25'b01100011_11000111_00101010_1;
      patterns[25546] = 25'b01100011_11001000_00101011_1;
      patterns[25547] = 25'b01100011_11001001_00101100_1;
      patterns[25548] = 25'b01100011_11001010_00101101_1;
      patterns[25549] = 25'b01100011_11001011_00101110_1;
      patterns[25550] = 25'b01100011_11001100_00101111_1;
      patterns[25551] = 25'b01100011_11001101_00110000_1;
      patterns[25552] = 25'b01100011_11001110_00110001_1;
      patterns[25553] = 25'b01100011_11001111_00110010_1;
      patterns[25554] = 25'b01100011_11010000_00110011_1;
      patterns[25555] = 25'b01100011_11010001_00110100_1;
      patterns[25556] = 25'b01100011_11010010_00110101_1;
      patterns[25557] = 25'b01100011_11010011_00110110_1;
      patterns[25558] = 25'b01100011_11010100_00110111_1;
      patterns[25559] = 25'b01100011_11010101_00111000_1;
      patterns[25560] = 25'b01100011_11010110_00111001_1;
      patterns[25561] = 25'b01100011_11010111_00111010_1;
      patterns[25562] = 25'b01100011_11011000_00111011_1;
      patterns[25563] = 25'b01100011_11011001_00111100_1;
      patterns[25564] = 25'b01100011_11011010_00111101_1;
      patterns[25565] = 25'b01100011_11011011_00111110_1;
      patterns[25566] = 25'b01100011_11011100_00111111_1;
      patterns[25567] = 25'b01100011_11011101_01000000_1;
      patterns[25568] = 25'b01100011_11011110_01000001_1;
      patterns[25569] = 25'b01100011_11011111_01000010_1;
      patterns[25570] = 25'b01100011_11100000_01000011_1;
      patterns[25571] = 25'b01100011_11100001_01000100_1;
      patterns[25572] = 25'b01100011_11100010_01000101_1;
      patterns[25573] = 25'b01100011_11100011_01000110_1;
      patterns[25574] = 25'b01100011_11100100_01000111_1;
      patterns[25575] = 25'b01100011_11100101_01001000_1;
      patterns[25576] = 25'b01100011_11100110_01001001_1;
      patterns[25577] = 25'b01100011_11100111_01001010_1;
      patterns[25578] = 25'b01100011_11101000_01001011_1;
      patterns[25579] = 25'b01100011_11101001_01001100_1;
      patterns[25580] = 25'b01100011_11101010_01001101_1;
      patterns[25581] = 25'b01100011_11101011_01001110_1;
      patterns[25582] = 25'b01100011_11101100_01001111_1;
      patterns[25583] = 25'b01100011_11101101_01010000_1;
      patterns[25584] = 25'b01100011_11101110_01010001_1;
      patterns[25585] = 25'b01100011_11101111_01010010_1;
      patterns[25586] = 25'b01100011_11110000_01010011_1;
      patterns[25587] = 25'b01100011_11110001_01010100_1;
      patterns[25588] = 25'b01100011_11110010_01010101_1;
      patterns[25589] = 25'b01100011_11110011_01010110_1;
      patterns[25590] = 25'b01100011_11110100_01010111_1;
      patterns[25591] = 25'b01100011_11110101_01011000_1;
      patterns[25592] = 25'b01100011_11110110_01011001_1;
      patterns[25593] = 25'b01100011_11110111_01011010_1;
      patterns[25594] = 25'b01100011_11111000_01011011_1;
      patterns[25595] = 25'b01100011_11111001_01011100_1;
      patterns[25596] = 25'b01100011_11111010_01011101_1;
      patterns[25597] = 25'b01100011_11111011_01011110_1;
      patterns[25598] = 25'b01100011_11111100_01011111_1;
      patterns[25599] = 25'b01100011_11111101_01100000_1;
      patterns[25600] = 25'b01100011_11111110_01100001_1;
      patterns[25601] = 25'b01100011_11111111_01100010_1;
      patterns[25602] = 25'b01100100_00000000_01100100_0;
      patterns[25603] = 25'b01100100_00000001_01100101_0;
      patterns[25604] = 25'b01100100_00000010_01100110_0;
      patterns[25605] = 25'b01100100_00000011_01100111_0;
      patterns[25606] = 25'b01100100_00000100_01101000_0;
      patterns[25607] = 25'b01100100_00000101_01101001_0;
      patterns[25608] = 25'b01100100_00000110_01101010_0;
      patterns[25609] = 25'b01100100_00000111_01101011_0;
      patterns[25610] = 25'b01100100_00001000_01101100_0;
      patterns[25611] = 25'b01100100_00001001_01101101_0;
      patterns[25612] = 25'b01100100_00001010_01101110_0;
      patterns[25613] = 25'b01100100_00001011_01101111_0;
      patterns[25614] = 25'b01100100_00001100_01110000_0;
      patterns[25615] = 25'b01100100_00001101_01110001_0;
      patterns[25616] = 25'b01100100_00001110_01110010_0;
      patterns[25617] = 25'b01100100_00001111_01110011_0;
      patterns[25618] = 25'b01100100_00010000_01110100_0;
      patterns[25619] = 25'b01100100_00010001_01110101_0;
      patterns[25620] = 25'b01100100_00010010_01110110_0;
      patterns[25621] = 25'b01100100_00010011_01110111_0;
      patterns[25622] = 25'b01100100_00010100_01111000_0;
      patterns[25623] = 25'b01100100_00010101_01111001_0;
      patterns[25624] = 25'b01100100_00010110_01111010_0;
      patterns[25625] = 25'b01100100_00010111_01111011_0;
      patterns[25626] = 25'b01100100_00011000_01111100_0;
      patterns[25627] = 25'b01100100_00011001_01111101_0;
      patterns[25628] = 25'b01100100_00011010_01111110_0;
      patterns[25629] = 25'b01100100_00011011_01111111_0;
      patterns[25630] = 25'b01100100_00011100_10000000_0;
      patterns[25631] = 25'b01100100_00011101_10000001_0;
      patterns[25632] = 25'b01100100_00011110_10000010_0;
      patterns[25633] = 25'b01100100_00011111_10000011_0;
      patterns[25634] = 25'b01100100_00100000_10000100_0;
      patterns[25635] = 25'b01100100_00100001_10000101_0;
      patterns[25636] = 25'b01100100_00100010_10000110_0;
      patterns[25637] = 25'b01100100_00100011_10000111_0;
      patterns[25638] = 25'b01100100_00100100_10001000_0;
      patterns[25639] = 25'b01100100_00100101_10001001_0;
      patterns[25640] = 25'b01100100_00100110_10001010_0;
      patterns[25641] = 25'b01100100_00100111_10001011_0;
      patterns[25642] = 25'b01100100_00101000_10001100_0;
      patterns[25643] = 25'b01100100_00101001_10001101_0;
      patterns[25644] = 25'b01100100_00101010_10001110_0;
      patterns[25645] = 25'b01100100_00101011_10001111_0;
      patterns[25646] = 25'b01100100_00101100_10010000_0;
      patterns[25647] = 25'b01100100_00101101_10010001_0;
      patterns[25648] = 25'b01100100_00101110_10010010_0;
      patterns[25649] = 25'b01100100_00101111_10010011_0;
      patterns[25650] = 25'b01100100_00110000_10010100_0;
      patterns[25651] = 25'b01100100_00110001_10010101_0;
      patterns[25652] = 25'b01100100_00110010_10010110_0;
      patterns[25653] = 25'b01100100_00110011_10010111_0;
      patterns[25654] = 25'b01100100_00110100_10011000_0;
      patterns[25655] = 25'b01100100_00110101_10011001_0;
      patterns[25656] = 25'b01100100_00110110_10011010_0;
      patterns[25657] = 25'b01100100_00110111_10011011_0;
      patterns[25658] = 25'b01100100_00111000_10011100_0;
      patterns[25659] = 25'b01100100_00111001_10011101_0;
      patterns[25660] = 25'b01100100_00111010_10011110_0;
      patterns[25661] = 25'b01100100_00111011_10011111_0;
      patterns[25662] = 25'b01100100_00111100_10100000_0;
      patterns[25663] = 25'b01100100_00111101_10100001_0;
      patterns[25664] = 25'b01100100_00111110_10100010_0;
      patterns[25665] = 25'b01100100_00111111_10100011_0;
      patterns[25666] = 25'b01100100_01000000_10100100_0;
      patterns[25667] = 25'b01100100_01000001_10100101_0;
      patterns[25668] = 25'b01100100_01000010_10100110_0;
      patterns[25669] = 25'b01100100_01000011_10100111_0;
      patterns[25670] = 25'b01100100_01000100_10101000_0;
      patterns[25671] = 25'b01100100_01000101_10101001_0;
      patterns[25672] = 25'b01100100_01000110_10101010_0;
      patterns[25673] = 25'b01100100_01000111_10101011_0;
      patterns[25674] = 25'b01100100_01001000_10101100_0;
      patterns[25675] = 25'b01100100_01001001_10101101_0;
      patterns[25676] = 25'b01100100_01001010_10101110_0;
      patterns[25677] = 25'b01100100_01001011_10101111_0;
      patterns[25678] = 25'b01100100_01001100_10110000_0;
      patterns[25679] = 25'b01100100_01001101_10110001_0;
      patterns[25680] = 25'b01100100_01001110_10110010_0;
      patterns[25681] = 25'b01100100_01001111_10110011_0;
      patterns[25682] = 25'b01100100_01010000_10110100_0;
      patterns[25683] = 25'b01100100_01010001_10110101_0;
      patterns[25684] = 25'b01100100_01010010_10110110_0;
      patterns[25685] = 25'b01100100_01010011_10110111_0;
      patterns[25686] = 25'b01100100_01010100_10111000_0;
      patterns[25687] = 25'b01100100_01010101_10111001_0;
      patterns[25688] = 25'b01100100_01010110_10111010_0;
      patterns[25689] = 25'b01100100_01010111_10111011_0;
      patterns[25690] = 25'b01100100_01011000_10111100_0;
      patterns[25691] = 25'b01100100_01011001_10111101_0;
      patterns[25692] = 25'b01100100_01011010_10111110_0;
      patterns[25693] = 25'b01100100_01011011_10111111_0;
      patterns[25694] = 25'b01100100_01011100_11000000_0;
      patterns[25695] = 25'b01100100_01011101_11000001_0;
      patterns[25696] = 25'b01100100_01011110_11000010_0;
      patterns[25697] = 25'b01100100_01011111_11000011_0;
      patterns[25698] = 25'b01100100_01100000_11000100_0;
      patterns[25699] = 25'b01100100_01100001_11000101_0;
      patterns[25700] = 25'b01100100_01100010_11000110_0;
      patterns[25701] = 25'b01100100_01100011_11000111_0;
      patterns[25702] = 25'b01100100_01100100_11001000_0;
      patterns[25703] = 25'b01100100_01100101_11001001_0;
      patterns[25704] = 25'b01100100_01100110_11001010_0;
      patterns[25705] = 25'b01100100_01100111_11001011_0;
      patterns[25706] = 25'b01100100_01101000_11001100_0;
      patterns[25707] = 25'b01100100_01101001_11001101_0;
      patterns[25708] = 25'b01100100_01101010_11001110_0;
      patterns[25709] = 25'b01100100_01101011_11001111_0;
      patterns[25710] = 25'b01100100_01101100_11010000_0;
      patterns[25711] = 25'b01100100_01101101_11010001_0;
      patterns[25712] = 25'b01100100_01101110_11010010_0;
      patterns[25713] = 25'b01100100_01101111_11010011_0;
      patterns[25714] = 25'b01100100_01110000_11010100_0;
      patterns[25715] = 25'b01100100_01110001_11010101_0;
      patterns[25716] = 25'b01100100_01110010_11010110_0;
      patterns[25717] = 25'b01100100_01110011_11010111_0;
      patterns[25718] = 25'b01100100_01110100_11011000_0;
      patterns[25719] = 25'b01100100_01110101_11011001_0;
      patterns[25720] = 25'b01100100_01110110_11011010_0;
      patterns[25721] = 25'b01100100_01110111_11011011_0;
      patterns[25722] = 25'b01100100_01111000_11011100_0;
      patterns[25723] = 25'b01100100_01111001_11011101_0;
      patterns[25724] = 25'b01100100_01111010_11011110_0;
      patterns[25725] = 25'b01100100_01111011_11011111_0;
      patterns[25726] = 25'b01100100_01111100_11100000_0;
      patterns[25727] = 25'b01100100_01111101_11100001_0;
      patterns[25728] = 25'b01100100_01111110_11100010_0;
      patterns[25729] = 25'b01100100_01111111_11100011_0;
      patterns[25730] = 25'b01100100_10000000_11100100_0;
      patterns[25731] = 25'b01100100_10000001_11100101_0;
      patterns[25732] = 25'b01100100_10000010_11100110_0;
      patterns[25733] = 25'b01100100_10000011_11100111_0;
      patterns[25734] = 25'b01100100_10000100_11101000_0;
      patterns[25735] = 25'b01100100_10000101_11101001_0;
      patterns[25736] = 25'b01100100_10000110_11101010_0;
      patterns[25737] = 25'b01100100_10000111_11101011_0;
      patterns[25738] = 25'b01100100_10001000_11101100_0;
      patterns[25739] = 25'b01100100_10001001_11101101_0;
      patterns[25740] = 25'b01100100_10001010_11101110_0;
      patterns[25741] = 25'b01100100_10001011_11101111_0;
      patterns[25742] = 25'b01100100_10001100_11110000_0;
      patterns[25743] = 25'b01100100_10001101_11110001_0;
      patterns[25744] = 25'b01100100_10001110_11110010_0;
      patterns[25745] = 25'b01100100_10001111_11110011_0;
      patterns[25746] = 25'b01100100_10010000_11110100_0;
      patterns[25747] = 25'b01100100_10010001_11110101_0;
      patterns[25748] = 25'b01100100_10010010_11110110_0;
      patterns[25749] = 25'b01100100_10010011_11110111_0;
      patterns[25750] = 25'b01100100_10010100_11111000_0;
      patterns[25751] = 25'b01100100_10010101_11111001_0;
      patterns[25752] = 25'b01100100_10010110_11111010_0;
      patterns[25753] = 25'b01100100_10010111_11111011_0;
      patterns[25754] = 25'b01100100_10011000_11111100_0;
      patterns[25755] = 25'b01100100_10011001_11111101_0;
      patterns[25756] = 25'b01100100_10011010_11111110_0;
      patterns[25757] = 25'b01100100_10011011_11111111_0;
      patterns[25758] = 25'b01100100_10011100_00000000_1;
      patterns[25759] = 25'b01100100_10011101_00000001_1;
      patterns[25760] = 25'b01100100_10011110_00000010_1;
      patterns[25761] = 25'b01100100_10011111_00000011_1;
      patterns[25762] = 25'b01100100_10100000_00000100_1;
      patterns[25763] = 25'b01100100_10100001_00000101_1;
      patterns[25764] = 25'b01100100_10100010_00000110_1;
      patterns[25765] = 25'b01100100_10100011_00000111_1;
      patterns[25766] = 25'b01100100_10100100_00001000_1;
      patterns[25767] = 25'b01100100_10100101_00001001_1;
      patterns[25768] = 25'b01100100_10100110_00001010_1;
      patterns[25769] = 25'b01100100_10100111_00001011_1;
      patterns[25770] = 25'b01100100_10101000_00001100_1;
      patterns[25771] = 25'b01100100_10101001_00001101_1;
      patterns[25772] = 25'b01100100_10101010_00001110_1;
      patterns[25773] = 25'b01100100_10101011_00001111_1;
      patterns[25774] = 25'b01100100_10101100_00010000_1;
      patterns[25775] = 25'b01100100_10101101_00010001_1;
      patterns[25776] = 25'b01100100_10101110_00010010_1;
      patterns[25777] = 25'b01100100_10101111_00010011_1;
      patterns[25778] = 25'b01100100_10110000_00010100_1;
      patterns[25779] = 25'b01100100_10110001_00010101_1;
      patterns[25780] = 25'b01100100_10110010_00010110_1;
      patterns[25781] = 25'b01100100_10110011_00010111_1;
      patterns[25782] = 25'b01100100_10110100_00011000_1;
      patterns[25783] = 25'b01100100_10110101_00011001_1;
      patterns[25784] = 25'b01100100_10110110_00011010_1;
      patterns[25785] = 25'b01100100_10110111_00011011_1;
      patterns[25786] = 25'b01100100_10111000_00011100_1;
      patterns[25787] = 25'b01100100_10111001_00011101_1;
      patterns[25788] = 25'b01100100_10111010_00011110_1;
      patterns[25789] = 25'b01100100_10111011_00011111_1;
      patterns[25790] = 25'b01100100_10111100_00100000_1;
      patterns[25791] = 25'b01100100_10111101_00100001_1;
      patterns[25792] = 25'b01100100_10111110_00100010_1;
      patterns[25793] = 25'b01100100_10111111_00100011_1;
      patterns[25794] = 25'b01100100_11000000_00100100_1;
      patterns[25795] = 25'b01100100_11000001_00100101_1;
      patterns[25796] = 25'b01100100_11000010_00100110_1;
      patterns[25797] = 25'b01100100_11000011_00100111_1;
      patterns[25798] = 25'b01100100_11000100_00101000_1;
      patterns[25799] = 25'b01100100_11000101_00101001_1;
      patterns[25800] = 25'b01100100_11000110_00101010_1;
      patterns[25801] = 25'b01100100_11000111_00101011_1;
      patterns[25802] = 25'b01100100_11001000_00101100_1;
      patterns[25803] = 25'b01100100_11001001_00101101_1;
      patterns[25804] = 25'b01100100_11001010_00101110_1;
      patterns[25805] = 25'b01100100_11001011_00101111_1;
      patterns[25806] = 25'b01100100_11001100_00110000_1;
      patterns[25807] = 25'b01100100_11001101_00110001_1;
      patterns[25808] = 25'b01100100_11001110_00110010_1;
      patterns[25809] = 25'b01100100_11001111_00110011_1;
      patterns[25810] = 25'b01100100_11010000_00110100_1;
      patterns[25811] = 25'b01100100_11010001_00110101_1;
      patterns[25812] = 25'b01100100_11010010_00110110_1;
      patterns[25813] = 25'b01100100_11010011_00110111_1;
      patterns[25814] = 25'b01100100_11010100_00111000_1;
      patterns[25815] = 25'b01100100_11010101_00111001_1;
      patterns[25816] = 25'b01100100_11010110_00111010_1;
      patterns[25817] = 25'b01100100_11010111_00111011_1;
      patterns[25818] = 25'b01100100_11011000_00111100_1;
      patterns[25819] = 25'b01100100_11011001_00111101_1;
      patterns[25820] = 25'b01100100_11011010_00111110_1;
      patterns[25821] = 25'b01100100_11011011_00111111_1;
      patterns[25822] = 25'b01100100_11011100_01000000_1;
      patterns[25823] = 25'b01100100_11011101_01000001_1;
      patterns[25824] = 25'b01100100_11011110_01000010_1;
      patterns[25825] = 25'b01100100_11011111_01000011_1;
      patterns[25826] = 25'b01100100_11100000_01000100_1;
      patterns[25827] = 25'b01100100_11100001_01000101_1;
      patterns[25828] = 25'b01100100_11100010_01000110_1;
      patterns[25829] = 25'b01100100_11100011_01000111_1;
      patterns[25830] = 25'b01100100_11100100_01001000_1;
      patterns[25831] = 25'b01100100_11100101_01001001_1;
      patterns[25832] = 25'b01100100_11100110_01001010_1;
      patterns[25833] = 25'b01100100_11100111_01001011_1;
      patterns[25834] = 25'b01100100_11101000_01001100_1;
      patterns[25835] = 25'b01100100_11101001_01001101_1;
      patterns[25836] = 25'b01100100_11101010_01001110_1;
      patterns[25837] = 25'b01100100_11101011_01001111_1;
      patterns[25838] = 25'b01100100_11101100_01010000_1;
      patterns[25839] = 25'b01100100_11101101_01010001_1;
      patterns[25840] = 25'b01100100_11101110_01010010_1;
      patterns[25841] = 25'b01100100_11101111_01010011_1;
      patterns[25842] = 25'b01100100_11110000_01010100_1;
      patterns[25843] = 25'b01100100_11110001_01010101_1;
      patterns[25844] = 25'b01100100_11110010_01010110_1;
      patterns[25845] = 25'b01100100_11110011_01010111_1;
      patterns[25846] = 25'b01100100_11110100_01011000_1;
      patterns[25847] = 25'b01100100_11110101_01011001_1;
      patterns[25848] = 25'b01100100_11110110_01011010_1;
      patterns[25849] = 25'b01100100_11110111_01011011_1;
      patterns[25850] = 25'b01100100_11111000_01011100_1;
      patterns[25851] = 25'b01100100_11111001_01011101_1;
      patterns[25852] = 25'b01100100_11111010_01011110_1;
      patterns[25853] = 25'b01100100_11111011_01011111_1;
      patterns[25854] = 25'b01100100_11111100_01100000_1;
      patterns[25855] = 25'b01100100_11111101_01100001_1;
      patterns[25856] = 25'b01100100_11111110_01100010_1;
      patterns[25857] = 25'b01100100_11111111_01100011_1;
      patterns[25858] = 25'b01100101_00000000_01100101_0;
      patterns[25859] = 25'b01100101_00000001_01100110_0;
      patterns[25860] = 25'b01100101_00000010_01100111_0;
      patterns[25861] = 25'b01100101_00000011_01101000_0;
      patterns[25862] = 25'b01100101_00000100_01101001_0;
      patterns[25863] = 25'b01100101_00000101_01101010_0;
      patterns[25864] = 25'b01100101_00000110_01101011_0;
      patterns[25865] = 25'b01100101_00000111_01101100_0;
      patterns[25866] = 25'b01100101_00001000_01101101_0;
      patterns[25867] = 25'b01100101_00001001_01101110_0;
      patterns[25868] = 25'b01100101_00001010_01101111_0;
      patterns[25869] = 25'b01100101_00001011_01110000_0;
      patterns[25870] = 25'b01100101_00001100_01110001_0;
      patterns[25871] = 25'b01100101_00001101_01110010_0;
      patterns[25872] = 25'b01100101_00001110_01110011_0;
      patterns[25873] = 25'b01100101_00001111_01110100_0;
      patterns[25874] = 25'b01100101_00010000_01110101_0;
      patterns[25875] = 25'b01100101_00010001_01110110_0;
      patterns[25876] = 25'b01100101_00010010_01110111_0;
      patterns[25877] = 25'b01100101_00010011_01111000_0;
      patterns[25878] = 25'b01100101_00010100_01111001_0;
      patterns[25879] = 25'b01100101_00010101_01111010_0;
      patterns[25880] = 25'b01100101_00010110_01111011_0;
      patterns[25881] = 25'b01100101_00010111_01111100_0;
      patterns[25882] = 25'b01100101_00011000_01111101_0;
      patterns[25883] = 25'b01100101_00011001_01111110_0;
      patterns[25884] = 25'b01100101_00011010_01111111_0;
      patterns[25885] = 25'b01100101_00011011_10000000_0;
      patterns[25886] = 25'b01100101_00011100_10000001_0;
      patterns[25887] = 25'b01100101_00011101_10000010_0;
      patterns[25888] = 25'b01100101_00011110_10000011_0;
      patterns[25889] = 25'b01100101_00011111_10000100_0;
      patterns[25890] = 25'b01100101_00100000_10000101_0;
      patterns[25891] = 25'b01100101_00100001_10000110_0;
      patterns[25892] = 25'b01100101_00100010_10000111_0;
      patterns[25893] = 25'b01100101_00100011_10001000_0;
      patterns[25894] = 25'b01100101_00100100_10001001_0;
      patterns[25895] = 25'b01100101_00100101_10001010_0;
      patterns[25896] = 25'b01100101_00100110_10001011_0;
      patterns[25897] = 25'b01100101_00100111_10001100_0;
      patterns[25898] = 25'b01100101_00101000_10001101_0;
      patterns[25899] = 25'b01100101_00101001_10001110_0;
      patterns[25900] = 25'b01100101_00101010_10001111_0;
      patterns[25901] = 25'b01100101_00101011_10010000_0;
      patterns[25902] = 25'b01100101_00101100_10010001_0;
      patterns[25903] = 25'b01100101_00101101_10010010_0;
      patterns[25904] = 25'b01100101_00101110_10010011_0;
      patterns[25905] = 25'b01100101_00101111_10010100_0;
      patterns[25906] = 25'b01100101_00110000_10010101_0;
      patterns[25907] = 25'b01100101_00110001_10010110_0;
      patterns[25908] = 25'b01100101_00110010_10010111_0;
      patterns[25909] = 25'b01100101_00110011_10011000_0;
      patterns[25910] = 25'b01100101_00110100_10011001_0;
      patterns[25911] = 25'b01100101_00110101_10011010_0;
      patterns[25912] = 25'b01100101_00110110_10011011_0;
      patterns[25913] = 25'b01100101_00110111_10011100_0;
      patterns[25914] = 25'b01100101_00111000_10011101_0;
      patterns[25915] = 25'b01100101_00111001_10011110_0;
      patterns[25916] = 25'b01100101_00111010_10011111_0;
      patterns[25917] = 25'b01100101_00111011_10100000_0;
      patterns[25918] = 25'b01100101_00111100_10100001_0;
      patterns[25919] = 25'b01100101_00111101_10100010_0;
      patterns[25920] = 25'b01100101_00111110_10100011_0;
      patterns[25921] = 25'b01100101_00111111_10100100_0;
      patterns[25922] = 25'b01100101_01000000_10100101_0;
      patterns[25923] = 25'b01100101_01000001_10100110_0;
      patterns[25924] = 25'b01100101_01000010_10100111_0;
      patterns[25925] = 25'b01100101_01000011_10101000_0;
      patterns[25926] = 25'b01100101_01000100_10101001_0;
      patterns[25927] = 25'b01100101_01000101_10101010_0;
      patterns[25928] = 25'b01100101_01000110_10101011_0;
      patterns[25929] = 25'b01100101_01000111_10101100_0;
      patterns[25930] = 25'b01100101_01001000_10101101_0;
      patterns[25931] = 25'b01100101_01001001_10101110_0;
      patterns[25932] = 25'b01100101_01001010_10101111_0;
      patterns[25933] = 25'b01100101_01001011_10110000_0;
      patterns[25934] = 25'b01100101_01001100_10110001_0;
      patterns[25935] = 25'b01100101_01001101_10110010_0;
      patterns[25936] = 25'b01100101_01001110_10110011_0;
      patterns[25937] = 25'b01100101_01001111_10110100_0;
      patterns[25938] = 25'b01100101_01010000_10110101_0;
      patterns[25939] = 25'b01100101_01010001_10110110_0;
      patterns[25940] = 25'b01100101_01010010_10110111_0;
      patterns[25941] = 25'b01100101_01010011_10111000_0;
      patterns[25942] = 25'b01100101_01010100_10111001_0;
      patterns[25943] = 25'b01100101_01010101_10111010_0;
      patterns[25944] = 25'b01100101_01010110_10111011_0;
      patterns[25945] = 25'b01100101_01010111_10111100_0;
      patterns[25946] = 25'b01100101_01011000_10111101_0;
      patterns[25947] = 25'b01100101_01011001_10111110_0;
      patterns[25948] = 25'b01100101_01011010_10111111_0;
      patterns[25949] = 25'b01100101_01011011_11000000_0;
      patterns[25950] = 25'b01100101_01011100_11000001_0;
      patterns[25951] = 25'b01100101_01011101_11000010_0;
      patterns[25952] = 25'b01100101_01011110_11000011_0;
      patterns[25953] = 25'b01100101_01011111_11000100_0;
      patterns[25954] = 25'b01100101_01100000_11000101_0;
      patterns[25955] = 25'b01100101_01100001_11000110_0;
      patterns[25956] = 25'b01100101_01100010_11000111_0;
      patterns[25957] = 25'b01100101_01100011_11001000_0;
      patterns[25958] = 25'b01100101_01100100_11001001_0;
      patterns[25959] = 25'b01100101_01100101_11001010_0;
      patterns[25960] = 25'b01100101_01100110_11001011_0;
      patterns[25961] = 25'b01100101_01100111_11001100_0;
      patterns[25962] = 25'b01100101_01101000_11001101_0;
      patterns[25963] = 25'b01100101_01101001_11001110_0;
      patterns[25964] = 25'b01100101_01101010_11001111_0;
      patterns[25965] = 25'b01100101_01101011_11010000_0;
      patterns[25966] = 25'b01100101_01101100_11010001_0;
      patterns[25967] = 25'b01100101_01101101_11010010_0;
      patterns[25968] = 25'b01100101_01101110_11010011_0;
      patterns[25969] = 25'b01100101_01101111_11010100_0;
      patterns[25970] = 25'b01100101_01110000_11010101_0;
      patterns[25971] = 25'b01100101_01110001_11010110_0;
      patterns[25972] = 25'b01100101_01110010_11010111_0;
      patterns[25973] = 25'b01100101_01110011_11011000_0;
      patterns[25974] = 25'b01100101_01110100_11011001_0;
      patterns[25975] = 25'b01100101_01110101_11011010_0;
      patterns[25976] = 25'b01100101_01110110_11011011_0;
      patterns[25977] = 25'b01100101_01110111_11011100_0;
      patterns[25978] = 25'b01100101_01111000_11011101_0;
      patterns[25979] = 25'b01100101_01111001_11011110_0;
      patterns[25980] = 25'b01100101_01111010_11011111_0;
      patterns[25981] = 25'b01100101_01111011_11100000_0;
      patterns[25982] = 25'b01100101_01111100_11100001_0;
      patterns[25983] = 25'b01100101_01111101_11100010_0;
      patterns[25984] = 25'b01100101_01111110_11100011_0;
      patterns[25985] = 25'b01100101_01111111_11100100_0;
      patterns[25986] = 25'b01100101_10000000_11100101_0;
      patterns[25987] = 25'b01100101_10000001_11100110_0;
      patterns[25988] = 25'b01100101_10000010_11100111_0;
      patterns[25989] = 25'b01100101_10000011_11101000_0;
      patterns[25990] = 25'b01100101_10000100_11101001_0;
      patterns[25991] = 25'b01100101_10000101_11101010_0;
      patterns[25992] = 25'b01100101_10000110_11101011_0;
      patterns[25993] = 25'b01100101_10000111_11101100_0;
      patterns[25994] = 25'b01100101_10001000_11101101_0;
      patterns[25995] = 25'b01100101_10001001_11101110_0;
      patterns[25996] = 25'b01100101_10001010_11101111_0;
      patterns[25997] = 25'b01100101_10001011_11110000_0;
      patterns[25998] = 25'b01100101_10001100_11110001_0;
      patterns[25999] = 25'b01100101_10001101_11110010_0;
      patterns[26000] = 25'b01100101_10001110_11110011_0;
      patterns[26001] = 25'b01100101_10001111_11110100_0;
      patterns[26002] = 25'b01100101_10010000_11110101_0;
      patterns[26003] = 25'b01100101_10010001_11110110_0;
      patterns[26004] = 25'b01100101_10010010_11110111_0;
      patterns[26005] = 25'b01100101_10010011_11111000_0;
      patterns[26006] = 25'b01100101_10010100_11111001_0;
      patterns[26007] = 25'b01100101_10010101_11111010_0;
      patterns[26008] = 25'b01100101_10010110_11111011_0;
      patterns[26009] = 25'b01100101_10010111_11111100_0;
      patterns[26010] = 25'b01100101_10011000_11111101_0;
      patterns[26011] = 25'b01100101_10011001_11111110_0;
      patterns[26012] = 25'b01100101_10011010_11111111_0;
      patterns[26013] = 25'b01100101_10011011_00000000_1;
      patterns[26014] = 25'b01100101_10011100_00000001_1;
      patterns[26015] = 25'b01100101_10011101_00000010_1;
      patterns[26016] = 25'b01100101_10011110_00000011_1;
      patterns[26017] = 25'b01100101_10011111_00000100_1;
      patterns[26018] = 25'b01100101_10100000_00000101_1;
      patterns[26019] = 25'b01100101_10100001_00000110_1;
      patterns[26020] = 25'b01100101_10100010_00000111_1;
      patterns[26021] = 25'b01100101_10100011_00001000_1;
      patterns[26022] = 25'b01100101_10100100_00001001_1;
      patterns[26023] = 25'b01100101_10100101_00001010_1;
      patterns[26024] = 25'b01100101_10100110_00001011_1;
      patterns[26025] = 25'b01100101_10100111_00001100_1;
      patterns[26026] = 25'b01100101_10101000_00001101_1;
      patterns[26027] = 25'b01100101_10101001_00001110_1;
      patterns[26028] = 25'b01100101_10101010_00001111_1;
      patterns[26029] = 25'b01100101_10101011_00010000_1;
      patterns[26030] = 25'b01100101_10101100_00010001_1;
      patterns[26031] = 25'b01100101_10101101_00010010_1;
      patterns[26032] = 25'b01100101_10101110_00010011_1;
      patterns[26033] = 25'b01100101_10101111_00010100_1;
      patterns[26034] = 25'b01100101_10110000_00010101_1;
      patterns[26035] = 25'b01100101_10110001_00010110_1;
      patterns[26036] = 25'b01100101_10110010_00010111_1;
      patterns[26037] = 25'b01100101_10110011_00011000_1;
      patterns[26038] = 25'b01100101_10110100_00011001_1;
      patterns[26039] = 25'b01100101_10110101_00011010_1;
      patterns[26040] = 25'b01100101_10110110_00011011_1;
      patterns[26041] = 25'b01100101_10110111_00011100_1;
      patterns[26042] = 25'b01100101_10111000_00011101_1;
      patterns[26043] = 25'b01100101_10111001_00011110_1;
      patterns[26044] = 25'b01100101_10111010_00011111_1;
      patterns[26045] = 25'b01100101_10111011_00100000_1;
      patterns[26046] = 25'b01100101_10111100_00100001_1;
      patterns[26047] = 25'b01100101_10111101_00100010_1;
      patterns[26048] = 25'b01100101_10111110_00100011_1;
      patterns[26049] = 25'b01100101_10111111_00100100_1;
      patterns[26050] = 25'b01100101_11000000_00100101_1;
      patterns[26051] = 25'b01100101_11000001_00100110_1;
      patterns[26052] = 25'b01100101_11000010_00100111_1;
      patterns[26053] = 25'b01100101_11000011_00101000_1;
      patterns[26054] = 25'b01100101_11000100_00101001_1;
      patterns[26055] = 25'b01100101_11000101_00101010_1;
      patterns[26056] = 25'b01100101_11000110_00101011_1;
      patterns[26057] = 25'b01100101_11000111_00101100_1;
      patterns[26058] = 25'b01100101_11001000_00101101_1;
      patterns[26059] = 25'b01100101_11001001_00101110_1;
      patterns[26060] = 25'b01100101_11001010_00101111_1;
      patterns[26061] = 25'b01100101_11001011_00110000_1;
      patterns[26062] = 25'b01100101_11001100_00110001_1;
      patterns[26063] = 25'b01100101_11001101_00110010_1;
      patterns[26064] = 25'b01100101_11001110_00110011_1;
      patterns[26065] = 25'b01100101_11001111_00110100_1;
      patterns[26066] = 25'b01100101_11010000_00110101_1;
      patterns[26067] = 25'b01100101_11010001_00110110_1;
      patterns[26068] = 25'b01100101_11010010_00110111_1;
      patterns[26069] = 25'b01100101_11010011_00111000_1;
      patterns[26070] = 25'b01100101_11010100_00111001_1;
      patterns[26071] = 25'b01100101_11010101_00111010_1;
      patterns[26072] = 25'b01100101_11010110_00111011_1;
      patterns[26073] = 25'b01100101_11010111_00111100_1;
      patterns[26074] = 25'b01100101_11011000_00111101_1;
      patterns[26075] = 25'b01100101_11011001_00111110_1;
      patterns[26076] = 25'b01100101_11011010_00111111_1;
      patterns[26077] = 25'b01100101_11011011_01000000_1;
      patterns[26078] = 25'b01100101_11011100_01000001_1;
      patterns[26079] = 25'b01100101_11011101_01000010_1;
      patterns[26080] = 25'b01100101_11011110_01000011_1;
      patterns[26081] = 25'b01100101_11011111_01000100_1;
      patterns[26082] = 25'b01100101_11100000_01000101_1;
      patterns[26083] = 25'b01100101_11100001_01000110_1;
      patterns[26084] = 25'b01100101_11100010_01000111_1;
      patterns[26085] = 25'b01100101_11100011_01001000_1;
      patterns[26086] = 25'b01100101_11100100_01001001_1;
      patterns[26087] = 25'b01100101_11100101_01001010_1;
      patterns[26088] = 25'b01100101_11100110_01001011_1;
      patterns[26089] = 25'b01100101_11100111_01001100_1;
      patterns[26090] = 25'b01100101_11101000_01001101_1;
      patterns[26091] = 25'b01100101_11101001_01001110_1;
      patterns[26092] = 25'b01100101_11101010_01001111_1;
      patterns[26093] = 25'b01100101_11101011_01010000_1;
      patterns[26094] = 25'b01100101_11101100_01010001_1;
      patterns[26095] = 25'b01100101_11101101_01010010_1;
      patterns[26096] = 25'b01100101_11101110_01010011_1;
      patterns[26097] = 25'b01100101_11101111_01010100_1;
      patterns[26098] = 25'b01100101_11110000_01010101_1;
      patterns[26099] = 25'b01100101_11110001_01010110_1;
      patterns[26100] = 25'b01100101_11110010_01010111_1;
      patterns[26101] = 25'b01100101_11110011_01011000_1;
      patterns[26102] = 25'b01100101_11110100_01011001_1;
      patterns[26103] = 25'b01100101_11110101_01011010_1;
      patterns[26104] = 25'b01100101_11110110_01011011_1;
      patterns[26105] = 25'b01100101_11110111_01011100_1;
      patterns[26106] = 25'b01100101_11111000_01011101_1;
      patterns[26107] = 25'b01100101_11111001_01011110_1;
      patterns[26108] = 25'b01100101_11111010_01011111_1;
      patterns[26109] = 25'b01100101_11111011_01100000_1;
      patterns[26110] = 25'b01100101_11111100_01100001_1;
      patterns[26111] = 25'b01100101_11111101_01100010_1;
      patterns[26112] = 25'b01100101_11111110_01100011_1;
      patterns[26113] = 25'b01100101_11111111_01100100_1;
      patterns[26114] = 25'b01100110_00000000_01100110_0;
      patterns[26115] = 25'b01100110_00000001_01100111_0;
      patterns[26116] = 25'b01100110_00000010_01101000_0;
      patterns[26117] = 25'b01100110_00000011_01101001_0;
      patterns[26118] = 25'b01100110_00000100_01101010_0;
      patterns[26119] = 25'b01100110_00000101_01101011_0;
      patterns[26120] = 25'b01100110_00000110_01101100_0;
      patterns[26121] = 25'b01100110_00000111_01101101_0;
      patterns[26122] = 25'b01100110_00001000_01101110_0;
      patterns[26123] = 25'b01100110_00001001_01101111_0;
      patterns[26124] = 25'b01100110_00001010_01110000_0;
      patterns[26125] = 25'b01100110_00001011_01110001_0;
      patterns[26126] = 25'b01100110_00001100_01110010_0;
      patterns[26127] = 25'b01100110_00001101_01110011_0;
      patterns[26128] = 25'b01100110_00001110_01110100_0;
      patterns[26129] = 25'b01100110_00001111_01110101_0;
      patterns[26130] = 25'b01100110_00010000_01110110_0;
      patterns[26131] = 25'b01100110_00010001_01110111_0;
      patterns[26132] = 25'b01100110_00010010_01111000_0;
      patterns[26133] = 25'b01100110_00010011_01111001_0;
      patterns[26134] = 25'b01100110_00010100_01111010_0;
      patterns[26135] = 25'b01100110_00010101_01111011_0;
      patterns[26136] = 25'b01100110_00010110_01111100_0;
      patterns[26137] = 25'b01100110_00010111_01111101_0;
      patterns[26138] = 25'b01100110_00011000_01111110_0;
      patterns[26139] = 25'b01100110_00011001_01111111_0;
      patterns[26140] = 25'b01100110_00011010_10000000_0;
      patterns[26141] = 25'b01100110_00011011_10000001_0;
      patterns[26142] = 25'b01100110_00011100_10000010_0;
      patterns[26143] = 25'b01100110_00011101_10000011_0;
      patterns[26144] = 25'b01100110_00011110_10000100_0;
      patterns[26145] = 25'b01100110_00011111_10000101_0;
      patterns[26146] = 25'b01100110_00100000_10000110_0;
      patterns[26147] = 25'b01100110_00100001_10000111_0;
      patterns[26148] = 25'b01100110_00100010_10001000_0;
      patterns[26149] = 25'b01100110_00100011_10001001_0;
      patterns[26150] = 25'b01100110_00100100_10001010_0;
      patterns[26151] = 25'b01100110_00100101_10001011_0;
      patterns[26152] = 25'b01100110_00100110_10001100_0;
      patterns[26153] = 25'b01100110_00100111_10001101_0;
      patterns[26154] = 25'b01100110_00101000_10001110_0;
      patterns[26155] = 25'b01100110_00101001_10001111_0;
      patterns[26156] = 25'b01100110_00101010_10010000_0;
      patterns[26157] = 25'b01100110_00101011_10010001_0;
      patterns[26158] = 25'b01100110_00101100_10010010_0;
      patterns[26159] = 25'b01100110_00101101_10010011_0;
      patterns[26160] = 25'b01100110_00101110_10010100_0;
      patterns[26161] = 25'b01100110_00101111_10010101_0;
      patterns[26162] = 25'b01100110_00110000_10010110_0;
      patterns[26163] = 25'b01100110_00110001_10010111_0;
      patterns[26164] = 25'b01100110_00110010_10011000_0;
      patterns[26165] = 25'b01100110_00110011_10011001_0;
      patterns[26166] = 25'b01100110_00110100_10011010_0;
      patterns[26167] = 25'b01100110_00110101_10011011_0;
      patterns[26168] = 25'b01100110_00110110_10011100_0;
      patterns[26169] = 25'b01100110_00110111_10011101_0;
      patterns[26170] = 25'b01100110_00111000_10011110_0;
      patterns[26171] = 25'b01100110_00111001_10011111_0;
      patterns[26172] = 25'b01100110_00111010_10100000_0;
      patterns[26173] = 25'b01100110_00111011_10100001_0;
      patterns[26174] = 25'b01100110_00111100_10100010_0;
      patterns[26175] = 25'b01100110_00111101_10100011_0;
      patterns[26176] = 25'b01100110_00111110_10100100_0;
      patterns[26177] = 25'b01100110_00111111_10100101_0;
      patterns[26178] = 25'b01100110_01000000_10100110_0;
      patterns[26179] = 25'b01100110_01000001_10100111_0;
      patterns[26180] = 25'b01100110_01000010_10101000_0;
      patterns[26181] = 25'b01100110_01000011_10101001_0;
      patterns[26182] = 25'b01100110_01000100_10101010_0;
      patterns[26183] = 25'b01100110_01000101_10101011_0;
      patterns[26184] = 25'b01100110_01000110_10101100_0;
      patterns[26185] = 25'b01100110_01000111_10101101_0;
      patterns[26186] = 25'b01100110_01001000_10101110_0;
      patterns[26187] = 25'b01100110_01001001_10101111_0;
      patterns[26188] = 25'b01100110_01001010_10110000_0;
      patterns[26189] = 25'b01100110_01001011_10110001_0;
      patterns[26190] = 25'b01100110_01001100_10110010_0;
      patterns[26191] = 25'b01100110_01001101_10110011_0;
      patterns[26192] = 25'b01100110_01001110_10110100_0;
      patterns[26193] = 25'b01100110_01001111_10110101_0;
      patterns[26194] = 25'b01100110_01010000_10110110_0;
      patterns[26195] = 25'b01100110_01010001_10110111_0;
      patterns[26196] = 25'b01100110_01010010_10111000_0;
      patterns[26197] = 25'b01100110_01010011_10111001_0;
      patterns[26198] = 25'b01100110_01010100_10111010_0;
      patterns[26199] = 25'b01100110_01010101_10111011_0;
      patterns[26200] = 25'b01100110_01010110_10111100_0;
      patterns[26201] = 25'b01100110_01010111_10111101_0;
      patterns[26202] = 25'b01100110_01011000_10111110_0;
      patterns[26203] = 25'b01100110_01011001_10111111_0;
      patterns[26204] = 25'b01100110_01011010_11000000_0;
      patterns[26205] = 25'b01100110_01011011_11000001_0;
      patterns[26206] = 25'b01100110_01011100_11000010_0;
      patterns[26207] = 25'b01100110_01011101_11000011_0;
      patterns[26208] = 25'b01100110_01011110_11000100_0;
      patterns[26209] = 25'b01100110_01011111_11000101_0;
      patterns[26210] = 25'b01100110_01100000_11000110_0;
      patterns[26211] = 25'b01100110_01100001_11000111_0;
      patterns[26212] = 25'b01100110_01100010_11001000_0;
      patterns[26213] = 25'b01100110_01100011_11001001_0;
      patterns[26214] = 25'b01100110_01100100_11001010_0;
      patterns[26215] = 25'b01100110_01100101_11001011_0;
      patterns[26216] = 25'b01100110_01100110_11001100_0;
      patterns[26217] = 25'b01100110_01100111_11001101_0;
      patterns[26218] = 25'b01100110_01101000_11001110_0;
      patterns[26219] = 25'b01100110_01101001_11001111_0;
      patterns[26220] = 25'b01100110_01101010_11010000_0;
      patterns[26221] = 25'b01100110_01101011_11010001_0;
      patterns[26222] = 25'b01100110_01101100_11010010_0;
      patterns[26223] = 25'b01100110_01101101_11010011_0;
      patterns[26224] = 25'b01100110_01101110_11010100_0;
      patterns[26225] = 25'b01100110_01101111_11010101_0;
      patterns[26226] = 25'b01100110_01110000_11010110_0;
      patterns[26227] = 25'b01100110_01110001_11010111_0;
      patterns[26228] = 25'b01100110_01110010_11011000_0;
      patterns[26229] = 25'b01100110_01110011_11011001_0;
      patterns[26230] = 25'b01100110_01110100_11011010_0;
      patterns[26231] = 25'b01100110_01110101_11011011_0;
      patterns[26232] = 25'b01100110_01110110_11011100_0;
      patterns[26233] = 25'b01100110_01110111_11011101_0;
      patterns[26234] = 25'b01100110_01111000_11011110_0;
      patterns[26235] = 25'b01100110_01111001_11011111_0;
      patterns[26236] = 25'b01100110_01111010_11100000_0;
      patterns[26237] = 25'b01100110_01111011_11100001_0;
      patterns[26238] = 25'b01100110_01111100_11100010_0;
      patterns[26239] = 25'b01100110_01111101_11100011_0;
      patterns[26240] = 25'b01100110_01111110_11100100_0;
      patterns[26241] = 25'b01100110_01111111_11100101_0;
      patterns[26242] = 25'b01100110_10000000_11100110_0;
      patterns[26243] = 25'b01100110_10000001_11100111_0;
      patterns[26244] = 25'b01100110_10000010_11101000_0;
      patterns[26245] = 25'b01100110_10000011_11101001_0;
      patterns[26246] = 25'b01100110_10000100_11101010_0;
      patterns[26247] = 25'b01100110_10000101_11101011_0;
      patterns[26248] = 25'b01100110_10000110_11101100_0;
      patterns[26249] = 25'b01100110_10000111_11101101_0;
      patterns[26250] = 25'b01100110_10001000_11101110_0;
      patterns[26251] = 25'b01100110_10001001_11101111_0;
      patterns[26252] = 25'b01100110_10001010_11110000_0;
      patterns[26253] = 25'b01100110_10001011_11110001_0;
      patterns[26254] = 25'b01100110_10001100_11110010_0;
      patterns[26255] = 25'b01100110_10001101_11110011_0;
      patterns[26256] = 25'b01100110_10001110_11110100_0;
      patterns[26257] = 25'b01100110_10001111_11110101_0;
      patterns[26258] = 25'b01100110_10010000_11110110_0;
      patterns[26259] = 25'b01100110_10010001_11110111_0;
      patterns[26260] = 25'b01100110_10010010_11111000_0;
      patterns[26261] = 25'b01100110_10010011_11111001_0;
      patterns[26262] = 25'b01100110_10010100_11111010_0;
      patterns[26263] = 25'b01100110_10010101_11111011_0;
      patterns[26264] = 25'b01100110_10010110_11111100_0;
      patterns[26265] = 25'b01100110_10010111_11111101_0;
      patterns[26266] = 25'b01100110_10011000_11111110_0;
      patterns[26267] = 25'b01100110_10011001_11111111_0;
      patterns[26268] = 25'b01100110_10011010_00000000_1;
      patterns[26269] = 25'b01100110_10011011_00000001_1;
      patterns[26270] = 25'b01100110_10011100_00000010_1;
      patterns[26271] = 25'b01100110_10011101_00000011_1;
      patterns[26272] = 25'b01100110_10011110_00000100_1;
      patterns[26273] = 25'b01100110_10011111_00000101_1;
      patterns[26274] = 25'b01100110_10100000_00000110_1;
      patterns[26275] = 25'b01100110_10100001_00000111_1;
      patterns[26276] = 25'b01100110_10100010_00001000_1;
      patterns[26277] = 25'b01100110_10100011_00001001_1;
      patterns[26278] = 25'b01100110_10100100_00001010_1;
      patterns[26279] = 25'b01100110_10100101_00001011_1;
      patterns[26280] = 25'b01100110_10100110_00001100_1;
      patterns[26281] = 25'b01100110_10100111_00001101_1;
      patterns[26282] = 25'b01100110_10101000_00001110_1;
      patterns[26283] = 25'b01100110_10101001_00001111_1;
      patterns[26284] = 25'b01100110_10101010_00010000_1;
      patterns[26285] = 25'b01100110_10101011_00010001_1;
      patterns[26286] = 25'b01100110_10101100_00010010_1;
      patterns[26287] = 25'b01100110_10101101_00010011_1;
      patterns[26288] = 25'b01100110_10101110_00010100_1;
      patterns[26289] = 25'b01100110_10101111_00010101_1;
      patterns[26290] = 25'b01100110_10110000_00010110_1;
      patterns[26291] = 25'b01100110_10110001_00010111_1;
      patterns[26292] = 25'b01100110_10110010_00011000_1;
      patterns[26293] = 25'b01100110_10110011_00011001_1;
      patterns[26294] = 25'b01100110_10110100_00011010_1;
      patterns[26295] = 25'b01100110_10110101_00011011_1;
      patterns[26296] = 25'b01100110_10110110_00011100_1;
      patterns[26297] = 25'b01100110_10110111_00011101_1;
      patterns[26298] = 25'b01100110_10111000_00011110_1;
      patterns[26299] = 25'b01100110_10111001_00011111_1;
      patterns[26300] = 25'b01100110_10111010_00100000_1;
      patterns[26301] = 25'b01100110_10111011_00100001_1;
      patterns[26302] = 25'b01100110_10111100_00100010_1;
      patterns[26303] = 25'b01100110_10111101_00100011_1;
      patterns[26304] = 25'b01100110_10111110_00100100_1;
      patterns[26305] = 25'b01100110_10111111_00100101_1;
      patterns[26306] = 25'b01100110_11000000_00100110_1;
      patterns[26307] = 25'b01100110_11000001_00100111_1;
      patterns[26308] = 25'b01100110_11000010_00101000_1;
      patterns[26309] = 25'b01100110_11000011_00101001_1;
      patterns[26310] = 25'b01100110_11000100_00101010_1;
      patterns[26311] = 25'b01100110_11000101_00101011_1;
      patterns[26312] = 25'b01100110_11000110_00101100_1;
      patterns[26313] = 25'b01100110_11000111_00101101_1;
      patterns[26314] = 25'b01100110_11001000_00101110_1;
      patterns[26315] = 25'b01100110_11001001_00101111_1;
      patterns[26316] = 25'b01100110_11001010_00110000_1;
      patterns[26317] = 25'b01100110_11001011_00110001_1;
      patterns[26318] = 25'b01100110_11001100_00110010_1;
      patterns[26319] = 25'b01100110_11001101_00110011_1;
      patterns[26320] = 25'b01100110_11001110_00110100_1;
      patterns[26321] = 25'b01100110_11001111_00110101_1;
      patterns[26322] = 25'b01100110_11010000_00110110_1;
      patterns[26323] = 25'b01100110_11010001_00110111_1;
      patterns[26324] = 25'b01100110_11010010_00111000_1;
      patterns[26325] = 25'b01100110_11010011_00111001_1;
      patterns[26326] = 25'b01100110_11010100_00111010_1;
      patterns[26327] = 25'b01100110_11010101_00111011_1;
      patterns[26328] = 25'b01100110_11010110_00111100_1;
      patterns[26329] = 25'b01100110_11010111_00111101_1;
      patterns[26330] = 25'b01100110_11011000_00111110_1;
      patterns[26331] = 25'b01100110_11011001_00111111_1;
      patterns[26332] = 25'b01100110_11011010_01000000_1;
      patterns[26333] = 25'b01100110_11011011_01000001_1;
      patterns[26334] = 25'b01100110_11011100_01000010_1;
      patterns[26335] = 25'b01100110_11011101_01000011_1;
      patterns[26336] = 25'b01100110_11011110_01000100_1;
      patterns[26337] = 25'b01100110_11011111_01000101_1;
      patterns[26338] = 25'b01100110_11100000_01000110_1;
      patterns[26339] = 25'b01100110_11100001_01000111_1;
      patterns[26340] = 25'b01100110_11100010_01001000_1;
      patterns[26341] = 25'b01100110_11100011_01001001_1;
      patterns[26342] = 25'b01100110_11100100_01001010_1;
      patterns[26343] = 25'b01100110_11100101_01001011_1;
      patterns[26344] = 25'b01100110_11100110_01001100_1;
      patterns[26345] = 25'b01100110_11100111_01001101_1;
      patterns[26346] = 25'b01100110_11101000_01001110_1;
      patterns[26347] = 25'b01100110_11101001_01001111_1;
      patterns[26348] = 25'b01100110_11101010_01010000_1;
      patterns[26349] = 25'b01100110_11101011_01010001_1;
      patterns[26350] = 25'b01100110_11101100_01010010_1;
      patterns[26351] = 25'b01100110_11101101_01010011_1;
      patterns[26352] = 25'b01100110_11101110_01010100_1;
      patterns[26353] = 25'b01100110_11101111_01010101_1;
      patterns[26354] = 25'b01100110_11110000_01010110_1;
      patterns[26355] = 25'b01100110_11110001_01010111_1;
      patterns[26356] = 25'b01100110_11110010_01011000_1;
      patterns[26357] = 25'b01100110_11110011_01011001_1;
      patterns[26358] = 25'b01100110_11110100_01011010_1;
      patterns[26359] = 25'b01100110_11110101_01011011_1;
      patterns[26360] = 25'b01100110_11110110_01011100_1;
      patterns[26361] = 25'b01100110_11110111_01011101_1;
      patterns[26362] = 25'b01100110_11111000_01011110_1;
      patterns[26363] = 25'b01100110_11111001_01011111_1;
      patterns[26364] = 25'b01100110_11111010_01100000_1;
      patterns[26365] = 25'b01100110_11111011_01100001_1;
      patterns[26366] = 25'b01100110_11111100_01100010_1;
      patterns[26367] = 25'b01100110_11111101_01100011_1;
      patterns[26368] = 25'b01100110_11111110_01100100_1;
      patterns[26369] = 25'b01100110_11111111_01100101_1;
      patterns[26370] = 25'b01100111_00000000_01100111_0;
      patterns[26371] = 25'b01100111_00000001_01101000_0;
      patterns[26372] = 25'b01100111_00000010_01101001_0;
      patterns[26373] = 25'b01100111_00000011_01101010_0;
      patterns[26374] = 25'b01100111_00000100_01101011_0;
      patterns[26375] = 25'b01100111_00000101_01101100_0;
      patterns[26376] = 25'b01100111_00000110_01101101_0;
      patterns[26377] = 25'b01100111_00000111_01101110_0;
      patterns[26378] = 25'b01100111_00001000_01101111_0;
      patterns[26379] = 25'b01100111_00001001_01110000_0;
      patterns[26380] = 25'b01100111_00001010_01110001_0;
      patterns[26381] = 25'b01100111_00001011_01110010_0;
      patterns[26382] = 25'b01100111_00001100_01110011_0;
      patterns[26383] = 25'b01100111_00001101_01110100_0;
      patterns[26384] = 25'b01100111_00001110_01110101_0;
      patterns[26385] = 25'b01100111_00001111_01110110_0;
      patterns[26386] = 25'b01100111_00010000_01110111_0;
      patterns[26387] = 25'b01100111_00010001_01111000_0;
      patterns[26388] = 25'b01100111_00010010_01111001_0;
      patterns[26389] = 25'b01100111_00010011_01111010_0;
      patterns[26390] = 25'b01100111_00010100_01111011_0;
      patterns[26391] = 25'b01100111_00010101_01111100_0;
      patterns[26392] = 25'b01100111_00010110_01111101_0;
      patterns[26393] = 25'b01100111_00010111_01111110_0;
      patterns[26394] = 25'b01100111_00011000_01111111_0;
      patterns[26395] = 25'b01100111_00011001_10000000_0;
      patterns[26396] = 25'b01100111_00011010_10000001_0;
      patterns[26397] = 25'b01100111_00011011_10000010_0;
      patterns[26398] = 25'b01100111_00011100_10000011_0;
      patterns[26399] = 25'b01100111_00011101_10000100_0;
      patterns[26400] = 25'b01100111_00011110_10000101_0;
      patterns[26401] = 25'b01100111_00011111_10000110_0;
      patterns[26402] = 25'b01100111_00100000_10000111_0;
      patterns[26403] = 25'b01100111_00100001_10001000_0;
      patterns[26404] = 25'b01100111_00100010_10001001_0;
      patterns[26405] = 25'b01100111_00100011_10001010_0;
      patterns[26406] = 25'b01100111_00100100_10001011_0;
      patterns[26407] = 25'b01100111_00100101_10001100_0;
      patterns[26408] = 25'b01100111_00100110_10001101_0;
      patterns[26409] = 25'b01100111_00100111_10001110_0;
      patterns[26410] = 25'b01100111_00101000_10001111_0;
      patterns[26411] = 25'b01100111_00101001_10010000_0;
      patterns[26412] = 25'b01100111_00101010_10010001_0;
      patterns[26413] = 25'b01100111_00101011_10010010_0;
      patterns[26414] = 25'b01100111_00101100_10010011_0;
      patterns[26415] = 25'b01100111_00101101_10010100_0;
      patterns[26416] = 25'b01100111_00101110_10010101_0;
      patterns[26417] = 25'b01100111_00101111_10010110_0;
      patterns[26418] = 25'b01100111_00110000_10010111_0;
      patterns[26419] = 25'b01100111_00110001_10011000_0;
      patterns[26420] = 25'b01100111_00110010_10011001_0;
      patterns[26421] = 25'b01100111_00110011_10011010_0;
      patterns[26422] = 25'b01100111_00110100_10011011_0;
      patterns[26423] = 25'b01100111_00110101_10011100_0;
      patterns[26424] = 25'b01100111_00110110_10011101_0;
      patterns[26425] = 25'b01100111_00110111_10011110_0;
      patterns[26426] = 25'b01100111_00111000_10011111_0;
      patterns[26427] = 25'b01100111_00111001_10100000_0;
      patterns[26428] = 25'b01100111_00111010_10100001_0;
      patterns[26429] = 25'b01100111_00111011_10100010_0;
      patterns[26430] = 25'b01100111_00111100_10100011_0;
      patterns[26431] = 25'b01100111_00111101_10100100_0;
      patterns[26432] = 25'b01100111_00111110_10100101_0;
      patterns[26433] = 25'b01100111_00111111_10100110_0;
      patterns[26434] = 25'b01100111_01000000_10100111_0;
      patterns[26435] = 25'b01100111_01000001_10101000_0;
      patterns[26436] = 25'b01100111_01000010_10101001_0;
      patterns[26437] = 25'b01100111_01000011_10101010_0;
      patterns[26438] = 25'b01100111_01000100_10101011_0;
      patterns[26439] = 25'b01100111_01000101_10101100_0;
      patterns[26440] = 25'b01100111_01000110_10101101_0;
      patterns[26441] = 25'b01100111_01000111_10101110_0;
      patterns[26442] = 25'b01100111_01001000_10101111_0;
      patterns[26443] = 25'b01100111_01001001_10110000_0;
      patterns[26444] = 25'b01100111_01001010_10110001_0;
      patterns[26445] = 25'b01100111_01001011_10110010_0;
      patterns[26446] = 25'b01100111_01001100_10110011_0;
      patterns[26447] = 25'b01100111_01001101_10110100_0;
      patterns[26448] = 25'b01100111_01001110_10110101_0;
      patterns[26449] = 25'b01100111_01001111_10110110_0;
      patterns[26450] = 25'b01100111_01010000_10110111_0;
      patterns[26451] = 25'b01100111_01010001_10111000_0;
      patterns[26452] = 25'b01100111_01010010_10111001_0;
      patterns[26453] = 25'b01100111_01010011_10111010_0;
      patterns[26454] = 25'b01100111_01010100_10111011_0;
      patterns[26455] = 25'b01100111_01010101_10111100_0;
      patterns[26456] = 25'b01100111_01010110_10111101_0;
      patterns[26457] = 25'b01100111_01010111_10111110_0;
      patterns[26458] = 25'b01100111_01011000_10111111_0;
      patterns[26459] = 25'b01100111_01011001_11000000_0;
      patterns[26460] = 25'b01100111_01011010_11000001_0;
      patterns[26461] = 25'b01100111_01011011_11000010_0;
      patterns[26462] = 25'b01100111_01011100_11000011_0;
      patterns[26463] = 25'b01100111_01011101_11000100_0;
      patterns[26464] = 25'b01100111_01011110_11000101_0;
      patterns[26465] = 25'b01100111_01011111_11000110_0;
      patterns[26466] = 25'b01100111_01100000_11000111_0;
      patterns[26467] = 25'b01100111_01100001_11001000_0;
      patterns[26468] = 25'b01100111_01100010_11001001_0;
      patterns[26469] = 25'b01100111_01100011_11001010_0;
      patterns[26470] = 25'b01100111_01100100_11001011_0;
      patterns[26471] = 25'b01100111_01100101_11001100_0;
      patterns[26472] = 25'b01100111_01100110_11001101_0;
      patterns[26473] = 25'b01100111_01100111_11001110_0;
      patterns[26474] = 25'b01100111_01101000_11001111_0;
      patterns[26475] = 25'b01100111_01101001_11010000_0;
      patterns[26476] = 25'b01100111_01101010_11010001_0;
      patterns[26477] = 25'b01100111_01101011_11010010_0;
      patterns[26478] = 25'b01100111_01101100_11010011_0;
      patterns[26479] = 25'b01100111_01101101_11010100_0;
      patterns[26480] = 25'b01100111_01101110_11010101_0;
      patterns[26481] = 25'b01100111_01101111_11010110_0;
      patterns[26482] = 25'b01100111_01110000_11010111_0;
      patterns[26483] = 25'b01100111_01110001_11011000_0;
      patterns[26484] = 25'b01100111_01110010_11011001_0;
      patterns[26485] = 25'b01100111_01110011_11011010_0;
      patterns[26486] = 25'b01100111_01110100_11011011_0;
      patterns[26487] = 25'b01100111_01110101_11011100_0;
      patterns[26488] = 25'b01100111_01110110_11011101_0;
      patterns[26489] = 25'b01100111_01110111_11011110_0;
      patterns[26490] = 25'b01100111_01111000_11011111_0;
      patterns[26491] = 25'b01100111_01111001_11100000_0;
      patterns[26492] = 25'b01100111_01111010_11100001_0;
      patterns[26493] = 25'b01100111_01111011_11100010_0;
      patterns[26494] = 25'b01100111_01111100_11100011_0;
      patterns[26495] = 25'b01100111_01111101_11100100_0;
      patterns[26496] = 25'b01100111_01111110_11100101_0;
      patterns[26497] = 25'b01100111_01111111_11100110_0;
      patterns[26498] = 25'b01100111_10000000_11100111_0;
      patterns[26499] = 25'b01100111_10000001_11101000_0;
      patterns[26500] = 25'b01100111_10000010_11101001_0;
      patterns[26501] = 25'b01100111_10000011_11101010_0;
      patterns[26502] = 25'b01100111_10000100_11101011_0;
      patterns[26503] = 25'b01100111_10000101_11101100_0;
      patterns[26504] = 25'b01100111_10000110_11101101_0;
      patterns[26505] = 25'b01100111_10000111_11101110_0;
      patterns[26506] = 25'b01100111_10001000_11101111_0;
      patterns[26507] = 25'b01100111_10001001_11110000_0;
      patterns[26508] = 25'b01100111_10001010_11110001_0;
      patterns[26509] = 25'b01100111_10001011_11110010_0;
      patterns[26510] = 25'b01100111_10001100_11110011_0;
      patterns[26511] = 25'b01100111_10001101_11110100_0;
      patterns[26512] = 25'b01100111_10001110_11110101_0;
      patterns[26513] = 25'b01100111_10001111_11110110_0;
      patterns[26514] = 25'b01100111_10010000_11110111_0;
      patterns[26515] = 25'b01100111_10010001_11111000_0;
      patterns[26516] = 25'b01100111_10010010_11111001_0;
      patterns[26517] = 25'b01100111_10010011_11111010_0;
      patterns[26518] = 25'b01100111_10010100_11111011_0;
      patterns[26519] = 25'b01100111_10010101_11111100_0;
      patterns[26520] = 25'b01100111_10010110_11111101_0;
      patterns[26521] = 25'b01100111_10010111_11111110_0;
      patterns[26522] = 25'b01100111_10011000_11111111_0;
      patterns[26523] = 25'b01100111_10011001_00000000_1;
      patterns[26524] = 25'b01100111_10011010_00000001_1;
      patterns[26525] = 25'b01100111_10011011_00000010_1;
      patterns[26526] = 25'b01100111_10011100_00000011_1;
      patterns[26527] = 25'b01100111_10011101_00000100_1;
      patterns[26528] = 25'b01100111_10011110_00000101_1;
      patterns[26529] = 25'b01100111_10011111_00000110_1;
      patterns[26530] = 25'b01100111_10100000_00000111_1;
      patterns[26531] = 25'b01100111_10100001_00001000_1;
      patterns[26532] = 25'b01100111_10100010_00001001_1;
      patterns[26533] = 25'b01100111_10100011_00001010_1;
      patterns[26534] = 25'b01100111_10100100_00001011_1;
      patterns[26535] = 25'b01100111_10100101_00001100_1;
      patterns[26536] = 25'b01100111_10100110_00001101_1;
      patterns[26537] = 25'b01100111_10100111_00001110_1;
      patterns[26538] = 25'b01100111_10101000_00001111_1;
      patterns[26539] = 25'b01100111_10101001_00010000_1;
      patterns[26540] = 25'b01100111_10101010_00010001_1;
      patterns[26541] = 25'b01100111_10101011_00010010_1;
      patterns[26542] = 25'b01100111_10101100_00010011_1;
      patterns[26543] = 25'b01100111_10101101_00010100_1;
      patterns[26544] = 25'b01100111_10101110_00010101_1;
      patterns[26545] = 25'b01100111_10101111_00010110_1;
      patterns[26546] = 25'b01100111_10110000_00010111_1;
      patterns[26547] = 25'b01100111_10110001_00011000_1;
      patterns[26548] = 25'b01100111_10110010_00011001_1;
      patterns[26549] = 25'b01100111_10110011_00011010_1;
      patterns[26550] = 25'b01100111_10110100_00011011_1;
      patterns[26551] = 25'b01100111_10110101_00011100_1;
      patterns[26552] = 25'b01100111_10110110_00011101_1;
      patterns[26553] = 25'b01100111_10110111_00011110_1;
      patterns[26554] = 25'b01100111_10111000_00011111_1;
      patterns[26555] = 25'b01100111_10111001_00100000_1;
      patterns[26556] = 25'b01100111_10111010_00100001_1;
      patterns[26557] = 25'b01100111_10111011_00100010_1;
      patterns[26558] = 25'b01100111_10111100_00100011_1;
      patterns[26559] = 25'b01100111_10111101_00100100_1;
      patterns[26560] = 25'b01100111_10111110_00100101_1;
      patterns[26561] = 25'b01100111_10111111_00100110_1;
      patterns[26562] = 25'b01100111_11000000_00100111_1;
      patterns[26563] = 25'b01100111_11000001_00101000_1;
      patterns[26564] = 25'b01100111_11000010_00101001_1;
      patterns[26565] = 25'b01100111_11000011_00101010_1;
      patterns[26566] = 25'b01100111_11000100_00101011_1;
      patterns[26567] = 25'b01100111_11000101_00101100_1;
      patterns[26568] = 25'b01100111_11000110_00101101_1;
      patterns[26569] = 25'b01100111_11000111_00101110_1;
      patterns[26570] = 25'b01100111_11001000_00101111_1;
      patterns[26571] = 25'b01100111_11001001_00110000_1;
      patterns[26572] = 25'b01100111_11001010_00110001_1;
      patterns[26573] = 25'b01100111_11001011_00110010_1;
      patterns[26574] = 25'b01100111_11001100_00110011_1;
      patterns[26575] = 25'b01100111_11001101_00110100_1;
      patterns[26576] = 25'b01100111_11001110_00110101_1;
      patterns[26577] = 25'b01100111_11001111_00110110_1;
      patterns[26578] = 25'b01100111_11010000_00110111_1;
      patterns[26579] = 25'b01100111_11010001_00111000_1;
      patterns[26580] = 25'b01100111_11010010_00111001_1;
      patterns[26581] = 25'b01100111_11010011_00111010_1;
      patterns[26582] = 25'b01100111_11010100_00111011_1;
      patterns[26583] = 25'b01100111_11010101_00111100_1;
      patterns[26584] = 25'b01100111_11010110_00111101_1;
      patterns[26585] = 25'b01100111_11010111_00111110_1;
      patterns[26586] = 25'b01100111_11011000_00111111_1;
      patterns[26587] = 25'b01100111_11011001_01000000_1;
      patterns[26588] = 25'b01100111_11011010_01000001_1;
      patterns[26589] = 25'b01100111_11011011_01000010_1;
      patterns[26590] = 25'b01100111_11011100_01000011_1;
      patterns[26591] = 25'b01100111_11011101_01000100_1;
      patterns[26592] = 25'b01100111_11011110_01000101_1;
      patterns[26593] = 25'b01100111_11011111_01000110_1;
      patterns[26594] = 25'b01100111_11100000_01000111_1;
      patterns[26595] = 25'b01100111_11100001_01001000_1;
      patterns[26596] = 25'b01100111_11100010_01001001_1;
      patterns[26597] = 25'b01100111_11100011_01001010_1;
      patterns[26598] = 25'b01100111_11100100_01001011_1;
      patterns[26599] = 25'b01100111_11100101_01001100_1;
      patterns[26600] = 25'b01100111_11100110_01001101_1;
      patterns[26601] = 25'b01100111_11100111_01001110_1;
      patterns[26602] = 25'b01100111_11101000_01001111_1;
      patterns[26603] = 25'b01100111_11101001_01010000_1;
      patterns[26604] = 25'b01100111_11101010_01010001_1;
      patterns[26605] = 25'b01100111_11101011_01010010_1;
      patterns[26606] = 25'b01100111_11101100_01010011_1;
      patterns[26607] = 25'b01100111_11101101_01010100_1;
      patterns[26608] = 25'b01100111_11101110_01010101_1;
      patterns[26609] = 25'b01100111_11101111_01010110_1;
      patterns[26610] = 25'b01100111_11110000_01010111_1;
      patterns[26611] = 25'b01100111_11110001_01011000_1;
      patterns[26612] = 25'b01100111_11110010_01011001_1;
      patterns[26613] = 25'b01100111_11110011_01011010_1;
      patterns[26614] = 25'b01100111_11110100_01011011_1;
      patterns[26615] = 25'b01100111_11110101_01011100_1;
      patterns[26616] = 25'b01100111_11110110_01011101_1;
      patterns[26617] = 25'b01100111_11110111_01011110_1;
      patterns[26618] = 25'b01100111_11111000_01011111_1;
      patterns[26619] = 25'b01100111_11111001_01100000_1;
      patterns[26620] = 25'b01100111_11111010_01100001_1;
      patterns[26621] = 25'b01100111_11111011_01100010_1;
      patterns[26622] = 25'b01100111_11111100_01100011_1;
      patterns[26623] = 25'b01100111_11111101_01100100_1;
      patterns[26624] = 25'b01100111_11111110_01100101_1;
      patterns[26625] = 25'b01100111_11111111_01100110_1;
      patterns[26626] = 25'b01101000_00000000_01101000_0;
      patterns[26627] = 25'b01101000_00000001_01101001_0;
      patterns[26628] = 25'b01101000_00000010_01101010_0;
      patterns[26629] = 25'b01101000_00000011_01101011_0;
      patterns[26630] = 25'b01101000_00000100_01101100_0;
      patterns[26631] = 25'b01101000_00000101_01101101_0;
      patterns[26632] = 25'b01101000_00000110_01101110_0;
      patterns[26633] = 25'b01101000_00000111_01101111_0;
      patterns[26634] = 25'b01101000_00001000_01110000_0;
      patterns[26635] = 25'b01101000_00001001_01110001_0;
      patterns[26636] = 25'b01101000_00001010_01110010_0;
      patterns[26637] = 25'b01101000_00001011_01110011_0;
      patterns[26638] = 25'b01101000_00001100_01110100_0;
      patterns[26639] = 25'b01101000_00001101_01110101_0;
      patterns[26640] = 25'b01101000_00001110_01110110_0;
      patterns[26641] = 25'b01101000_00001111_01110111_0;
      patterns[26642] = 25'b01101000_00010000_01111000_0;
      patterns[26643] = 25'b01101000_00010001_01111001_0;
      patterns[26644] = 25'b01101000_00010010_01111010_0;
      patterns[26645] = 25'b01101000_00010011_01111011_0;
      patterns[26646] = 25'b01101000_00010100_01111100_0;
      patterns[26647] = 25'b01101000_00010101_01111101_0;
      patterns[26648] = 25'b01101000_00010110_01111110_0;
      patterns[26649] = 25'b01101000_00010111_01111111_0;
      patterns[26650] = 25'b01101000_00011000_10000000_0;
      patterns[26651] = 25'b01101000_00011001_10000001_0;
      patterns[26652] = 25'b01101000_00011010_10000010_0;
      patterns[26653] = 25'b01101000_00011011_10000011_0;
      patterns[26654] = 25'b01101000_00011100_10000100_0;
      patterns[26655] = 25'b01101000_00011101_10000101_0;
      patterns[26656] = 25'b01101000_00011110_10000110_0;
      patterns[26657] = 25'b01101000_00011111_10000111_0;
      patterns[26658] = 25'b01101000_00100000_10001000_0;
      patterns[26659] = 25'b01101000_00100001_10001001_0;
      patterns[26660] = 25'b01101000_00100010_10001010_0;
      patterns[26661] = 25'b01101000_00100011_10001011_0;
      patterns[26662] = 25'b01101000_00100100_10001100_0;
      patterns[26663] = 25'b01101000_00100101_10001101_0;
      patterns[26664] = 25'b01101000_00100110_10001110_0;
      patterns[26665] = 25'b01101000_00100111_10001111_0;
      patterns[26666] = 25'b01101000_00101000_10010000_0;
      patterns[26667] = 25'b01101000_00101001_10010001_0;
      patterns[26668] = 25'b01101000_00101010_10010010_0;
      patterns[26669] = 25'b01101000_00101011_10010011_0;
      patterns[26670] = 25'b01101000_00101100_10010100_0;
      patterns[26671] = 25'b01101000_00101101_10010101_0;
      patterns[26672] = 25'b01101000_00101110_10010110_0;
      patterns[26673] = 25'b01101000_00101111_10010111_0;
      patterns[26674] = 25'b01101000_00110000_10011000_0;
      patterns[26675] = 25'b01101000_00110001_10011001_0;
      patterns[26676] = 25'b01101000_00110010_10011010_0;
      patterns[26677] = 25'b01101000_00110011_10011011_0;
      patterns[26678] = 25'b01101000_00110100_10011100_0;
      patterns[26679] = 25'b01101000_00110101_10011101_0;
      patterns[26680] = 25'b01101000_00110110_10011110_0;
      patterns[26681] = 25'b01101000_00110111_10011111_0;
      patterns[26682] = 25'b01101000_00111000_10100000_0;
      patterns[26683] = 25'b01101000_00111001_10100001_0;
      patterns[26684] = 25'b01101000_00111010_10100010_0;
      patterns[26685] = 25'b01101000_00111011_10100011_0;
      patterns[26686] = 25'b01101000_00111100_10100100_0;
      patterns[26687] = 25'b01101000_00111101_10100101_0;
      patterns[26688] = 25'b01101000_00111110_10100110_0;
      patterns[26689] = 25'b01101000_00111111_10100111_0;
      patterns[26690] = 25'b01101000_01000000_10101000_0;
      patterns[26691] = 25'b01101000_01000001_10101001_0;
      patterns[26692] = 25'b01101000_01000010_10101010_0;
      patterns[26693] = 25'b01101000_01000011_10101011_0;
      patterns[26694] = 25'b01101000_01000100_10101100_0;
      patterns[26695] = 25'b01101000_01000101_10101101_0;
      patterns[26696] = 25'b01101000_01000110_10101110_0;
      patterns[26697] = 25'b01101000_01000111_10101111_0;
      patterns[26698] = 25'b01101000_01001000_10110000_0;
      patterns[26699] = 25'b01101000_01001001_10110001_0;
      patterns[26700] = 25'b01101000_01001010_10110010_0;
      patterns[26701] = 25'b01101000_01001011_10110011_0;
      patterns[26702] = 25'b01101000_01001100_10110100_0;
      patterns[26703] = 25'b01101000_01001101_10110101_0;
      patterns[26704] = 25'b01101000_01001110_10110110_0;
      patterns[26705] = 25'b01101000_01001111_10110111_0;
      patterns[26706] = 25'b01101000_01010000_10111000_0;
      patterns[26707] = 25'b01101000_01010001_10111001_0;
      patterns[26708] = 25'b01101000_01010010_10111010_0;
      patterns[26709] = 25'b01101000_01010011_10111011_0;
      patterns[26710] = 25'b01101000_01010100_10111100_0;
      patterns[26711] = 25'b01101000_01010101_10111101_0;
      patterns[26712] = 25'b01101000_01010110_10111110_0;
      patterns[26713] = 25'b01101000_01010111_10111111_0;
      patterns[26714] = 25'b01101000_01011000_11000000_0;
      patterns[26715] = 25'b01101000_01011001_11000001_0;
      patterns[26716] = 25'b01101000_01011010_11000010_0;
      patterns[26717] = 25'b01101000_01011011_11000011_0;
      patterns[26718] = 25'b01101000_01011100_11000100_0;
      patterns[26719] = 25'b01101000_01011101_11000101_0;
      patterns[26720] = 25'b01101000_01011110_11000110_0;
      patterns[26721] = 25'b01101000_01011111_11000111_0;
      patterns[26722] = 25'b01101000_01100000_11001000_0;
      patterns[26723] = 25'b01101000_01100001_11001001_0;
      patterns[26724] = 25'b01101000_01100010_11001010_0;
      patterns[26725] = 25'b01101000_01100011_11001011_0;
      patterns[26726] = 25'b01101000_01100100_11001100_0;
      patterns[26727] = 25'b01101000_01100101_11001101_0;
      patterns[26728] = 25'b01101000_01100110_11001110_0;
      patterns[26729] = 25'b01101000_01100111_11001111_0;
      patterns[26730] = 25'b01101000_01101000_11010000_0;
      patterns[26731] = 25'b01101000_01101001_11010001_0;
      patterns[26732] = 25'b01101000_01101010_11010010_0;
      patterns[26733] = 25'b01101000_01101011_11010011_0;
      patterns[26734] = 25'b01101000_01101100_11010100_0;
      patterns[26735] = 25'b01101000_01101101_11010101_0;
      patterns[26736] = 25'b01101000_01101110_11010110_0;
      patterns[26737] = 25'b01101000_01101111_11010111_0;
      patterns[26738] = 25'b01101000_01110000_11011000_0;
      patterns[26739] = 25'b01101000_01110001_11011001_0;
      patterns[26740] = 25'b01101000_01110010_11011010_0;
      patterns[26741] = 25'b01101000_01110011_11011011_0;
      patterns[26742] = 25'b01101000_01110100_11011100_0;
      patterns[26743] = 25'b01101000_01110101_11011101_0;
      patterns[26744] = 25'b01101000_01110110_11011110_0;
      patterns[26745] = 25'b01101000_01110111_11011111_0;
      patterns[26746] = 25'b01101000_01111000_11100000_0;
      patterns[26747] = 25'b01101000_01111001_11100001_0;
      patterns[26748] = 25'b01101000_01111010_11100010_0;
      patterns[26749] = 25'b01101000_01111011_11100011_0;
      patterns[26750] = 25'b01101000_01111100_11100100_0;
      patterns[26751] = 25'b01101000_01111101_11100101_0;
      patterns[26752] = 25'b01101000_01111110_11100110_0;
      patterns[26753] = 25'b01101000_01111111_11100111_0;
      patterns[26754] = 25'b01101000_10000000_11101000_0;
      patterns[26755] = 25'b01101000_10000001_11101001_0;
      patterns[26756] = 25'b01101000_10000010_11101010_0;
      patterns[26757] = 25'b01101000_10000011_11101011_0;
      patterns[26758] = 25'b01101000_10000100_11101100_0;
      patterns[26759] = 25'b01101000_10000101_11101101_0;
      patterns[26760] = 25'b01101000_10000110_11101110_0;
      patterns[26761] = 25'b01101000_10000111_11101111_0;
      patterns[26762] = 25'b01101000_10001000_11110000_0;
      patterns[26763] = 25'b01101000_10001001_11110001_0;
      patterns[26764] = 25'b01101000_10001010_11110010_0;
      patterns[26765] = 25'b01101000_10001011_11110011_0;
      patterns[26766] = 25'b01101000_10001100_11110100_0;
      patterns[26767] = 25'b01101000_10001101_11110101_0;
      patterns[26768] = 25'b01101000_10001110_11110110_0;
      patterns[26769] = 25'b01101000_10001111_11110111_0;
      patterns[26770] = 25'b01101000_10010000_11111000_0;
      patterns[26771] = 25'b01101000_10010001_11111001_0;
      patterns[26772] = 25'b01101000_10010010_11111010_0;
      patterns[26773] = 25'b01101000_10010011_11111011_0;
      patterns[26774] = 25'b01101000_10010100_11111100_0;
      patterns[26775] = 25'b01101000_10010101_11111101_0;
      patterns[26776] = 25'b01101000_10010110_11111110_0;
      patterns[26777] = 25'b01101000_10010111_11111111_0;
      patterns[26778] = 25'b01101000_10011000_00000000_1;
      patterns[26779] = 25'b01101000_10011001_00000001_1;
      patterns[26780] = 25'b01101000_10011010_00000010_1;
      patterns[26781] = 25'b01101000_10011011_00000011_1;
      patterns[26782] = 25'b01101000_10011100_00000100_1;
      patterns[26783] = 25'b01101000_10011101_00000101_1;
      patterns[26784] = 25'b01101000_10011110_00000110_1;
      patterns[26785] = 25'b01101000_10011111_00000111_1;
      patterns[26786] = 25'b01101000_10100000_00001000_1;
      patterns[26787] = 25'b01101000_10100001_00001001_1;
      patterns[26788] = 25'b01101000_10100010_00001010_1;
      patterns[26789] = 25'b01101000_10100011_00001011_1;
      patterns[26790] = 25'b01101000_10100100_00001100_1;
      patterns[26791] = 25'b01101000_10100101_00001101_1;
      patterns[26792] = 25'b01101000_10100110_00001110_1;
      patterns[26793] = 25'b01101000_10100111_00001111_1;
      patterns[26794] = 25'b01101000_10101000_00010000_1;
      patterns[26795] = 25'b01101000_10101001_00010001_1;
      patterns[26796] = 25'b01101000_10101010_00010010_1;
      patterns[26797] = 25'b01101000_10101011_00010011_1;
      patterns[26798] = 25'b01101000_10101100_00010100_1;
      patterns[26799] = 25'b01101000_10101101_00010101_1;
      patterns[26800] = 25'b01101000_10101110_00010110_1;
      patterns[26801] = 25'b01101000_10101111_00010111_1;
      patterns[26802] = 25'b01101000_10110000_00011000_1;
      patterns[26803] = 25'b01101000_10110001_00011001_1;
      patterns[26804] = 25'b01101000_10110010_00011010_1;
      patterns[26805] = 25'b01101000_10110011_00011011_1;
      patterns[26806] = 25'b01101000_10110100_00011100_1;
      patterns[26807] = 25'b01101000_10110101_00011101_1;
      patterns[26808] = 25'b01101000_10110110_00011110_1;
      patterns[26809] = 25'b01101000_10110111_00011111_1;
      patterns[26810] = 25'b01101000_10111000_00100000_1;
      patterns[26811] = 25'b01101000_10111001_00100001_1;
      patterns[26812] = 25'b01101000_10111010_00100010_1;
      patterns[26813] = 25'b01101000_10111011_00100011_1;
      patterns[26814] = 25'b01101000_10111100_00100100_1;
      patterns[26815] = 25'b01101000_10111101_00100101_1;
      patterns[26816] = 25'b01101000_10111110_00100110_1;
      patterns[26817] = 25'b01101000_10111111_00100111_1;
      patterns[26818] = 25'b01101000_11000000_00101000_1;
      patterns[26819] = 25'b01101000_11000001_00101001_1;
      patterns[26820] = 25'b01101000_11000010_00101010_1;
      patterns[26821] = 25'b01101000_11000011_00101011_1;
      patterns[26822] = 25'b01101000_11000100_00101100_1;
      patterns[26823] = 25'b01101000_11000101_00101101_1;
      patterns[26824] = 25'b01101000_11000110_00101110_1;
      patterns[26825] = 25'b01101000_11000111_00101111_1;
      patterns[26826] = 25'b01101000_11001000_00110000_1;
      patterns[26827] = 25'b01101000_11001001_00110001_1;
      patterns[26828] = 25'b01101000_11001010_00110010_1;
      patterns[26829] = 25'b01101000_11001011_00110011_1;
      patterns[26830] = 25'b01101000_11001100_00110100_1;
      patterns[26831] = 25'b01101000_11001101_00110101_1;
      patterns[26832] = 25'b01101000_11001110_00110110_1;
      patterns[26833] = 25'b01101000_11001111_00110111_1;
      patterns[26834] = 25'b01101000_11010000_00111000_1;
      patterns[26835] = 25'b01101000_11010001_00111001_1;
      patterns[26836] = 25'b01101000_11010010_00111010_1;
      patterns[26837] = 25'b01101000_11010011_00111011_1;
      patterns[26838] = 25'b01101000_11010100_00111100_1;
      patterns[26839] = 25'b01101000_11010101_00111101_1;
      patterns[26840] = 25'b01101000_11010110_00111110_1;
      patterns[26841] = 25'b01101000_11010111_00111111_1;
      patterns[26842] = 25'b01101000_11011000_01000000_1;
      patterns[26843] = 25'b01101000_11011001_01000001_1;
      patterns[26844] = 25'b01101000_11011010_01000010_1;
      patterns[26845] = 25'b01101000_11011011_01000011_1;
      patterns[26846] = 25'b01101000_11011100_01000100_1;
      patterns[26847] = 25'b01101000_11011101_01000101_1;
      patterns[26848] = 25'b01101000_11011110_01000110_1;
      patterns[26849] = 25'b01101000_11011111_01000111_1;
      patterns[26850] = 25'b01101000_11100000_01001000_1;
      patterns[26851] = 25'b01101000_11100001_01001001_1;
      patterns[26852] = 25'b01101000_11100010_01001010_1;
      patterns[26853] = 25'b01101000_11100011_01001011_1;
      patterns[26854] = 25'b01101000_11100100_01001100_1;
      patterns[26855] = 25'b01101000_11100101_01001101_1;
      patterns[26856] = 25'b01101000_11100110_01001110_1;
      patterns[26857] = 25'b01101000_11100111_01001111_1;
      patterns[26858] = 25'b01101000_11101000_01010000_1;
      patterns[26859] = 25'b01101000_11101001_01010001_1;
      patterns[26860] = 25'b01101000_11101010_01010010_1;
      patterns[26861] = 25'b01101000_11101011_01010011_1;
      patterns[26862] = 25'b01101000_11101100_01010100_1;
      patterns[26863] = 25'b01101000_11101101_01010101_1;
      patterns[26864] = 25'b01101000_11101110_01010110_1;
      patterns[26865] = 25'b01101000_11101111_01010111_1;
      patterns[26866] = 25'b01101000_11110000_01011000_1;
      patterns[26867] = 25'b01101000_11110001_01011001_1;
      patterns[26868] = 25'b01101000_11110010_01011010_1;
      patterns[26869] = 25'b01101000_11110011_01011011_1;
      patterns[26870] = 25'b01101000_11110100_01011100_1;
      patterns[26871] = 25'b01101000_11110101_01011101_1;
      patterns[26872] = 25'b01101000_11110110_01011110_1;
      patterns[26873] = 25'b01101000_11110111_01011111_1;
      patterns[26874] = 25'b01101000_11111000_01100000_1;
      patterns[26875] = 25'b01101000_11111001_01100001_1;
      patterns[26876] = 25'b01101000_11111010_01100010_1;
      patterns[26877] = 25'b01101000_11111011_01100011_1;
      patterns[26878] = 25'b01101000_11111100_01100100_1;
      patterns[26879] = 25'b01101000_11111101_01100101_1;
      patterns[26880] = 25'b01101000_11111110_01100110_1;
      patterns[26881] = 25'b01101000_11111111_01100111_1;
      patterns[26882] = 25'b01101001_00000000_01101001_0;
      patterns[26883] = 25'b01101001_00000001_01101010_0;
      patterns[26884] = 25'b01101001_00000010_01101011_0;
      patterns[26885] = 25'b01101001_00000011_01101100_0;
      patterns[26886] = 25'b01101001_00000100_01101101_0;
      patterns[26887] = 25'b01101001_00000101_01101110_0;
      patterns[26888] = 25'b01101001_00000110_01101111_0;
      patterns[26889] = 25'b01101001_00000111_01110000_0;
      patterns[26890] = 25'b01101001_00001000_01110001_0;
      patterns[26891] = 25'b01101001_00001001_01110010_0;
      patterns[26892] = 25'b01101001_00001010_01110011_0;
      patterns[26893] = 25'b01101001_00001011_01110100_0;
      patterns[26894] = 25'b01101001_00001100_01110101_0;
      patterns[26895] = 25'b01101001_00001101_01110110_0;
      patterns[26896] = 25'b01101001_00001110_01110111_0;
      patterns[26897] = 25'b01101001_00001111_01111000_0;
      patterns[26898] = 25'b01101001_00010000_01111001_0;
      patterns[26899] = 25'b01101001_00010001_01111010_0;
      patterns[26900] = 25'b01101001_00010010_01111011_0;
      patterns[26901] = 25'b01101001_00010011_01111100_0;
      patterns[26902] = 25'b01101001_00010100_01111101_0;
      patterns[26903] = 25'b01101001_00010101_01111110_0;
      patterns[26904] = 25'b01101001_00010110_01111111_0;
      patterns[26905] = 25'b01101001_00010111_10000000_0;
      patterns[26906] = 25'b01101001_00011000_10000001_0;
      patterns[26907] = 25'b01101001_00011001_10000010_0;
      patterns[26908] = 25'b01101001_00011010_10000011_0;
      patterns[26909] = 25'b01101001_00011011_10000100_0;
      patterns[26910] = 25'b01101001_00011100_10000101_0;
      patterns[26911] = 25'b01101001_00011101_10000110_0;
      patterns[26912] = 25'b01101001_00011110_10000111_0;
      patterns[26913] = 25'b01101001_00011111_10001000_0;
      patterns[26914] = 25'b01101001_00100000_10001001_0;
      patterns[26915] = 25'b01101001_00100001_10001010_0;
      patterns[26916] = 25'b01101001_00100010_10001011_0;
      patterns[26917] = 25'b01101001_00100011_10001100_0;
      patterns[26918] = 25'b01101001_00100100_10001101_0;
      patterns[26919] = 25'b01101001_00100101_10001110_0;
      patterns[26920] = 25'b01101001_00100110_10001111_0;
      patterns[26921] = 25'b01101001_00100111_10010000_0;
      patterns[26922] = 25'b01101001_00101000_10010001_0;
      patterns[26923] = 25'b01101001_00101001_10010010_0;
      patterns[26924] = 25'b01101001_00101010_10010011_0;
      patterns[26925] = 25'b01101001_00101011_10010100_0;
      patterns[26926] = 25'b01101001_00101100_10010101_0;
      patterns[26927] = 25'b01101001_00101101_10010110_0;
      patterns[26928] = 25'b01101001_00101110_10010111_0;
      patterns[26929] = 25'b01101001_00101111_10011000_0;
      patterns[26930] = 25'b01101001_00110000_10011001_0;
      patterns[26931] = 25'b01101001_00110001_10011010_0;
      patterns[26932] = 25'b01101001_00110010_10011011_0;
      patterns[26933] = 25'b01101001_00110011_10011100_0;
      patterns[26934] = 25'b01101001_00110100_10011101_0;
      patterns[26935] = 25'b01101001_00110101_10011110_0;
      patterns[26936] = 25'b01101001_00110110_10011111_0;
      patterns[26937] = 25'b01101001_00110111_10100000_0;
      patterns[26938] = 25'b01101001_00111000_10100001_0;
      patterns[26939] = 25'b01101001_00111001_10100010_0;
      patterns[26940] = 25'b01101001_00111010_10100011_0;
      patterns[26941] = 25'b01101001_00111011_10100100_0;
      patterns[26942] = 25'b01101001_00111100_10100101_0;
      patterns[26943] = 25'b01101001_00111101_10100110_0;
      patterns[26944] = 25'b01101001_00111110_10100111_0;
      patterns[26945] = 25'b01101001_00111111_10101000_0;
      patterns[26946] = 25'b01101001_01000000_10101001_0;
      patterns[26947] = 25'b01101001_01000001_10101010_0;
      patterns[26948] = 25'b01101001_01000010_10101011_0;
      patterns[26949] = 25'b01101001_01000011_10101100_0;
      patterns[26950] = 25'b01101001_01000100_10101101_0;
      patterns[26951] = 25'b01101001_01000101_10101110_0;
      patterns[26952] = 25'b01101001_01000110_10101111_0;
      patterns[26953] = 25'b01101001_01000111_10110000_0;
      patterns[26954] = 25'b01101001_01001000_10110001_0;
      patterns[26955] = 25'b01101001_01001001_10110010_0;
      patterns[26956] = 25'b01101001_01001010_10110011_0;
      patterns[26957] = 25'b01101001_01001011_10110100_0;
      patterns[26958] = 25'b01101001_01001100_10110101_0;
      patterns[26959] = 25'b01101001_01001101_10110110_0;
      patterns[26960] = 25'b01101001_01001110_10110111_0;
      patterns[26961] = 25'b01101001_01001111_10111000_0;
      patterns[26962] = 25'b01101001_01010000_10111001_0;
      patterns[26963] = 25'b01101001_01010001_10111010_0;
      patterns[26964] = 25'b01101001_01010010_10111011_0;
      patterns[26965] = 25'b01101001_01010011_10111100_0;
      patterns[26966] = 25'b01101001_01010100_10111101_0;
      patterns[26967] = 25'b01101001_01010101_10111110_0;
      patterns[26968] = 25'b01101001_01010110_10111111_0;
      patterns[26969] = 25'b01101001_01010111_11000000_0;
      patterns[26970] = 25'b01101001_01011000_11000001_0;
      patterns[26971] = 25'b01101001_01011001_11000010_0;
      patterns[26972] = 25'b01101001_01011010_11000011_0;
      patterns[26973] = 25'b01101001_01011011_11000100_0;
      patterns[26974] = 25'b01101001_01011100_11000101_0;
      patterns[26975] = 25'b01101001_01011101_11000110_0;
      patterns[26976] = 25'b01101001_01011110_11000111_0;
      patterns[26977] = 25'b01101001_01011111_11001000_0;
      patterns[26978] = 25'b01101001_01100000_11001001_0;
      patterns[26979] = 25'b01101001_01100001_11001010_0;
      patterns[26980] = 25'b01101001_01100010_11001011_0;
      patterns[26981] = 25'b01101001_01100011_11001100_0;
      patterns[26982] = 25'b01101001_01100100_11001101_0;
      patterns[26983] = 25'b01101001_01100101_11001110_0;
      patterns[26984] = 25'b01101001_01100110_11001111_0;
      patterns[26985] = 25'b01101001_01100111_11010000_0;
      patterns[26986] = 25'b01101001_01101000_11010001_0;
      patterns[26987] = 25'b01101001_01101001_11010010_0;
      patterns[26988] = 25'b01101001_01101010_11010011_0;
      patterns[26989] = 25'b01101001_01101011_11010100_0;
      patterns[26990] = 25'b01101001_01101100_11010101_0;
      patterns[26991] = 25'b01101001_01101101_11010110_0;
      patterns[26992] = 25'b01101001_01101110_11010111_0;
      patterns[26993] = 25'b01101001_01101111_11011000_0;
      patterns[26994] = 25'b01101001_01110000_11011001_0;
      patterns[26995] = 25'b01101001_01110001_11011010_0;
      patterns[26996] = 25'b01101001_01110010_11011011_0;
      patterns[26997] = 25'b01101001_01110011_11011100_0;
      patterns[26998] = 25'b01101001_01110100_11011101_0;
      patterns[26999] = 25'b01101001_01110101_11011110_0;
      patterns[27000] = 25'b01101001_01110110_11011111_0;
      patterns[27001] = 25'b01101001_01110111_11100000_0;
      patterns[27002] = 25'b01101001_01111000_11100001_0;
      patterns[27003] = 25'b01101001_01111001_11100010_0;
      patterns[27004] = 25'b01101001_01111010_11100011_0;
      patterns[27005] = 25'b01101001_01111011_11100100_0;
      patterns[27006] = 25'b01101001_01111100_11100101_0;
      patterns[27007] = 25'b01101001_01111101_11100110_0;
      patterns[27008] = 25'b01101001_01111110_11100111_0;
      patterns[27009] = 25'b01101001_01111111_11101000_0;
      patterns[27010] = 25'b01101001_10000000_11101001_0;
      patterns[27011] = 25'b01101001_10000001_11101010_0;
      patterns[27012] = 25'b01101001_10000010_11101011_0;
      patterns[27013] = 25'b01101001_10000011_11101100_0;
      patterns[27014] = 25'b01101001_10000100_11101101_0;
      patterns[27015] = 25'b01101001_10000101_11101110_0;
      patterns[27016] = 25'b01101001_10000110_11101111_0;
      patterns[27017] = 25'b01101001_10000111_11110000_0;
      patterns[27018] = 25'b01101001_10001000_11110001_0;
      patterns[27019] = 25'b01101001_10001001_11110010_0;
      patterns[27020] = 25'b01101001_10001010_11110011_0;
      patterns[27021] = 25'b01101001_10001011_11110100_0;
      patterns[27022] = 25'b01101001_10001100_11110101_0;
      patterns[27023] = 25'b01101001_10001101_11110110_0;
      patterns[27024] = 25'b01101001_10001110_11110111_0;
      patterns[27025] = 25'b01101001_10001111_11111000_0;
      patterns[27026] = 25'b01101001_10010000_11111001_0;
      patterns[27027] = 25'b01101001_10010001_11111010_0;
      patterns[27028] = 25'b01101001_10010010_11111011_0;
      patterns[27029] = 25'b01101001_10010011_11111100_0;
      patterns[27030] = 25'b01101001_10010100_11111101_0;
      patterns[27031] = 25'b01101001_10010101_11111110_0;
      patterns[27032] = 25'b01101001_10010110_11111111_0;
      patterns[27033] = 25'b01101001_10010111_00000000_1;
      patterns[27034] = 25'b01101001_10011000_00000001_1;
      patterns[27035] = 25'b01101001_10011001_00000010_1;
      patterns[27036] = 25'b01101001_10011010_00000011_1;
      patterns[27037] = 25'b01101001_10011011_00000100_1;
      patterns[27038] = 25'b01101001_10011100_00000101_1;
      patterns[27039] = 25'b01101001_10011101_00000110_1;
      patterns[27040] = 25'b01101001_10011110_00000111_1;
      patterns[27041] = 25'b01101001_10011111_00001000_1;
      patterns[27042] = 25'b01101001_10100000_00001001_1;
      patterns[27043] = 25'b01101001_10100001_00001010_1;
      patterns[27044] = 25'b01101001_10100010_00001011_1;
      patterns[27045] = 25'b01101001_10100011_00001100_1;
      patterns[27046] = 25'b01101001_10100100_00001101_1;
      patterns[27047] = 25'b01101001_10100101_00001110_1;
      patterns[27048] = 25'b01101001_10100110_00001111_1;
      patterns[27049] = 25'b01101001_10100111_00010000_1;
      patterns[27050] = 25'b01101001_10101000_00010001_1;
      patterns[27051] = 25'b01101001_10101001_00010010_1;
      patterns[27052] = 25'b01101001_10101010_00010011_1;
      patterns[27053] = 25'b01101001_10101011_00010100_1;
      patterns[27054] = 25'b01101001_10101100_00010101_1;
      patterns[27055] = 25'b01101001_10101101_00010110_1;
      patterns[27056] = 25'b01101001_10101110_00010111_1;
      patterns[27057] = 25'b01101001_10101111_00011000_1;
      patterns[27058] = 25'b01101001_10110000_00011001_1;
      patterns[27059] = 25'b01101001_10110001_00011010_1;
      patterns[27060] = 25'b01101001_10110010_00011011_1;
      patterns[27061] = 25'b01101001_10110011_00011100_1;
      patterns[27062] = 25'b01101001_10110100_00011101_1;
      patterns[27063] = 25'b01101001_10110101_00011110_1;
      patterns[27064] = 25'b01101001_10110110_00011111_1;
      patterns[27065] = 25'b01101001_10110111_00100000_1;
      patterns[27066] = 25'b01101001_10111000_00100001_1;
      patterns[27067] = 25'b01101001_10111001_00100010_1;
      patterns[27068] = 25'b01101001_10111010_00100011_1;
      patterns[27069] = 25'b01101001_10111011_00100100_1;
      patterns[27070] = 25'b01101001_10111100_00100101_1;
      patterns[27071] = 25'b01101001_10111101_00100110_1;
      patterns[27072] = 25'b01101001_10111110_00100111_1;
      patterns[27073] = 25'b01101001_10111111_00101000_1;
      patterns[27074] = 25'b01101001_11000000_00101001_1;
      patterns[27075] = 25'b01101001_11000001_00101010_1;
      patterns[27076] = 25'b01101001_11000010_00101011_1;
      patterns[27077] = 25'b01101001_11000011_00101100_1;
      patterns[27078] = 25'b01101001_11000100_00101101_1;
      patterns[27079] = 25'b01101001_11000101_00101110_1;
      patterns[27080] = 25'b01101001_11000110_00101111_1;
      patterns[27081] = 25'b01101001_11000111_00110000_1;
      patterns[27082] = 25'b01101001_11001000_00110001_1;
      patterns[27083] = 25'b01101001_11001001_00110010_1;
      patterns[27084] = 25'b01101001_11001010_00110011_1;
      patterns[27085] = 25'b01101001_11001011_00110100_1;
      patterns[27086] = 25'b01101001_11001100_00110101_1;
      patterns[27087] = 25'b01101001_11001101_00110110_1;
      patterns[27088] = 25'b01101001_11001110_00110111_1;
      patterns[27089] = 25'b01101001_11001111_00111000_1;
      patterns[27090] = 25'b01101001_11010000_00111001_1;
      patterns[27091] = 25'b01101001_11010001_00111010_1;
      patterns[27092] = 25'b01101001_11010010_00111011_1;
      patterns[27093] = 25'b01101001_11010011_00111100_1;
      patterns[27094] = 25'b01101001_11010100_00111101_1;
      patterns[27095] = 25'b01101001_11010101_00111110_1;
      patterns[27096] = 25'b01101001_11010110_00111111_1;
      patterns[27097] = 25'b01101001_11010111_01000000_1;
      patterns[27098] = 25'b01101001_11011000_01000001_1;
      patterns[27099] = 25'b01101001_11011001_01000010_1;
      patterns[27100] = 25'b01101001_11011010_01000011_1;
      patterns[27101] = 25'b01101001_11011011_01000100_1;
      patterns[27102] = 25'b01101001_11011100_01000101_1;
      patterns[27103] = 25'b01101001_11011101_01000110_1;
      patterns[27104] = 25'b01101001_11011110_01000111_1;
      patterns[27105] = 25'b01101001_11011111_01001000_1;
      patterns[27106] = 25'b01101001_11100000_01001001_1;
      patterns[27107] = 25'b01101001_11100001_01001010_1;
      patterns[27108] = 25'b01101001_11100010_01001011_1;
      patterns[27109] = 25'b01101001_11100011_01001100_1;
      patterns[27110] = 25'b01101001_11100100_01001101_1;
      patterns[27111] = 25'b01101001_11100101_01001110_1;
      patterns[27112] = 25'b01101001_11100110_01001111_1;
      patterns[27113] = 25'b01101001_11100111_01010000_1;
      patterns[27114] = 25'b01101001_11101000_01010001_1;
      patterns[27115] = 25'b01101001_11101001_01010010_1;
      patterns[27116] = 25'b01101001_11101010_01010011_1;
      patterns[27117] = 25'b01101001_11101011_01010100_1;
      patterns[27118] = 25'b01101001_11101100_01010101_1;
      patterns[27119] = 25'b01101001_11101101_01010110_1;
      patterns[27120] = 25'b01101001_11101110_01010111_1;
      patterns[27121] = 25'b01101001_11101111_01011000_1;
      patterns[27122] = 25'b01101001_11110000_01011001_1;
      patterns[27123] = 25'b01101001_11110001_01011010_1;
      patterns[27124] = 25'b01101001_11110010_01011011_1;
      patterns[27125] = 25'b01101001_11110011_01011100_1;
      patterns[27126] = 25'b01101001_11110100_01011101_1;
      patterns[27127] = 25'b01101001_11110101_01011110_1;
      patterns[27128] = 25'b01101001_11110110_01011111_1;
      patterns[27129] = 25'b01101001_11110111_01100000_1;
      patterns[27130] = 25'b01101001_11111000_01100001_1;
      patterns[27131] = 25'b01101001_11111001_01100010_1;
      patterns[27132] = 25'b01101001_11111010_01100011_1;
      patterns[27133] = 25'b01101001_11111011_01100100_1;
      patterns[27134] = 25'b01101001_11111100_01100101_1;
      patterns[27135] = 25'b01101001_11111101_01100110_1;
      patterns[27136] = 25'b01101001_11111110_01100111_1;
      patterns[27137] = 25'b01101001_11111111_01101000_1;
      patterns[27138] = 25'b01101010_00000000_01101010_0;
      patterns[27139] = 25'b01101010_00000001_01101011_0;
      patterns[27140] = 25'b01101010_00000010_01101100_0;
      patterns[27141] = 25'b01101010_00000011_01101101_0;
      patterns[27142] = 25'b01101010_00000100_01101110_0;
      patterns[27143] = 25'b01101010_00000101_01101111_0;
      patterns[27144] = 25'b01101010_00000110_01110000_0;
      patterns[27145] = 25'b01101010_00000111_01110001_0;
      patterns[27146] = 25'b01101010_00001000_01110010_0;
      patterns[27147] = 25'b01101010_00001001_01110011_0;
      patterns[27148] = 25'b01101010_00001010_01110100_0;
      patterns[27149] = 25'b01101010_00001011_01110101_0;
      patterns[27150] = 25'b01101010_00001100_01110110_0;
      patterns[27151] = 25'b01101010_00001101_01110111_0;
      patterns[27152] = 25'b01101010_00001110_01111000_0;
      patterns[27153] = 25'b01101010_00001111_01111001_0;
      patterns[27154] = 25'b01101010_00010000_01111010_0;
      patterns[27155] = 25'b01101010_00010001_01111011_0;
      patterns[27156] = 25'b01101010_00010010_01111100_0;
      patterns[27157] = 25'b01101010_00010011_01111101_0;
      patterns[27158] = 25'b01101010_00010100_01111110_0;
      patterns[27159] = 25'b01101010_00010101_01111111_0;
      patterns[27160] = 25'b01101010_00010110_10000000_0;
      patterns[27161] = 25'b01101010_00010111_10000001_0;
      patterns[27162] = 25'b01101010_00011000_10000010_0;
      patterns[27163] = 25'b01101010_00011001_10000011_0;
      patterns[27164] = 25'b01101010_00011010_10000100_0;
      patterns[27165] = 25'b01101010_00011011_10000101_0;
      patterns[27166] = 25'b01101010_00011100_10000110_0;
      patterns[27167] = 25'b01101010_00011101_10000111_0;
      patterns[27168] = 25'b01101010_00011110_10001000_0;
      patterns[27169] = 25'b01101010_00011111_10001001_0;
      patterns[27170] = 25'b01101010_00100000_10001010_0;
      patterns[27171] = 25'b01101010_00100001_10001011_0;
      patterns[27172] = 25'b01101010_00100010_10001100_0;
      patterns[27173] = 25'b01101010_00100011_10001101_0;
      patterns[27174] = 25'b01101010_00100100_10001110_0;
      patterns[27175] = 25'b01101010_00100101_10001111_0;
      patterns[27176] = 25'b01101010_00100110_10010000_0;
      patterns[27177] = 25'b01101010_00100111_10010001_0;
      patterns[27178] = 25'b01101010_00101000_10010010_0;
      patterns[27179] = 25'b01101010_00101001_10010011_0;
      patterns[27180] = 25'b01101010_00101010_10010100_0;
      patterns[27181] = 25'b01101010_00101011_10010101_0;
      patterns[27182] = 25'b01101010_00101100_10010110_0;
      patterns[27183] = 25'b01101010_00101101_10010111_0;
      patterns[27184] = 25'b01101010_00101110_10011000_0;
      patterns[27185] = 25'b01101010_00101111_10011001_0;
      patterns[27186] = 25'b01101010_00110000_10011010_0;
      patterns[27187] = 25'b01101010_00110001_10011011_0;
      patterns[27188] = 25'b01101010_00110010_10011100_0;
      patterns[27189] = 25'b01101010_00110011_10011101_0;
      patterns[27190] = 25'b01101010_00110100_10011110_0;
      patterns[27191] = 25'b01101010_00110101_10011111_0;
      patterns[27192] = 25'b01101010_00110110_10100000_0;
      patterns[27193] = 25'b01101010_00110111_10100001_0;
      patterns[27194] = 25'b01101010_00111000_10100010_0;
      patterns[27195] = 25'b01101010_00111001_10100011_0;
      patterns[27196] = 25'b01101010_00111010_10100100_0;
      patterns[27197] = 25'b01101010_00111011_10100101_0;
      patterns[27198] = 25'b01101010_00111100_10100110_0;
      patterns[27199] = 25'b01101010_00111101_10100111_0;
      patterns[27200] = 25'b01101010_00111110_10101000_0;
      patterns[27201] = 25'b01101010_00111111_10101001_0;
      patterns[27202] = 25'b01101010_01000000_10101010_0;
      patterns[27203] = 25'b01101010_01000001_10101011_0;
      patterns[27204] = 25'b01101010_01000010_10101100_0;
      patterns[27205] = 25'b01101010_01000011_10101101_0;
      patterns[27206] = 25'b01101010_01000100_10101110_0;
      patterns[27207] = 25'b01101010_01000101_10101111_0;
      patterns[27208] = 25'b01101010_01000110_10110000_0;
      patterns[27209] = 25'b01101010_01000111_10110001_0;
      patterns[27210] = 25'b01101010_01001000_10110010_0;
      patterns[27211] = 25'b01101010_01001001_10110011_0;
      patterns[27212] = 25'b01101010_01001010_10110100_0;
      patterns[27213] = 25'b01101010_01001011_10110101_0;
      patterns[27214] = 25'b01101010_01001100_10110110_0;
      patterns[27215] = 25'b01101010_01001101_10110111_0;
      patterns[27216] = 25'b01101010_01001110_10111000_0;
      patterns[27217] = 25'b01101010_01001111_10111001_0;
      patterns[27218] = 25'b01101010_01010000_10111010_0;
      patterns[27219] = 25'b01101010_01010001_10111011_0;
      patterns[27220] = 25'b01101010_01010010_10111100_0;
      patterns[27221] = 25'b01101010_01010011_10111101_0;
      patterns[27222] = 25'b01101010_01010100_10111110_0;
      patterns[27223] = 25'b01101010_01010101_10111111_0;
      patterns[27224] = 25'b01101010_01010110_11000000_0;
      patterns[27225] = 25'b01101010_01010111_11000001_0;
      patterns[27226] = 25'b01101010_01011000_11000010_0;
      patterns[27227] = 25'b01101010_01011001_11000011_0;
      patterns[27228] = 25'b01101010_01011010_11000100_0;
      patterns[27229] = 25'b01101010_01011011_11000101_0;
      patterns[27230] = 25'b01101010_01011100_11000110_0;
      patterns[27231] = 25'b01101010_01011101_11000111_0;
      patterns[27232] = 25'b01101010_01011110_11001000_0;
      patterns[27233] = 25'b01101010_01011111_11001001_0;
      patterns[27234] = 25'b01101010_01100000_11001010_0;
      patterns[27235] = 25'b01101010_01100001_11001011_0;
      patterns[27236] = 25'b01101010_01100010_11001100_0;
      patterns[27237] = 25'b01101010_01100011_11001101_0;
      patterns[27238] = 25'b01101010_01100100_11001110_0;
      patterns[27239] = 25'b01101010_01100101_11001111_0;
      patterns[27240] = 25'b01101010_01100110_11010000_0;
      patterns[27241] = 25'b01101010_01100111_11010001_0;
      patterns[27242] = 25'b01101010_01101000_11010010_0;
      patterns[27243] = 25'b01101010_01101001_11010011_0;
      patterns[27244] = 25'b01101010_01101010_11010100_0;
      patterns[27245] = 25'b01101010_01101011_11010101_0;
      patterns[27246] = 25'b01101010_01101100_11010110_0;
      patterns[27247] = 25'b01101010_01101101_11010111_0;
      patterns[27248] = 25'b01101010_01101110_11011000_0;
      patterns[27249] = 25'b01101010_01101111_11011001_0;
      patterns[27250] = 25'b01101010_01110000_11011010_0;
      patterns[27251] = 25'b01101010_01110001_11011011_0;
      patterns[27252] = 25'b01101010_01110010_11011100_0;
      patterns[27253] = 25'b01101010_01110011_11011101_0;
      patterns[27254] = 25'b01101010_01110100_11011110_0;
      patterns[27255] = 25'b01101010_01110101_11011111_0;
      patterns[27256] = 25'b01101010_01110110_11100000_0;
      patterns[27257] = 25'b01101010_01110111_11100001_0;
      patterns[27258] = 25'b01101010_01111000_11100010_0;
      patterns[27259] = 25'b01101010_01111001_11100011_0;
      patterns[27260] = 25'b01101010_01111010_11100100_0;
      patterns[27261] = 25'b01101010_01111011_11100101_0;
      patterns[27262] = 25'b01101010_01111100_11100110_0;
      patterns[27263] = 25'b01101010_01111101_11100111_0;
      patterns[27264] = 25'b01101010_01111110_11101000_0;
      patterns[27265] = 25'b01101010_01111111_11101001_0;
      patterns[27266] = 25'b01101010_10000000_11101010_0;
      patterns[27267] = 25'b01101010_10000001_11101011_0;
      patterns[27268] = 25'b01101010_10000010_11101100_0;
      patterns[27269] = 25'b01101010_10000011_11101101_0;
      patterns[27270] = 25'b01101010_10000100_11101110_0;
      patterns[27271] = 25'b01101010_10000101_11101111_0;
      patterns[27272] = 25'b01101010_10000110_11110000_0;
      patterns[27273] = 25'b01101010_10000111_11110001_0;
      patterns[27274] = 25'b01101010_10001000_11110010_0;
      patterns[27275] = 25'b01101010_10001001_11110011_0;
      patterns[27276] = 25'b01101010_10001010_11110100_0;
      patterns[27277] = 25'b01101010_10001011_11110101_0;
      patterns[27278] = 25'b01101010_10001100_11110110_0;
      patterns[27279] = 25'b01101010_10001101_11110111_0;
      patterns[27280] = 25'b01101010_10001110_11111000_0;
      patterns[27281] = 25'b01101010_10001111_11111001_0;
      patterns[27282] = 25'b01101010_10010000_11111010_0;
      patterns[27283] = 25'b01101010_10010001_11111011_0;
      patterns[27284] = 25'b01101010_10010010_11111100_0;
      patterns[27285] = 25'b01101010_10010011_11111101_0;
      patterns[27286] = 25'b01101010_10010100_11111110_0;
      patterns[27287] = 25'b01101010_10010101_11111111_0;
      patterns[27288] = 25'b01101010_10010110_00000000_1;
      patterns[27289] = 25'b01101010_10010111_00000001_1;
      patterns[27290] = 25'b01101010_10011000_00000010_1;
      patterns[27291] = 25'b01101010_10011001_00000011_1;
      patterns[27292] = 25'b01101010_10011010_00000100_1;
      patterns[27293] = 25'b01101010_10011011_00000101_1;
      patterns[27294] = 25'b01101010_10011100_00000110_1;
      patterns[27295] = 25'b01101010_10011101_00000111_1;
      patterns[27296] = 25'b01101010_10011110_00001000_1;
      patterns[27297] = 25'b01101010_10011111_00001001_1;
      patterns[27298] = 25'b01101010_10100000_00001010_1;
      patterns[27299] = 25'b01101010_10100001_00001011_1;
      patterns[27300] = 25'b01101010_10100010_00001100_1;
      patterns[27301] = 25'b01101010_10100011_00001101_1;
      patterns[27302] = 25'b01101010_10100100_00001110_1;
      patterns[27303] = 25'b01101010_10100101_00001111_1;
      patterns[27304] = 25'b01101010_10100110_00010000_1;
      patterns[27305] = 25'b01101010_10100111_00010001_1;
      patterns[27306] = 25'b01101010_10101000_00010010_1;
      patterns[27307] = 25'b01101010_10101001_00010011_1;
      patterns[27308] = 25'b01101010_10101010_00010100_1;
      patterns[27309] = 25'b01101010_10101011_00010101_1;
      patterns[27310] = 25'b01101010_10101100_00010110_1;
      patterns[27311] = 25'b01101010_10101101_00010111_1;
      patterns[27312] = 25'b01101010_10101110_00011000_1;
      patterns[27313] = 25'b01101010_10101111_00011001_1;
      patterns[27314] = 25'b01101010_10110000_00011010_1;
      patterns[27315] = 25'b01101010_10110001_00011011_1;
      patterns[27316] = 25'b01101010_10110010_00011100_1;
      patterns[27317] = 25'b01101010_10110011_00011101_1;
      patterns[27318] = 25'b01101010_10110100_00011110_1;
      patterns[27319] = 25'b01101010_10110101_00011111_1;
      patterns[27320] = 25'b01101010_10110110_00100000_1;
      patterns[27321] = 25'b01101010_10110111_00100001_1;
      patterns[27322] = 25'b01101010_10111000_00100010_1;
      patterns[27323] = 25'b01101010_10111001_00100011_1;
      patterns[27324] = 25'b01101010_10111010_00100100_1;
      patterns[27325] = 25'b01101010_10111011_00100101_1;
      patterns[27326] = 25'b01101010_10111100_00100110_1;
      patterns[27327] = 25'b01101010_10111101_00100111_1;
      patterns[27328] = 25'b01101010_10111110_00101000_1;
      patterns[27329] = 25'b01101010_10111111_00101001_1;
      patterns[27330] = 25'b01101010_11000000_00101010_1;
      patterns[27331] = 25'b01101010_11000001_00101011_1;
      patterns[27332] = 25'b01101010_11000010_00101100_1;
      patterns[27333] = 25'b01101010_11000011_00101101_1;
      patterns[27334] = 25'b01101010_11000100_00101110_1;
      patterns[27335] = 25'b01101010_11000101_00101111_1;
      patterns[27336] = 25'b01101010_11000110_00110000_1;
      patterns[27337] = 25'b01101010_11000111_00110001_1;
      patterns[27338] = 25'b01101010_11001000_00110010_1;
      patterns[27339] = 25'b01101010_11001001_00110011_1;
      patterns[27340] = 25'b01101010_11001010_00110100_1;
      patterns[27341] = 25'b01101010_11001011_00110101_1;
      patterns[27342] = 25'b01101010_11001100_00110110_1;
      patterns[27343] = 25'b01101010_11001101_00110111_1;
      patterns[27344] = 25'b01101010_11001110_00111000_1;
      patterns[27345] = 25'b01101010_11001111_00111001_1;
      patterns[27346] = 25'b01101010_11010000_00111010_1;
      patterns[27347] = 25'b01101010_11010001_00111011_1;
      patterns[27348] = 25'b01101010_11010010_00111100_1;
      patterns[27349] = 25'b01101010_11010011_00111101_1;
      patterns[27350] = 25'b01101010_11010100_00111110_1;
      patterns[27351] = 25'b01101010_11010101_00111111_1;
      patterns[27352] = 25'b01101010_11010110_01000000_1;
      patterns[27353] = 25'b01101010_11010111_01000001_1;
      patterns[27354] = 25'b01101010_11011000_01000010_1;
      patterns[27355] = 25'b01101010_11011001_01000011_1;
      patterns[27356] = 25'b01101010_11011010_01000100_1;
      patterns[27357] = 25'b01101010_11011011_01000101_1;
      patterns[27358] = 25'b01101010_11011100_01000110_1;
      patterns[27359] = 25'b01101010_11011101_01000111_1;
      patterns[27360] = 25'b01101010_11011110_01001000_1;
      patterns[27361] = 25'b01101010_11011111_01001001_1;
      patterns[27362] = 25'b01101010_11100000_01001010_1;
      patterns[27363] = 25'b01101010_11100001_01001011_1;
      patterns[27364] = 25'b01101010_11100010_01001100_1;
      patterns[27365] = 25'b01101010_11100011_01001101_1;
      patterns[27366] = 25'b01101010_11100100_01001110_1;
      patterns[27367] = 25'b01101010_11100101_01001111_1;
      patterns[27368] = 25'b01101010_11100110_01010000_1;
      patterns[27369] = 25'b01101010_11100111_01010001_1;
      patterns[27370] = 25'b01101010_11101000_01010010_1;
      patterns[27371] = 25'b01101010_11101001_01010011_1;
      patterns[27372] = 25'b01101010_11101010_01010100_1;
      patterns[27373] = 25'b01101010_11101011_01010101_1;
      patterns[27374] = 25'b01101010_11101100_01010110_1;
      patterns[27375] = 25'b01101010_11101101_01010111_1;
      patterns[27376] = 25'b01101010_11101110_01011000_1;
      patterns[27377] = 25'b01101010_11101111_01011001_1;
      patterns[27378] = 25'b01101010_11110000_01011010_1;
      patterns[27379] = 25'b01101010_11110001_01011011_1;
      patterns[27380] = 25'b01101010_11110010_01011100_1;
      patterns[27381] = 25'b01101010_11110011_01011101_1;
      patterns[27382] = 25'b01101010_11110100_01011110_1;
      patterns[27383] = 25'b01101010_11110101_01011111_1;
      patterns[27384] = 25'b01101010_11110110_01100000_1;
      patterns[27385] = 25'b01101010_11110111_01100001_1;
      patterns[27386] = 25'b01101010_11111000_01100010_1;
      patterns[27387] = 25'b01101010_11111001_01100011_1;
      patterns[27388] = 25'b01101010_11111010_01100100_1;
      patterns[27389] = 25'b01101010_11111011_01100101_1;
      patterns[27390] = 25'b01101010_11111100_01100110_1;
      patterns[27391] = 25'b01101010_11111101_01100111_1;
      patterns[27392] = 25'b01101010_11111110_01101000_1;
      patterns[27393] = 25'b01101010_11111111_01101001_1;
      patterns[27394] = 25'b01101011_00000000_01101011_0;
      patterns[27395] = 25'b01101011_00000001_01101100_0;
      patterns[27396] = 25'b01101011_00000010_01101101_0;
      patterns[27397] = 25'b01101011_00000011_01101110_0;
      patterns[27398] = 25'b01101011_00000100_01101111_0;
      patterns[27399] = 25'b01101011_00000101_01110000_0;
      patterns[27400] = 25'b01101011_00000110_01110001_0;
      patterns[27401] = 25'b01101011_00000111_01110010_0;
      patterns[27402] = 25'b01101011_00001000_01110011_0;
      patterns[27403] = 25'b01101011_00001001_01110100_0;
      patterns[27404] = 25'b01101011_00001010_01110101_0;
      patterns[27405] = 25'b01101011_00001011_01110110_0;
      patterns[27406] = 25'b01101011_00001100_01110111_0;
      patterns[27407] = 25'b01101011_00001101_01111000_0;
      patterns[27408] = 25'b01101011_00001110_01111001_0;
      patterns[27409] = 25'b01101011_00001111_01111010_0;
      patterns[27410] = 25'b01101011_00010000_01111011_0;
      patterns[27411] = 25'b01101011_00010001_01111100_0;
      patterns[27412] = 25'b01101011_00010010_01111101_0;
      patterns[27413] = 25'b01101011_00010011_01111110_0;
      patterns[27414] = 25'b01101011_00010100_01111111_0;
      patterns[27415] = 25'b01101011_00010101_10000000_0;
      patterns[27416] = 25'b01101011_00010110_10000001_0;
      patterns[27417] = 25'b01101011_00010111_10000010_0;
      patterns[27418] = 25'b01101011_00011000_10000011_0;
      patterns[27419] = 25'b01101011_00011001_10000100_0;
      patterns[27420] = 25'b01101011_00011010_10000101_0;
      patterns[27421] = 25'b01101011_00011011_10000110_0;
      patterns[27422] = 25'b01101011_00011100_10000111_0;
      patterns[27423] = 25'b01101011_00011101_10001000_0;
      patterns[27424] = 25'b01101011_00011110_10001001_0;
      patterns[27425] = 25'b01101011_00011111_10001010_0;
      patterns[27426] = 25'b01101011_00100000_10001011_0;
      patterns[27427] = 25'b01101011_00100001_10001100_0;
      patterns[27428] = 25'b01101011_00100010_10001101_0;
      patterns[27429] = 25'b01101011_00100011_10001110_0;
      patterns[27430] = 25'b01101011_00100100_10001111_0;
      patterns[27431] = 25'b01101011_00100101_10010000_0;
      patterns[27432] = 25'b01101011_00100110_10010001_0;
      patterns[27433] = 25'b01101011_00100111_10010010_0;
      patterns[27434] = 25'b01101011_00101000_10010011_0;
      patterns[27435] = 25'b01101011_00101001_10010100_0;
      patterns[27436] = 25'b01101011_00101010_10010101_0;
      patterns[27437] = 25'b01101011_00101011_10010110_0;
      patterns[27438] = 25'b01101011_00101100_10010111_0;
      patterns[27439] = 25'b01101011_00101101_10011000_0;
      patterns[27440] = 25'b01101011_00101110_10011001_0;
      patterns[27441] = 25'b01101011_00101111_10011010_0;
      patterns[27442] = 25'b01101011_00110000_10011011_0;
      patterns[27443] = 25'b01101011_00110001_10011100_0;
      patterns[27444] = 25'b01101011_00110010_10011101_0;
      patterns[27445] = 25'b01101011_00110011_10011110_0;
      patterns[27446] = 25'b01101011_00110100_10011111_0;
      patterns[27447] = 25'b01101011_00110101_10100000_0;
      patterns[27448] = 25'b01101011_00110110_10100001_0;
      patterns[27449] = 25'b01101011_00110111_10100010_0;
      patterns[27450] = 25'b01101011_00111000_10100011_0;
      patterns[27451] = 25'b01101011_00111001_10100100_0;
      patterns[27452] = 25'b01101011_00111010_10100101_0;
      patterns[27453] = 25'b01101011_00111011_10100110_0;
      patterns[27454] = 25'b01101011_00111100_10100111_0;
      patterns[27455] = 25'b01101011_00111101_10101000_0;
      patterns[27456] = 25'b01101011_00111110_10101001_0;
      patterns[27457] = 25'b01101011_00111111_10101010_0;
      patterns[27458] = 25'b01101011_01000000_10101011_0;
      patterns[27459] = 25'b01101011_01000001_10101100_0;
      patterns[27460] = 25'b01101011_01000010_10101101_0;
      patterns[27461] = 25'b01101011_01000011_10101110_0;
      patterns[27462] = 25'b01101011_01000100_10101111_0;
      patterns[27463] = 25'b01101011_01000101_10110000_0;
      patterns[27464] = 25'b01101011_01000110_10110001_0;
      patterns[27465] = 25'b01101011_01000111_10110010_0;
      patterns[27466] = 25'b01101011_01001000_10110011_0;
      patterns[27467] = 25'b01101011_01001001_10110100_0;
      patterns[27468] = 25'b01101011_01001010_10110101_0;
      patterns[27469] = 25'b01101011_01001011_10110110_0;
      patterns[27470] = 25'b01101011_01001100_10110111_0;
      patterns[27471] = 25'b01101011_01001101_10111000_0;
      patterns[27472] = 25'b01101011_01001110_10111001_0;
      patterns[27473] = 25'b01101011_01001111_10111010_0;
      patterns[27474] = 25'b01101011_01010000_10111011_0;
      patterns[27475] = 25'b01101011_01010001_10111100_0;
      patterns[27476] = 25'b01101011_01010010_10111101_0;
      patterns[27477] = 25'b01101011_01010011_10111110_0;
      patterns[27478] = 25'b01101011_01010100_10111111_0;
      patterns[27479] = 25'b01101011_01010101_11000000_0;
      patterns[27480] = 25'b01101011_01010110_11000001_0;
      patterns[27481] = 25'b01101011_01010111_11000010_0;
      patterns[27482] = 25'b01101011_01011000_11000011_0;
      patterns[27483] = 25'b01101011_01011001_11000100_0;
      patterns[27484] = 25'b01101011_01011010_11000101_0;
      patterns[27485] = 25'b01101011_01011011_11000110_0;
      patterns[27486] = 25'b01101011_01011100_11000111_0;
      patterns[27487] = 25'b01101011_01011101_11001000_0;
      patterns[27488] = 25'b01101011_01011110_11001001_0;
      patterns[27489] = 25'b01101011_01011111_11001010_0;
      patterns[27490] = 25'b01101011_01100000_11001011_0;
      patterns[27491] = 25'b01101011_01100001_11001100_0;
      patterns[27492] = 25'b01101011_01100010_11001101_0;
      patterns[27493] = 25'b01101011_01100011_11001110_0;
      patterns[27494] = 25'b01101011_01100100_11001111_0;
      patterns[27495] = 25'b01101011_01100101_11010000_0;
      patterns[27496] = 25'b01101011_01100110_11010001_0;
      patterns[27497] = 25'b01101011_01100111_11010010_0;
      patterns[27498] = 25'b01101011_01101000_11010011_0;
      patterns[27499] = 25'b01101011_01101001_11010100_0;
      patterns[27500] = 25'b01101011_01101010_11010101_0;
      patterns[27501] = 25'b01101011_01101011_11010110_0;
      patterns[27502] = 25'b01101011_01101100_11010111_0;
      patterns[27503] = 25'b01101011_01101101_11011000_0;
      patterns[27504] = 25'b01101011_01101110_11011001_0;
      patterns[27505] = 25'b01101011_01101111_11011010_0;
      patterns[27506] = 25'b01101011_01110000_11011011_0;
      patterns[27507] = 25'b01101011_01110001_11011100_0;
      patterns[27508] = 25'b01101011_01110010_11011101_0;
      patterns[27509] = 25'b01101011_01110011_11011110_0;
      patterns[27510] = 25'b01101011_01110100_11011111_0;
      patterns[27511] = 25'b01101011_01110101_11100000_0;
      patterns[27512] = 25'b01101011_01110110_11100001_0;
      patterns[27513] = 25'b01101011_01110111_11100010_0;
      patterns[27514] = 25'b01101011_01111000_11100011_0;
      patterns[27515] = 25'b01101011_01111001_11100100_0;
      patterns[27516] = 25'b01101011_01111010_11100101_0;
      patterns[27517] = 25'b01101011_01111011_11100110_0;
      patterns[27518] = 25'b01101011_01111100_11100111_0;
      patterns[27519] = 25'b01101011_01111101_11101000_0;
      patterns[27520] = 25'b01101011_01111110_11101001_0;
      patterns[27521] = 25'b01101011_01111111_11101010_0;
      patterns[27522] = 25'b01101011_10000000_11101011_0;
      patterns[27523] = 25'b01101011_10000001_11101100_0;
      patterns[27524] = 25'b01101011_10000010_11101101_0;
      patterns[27525] = 25'b01101011_10000011_11101110_0;
      patterns[27526] = 25'b01101011_10000100_11101111_0;
      patterns[27527] = 25'b01101011_10000101_11110000_0;
      patterns[27528] = 25'b01101011_10000110_11110001_0;
      patterns[27529] = 25'b01101011_10000111_11110010_0;
      patterns[27530] = 25'b01101011_10001000_11110011_0;
      patterns[27531] = 25'b01101011_10001001_11110100_0;
      patterns[27532] = 25'b01101011_10001010_11110101_0;
      patterns[27533] = 25'b01101011_10001011_11110110_0;
      patterns[27534] = 25'b01101011_10001100_11110111_0;
      patterns[27535] = 25'b01101011_10001101_11111000_0;
      patterns[27536] = 25'b01101011_10001110_11111001_0;
      patterns[27537] = 25'b01101011_10001111_11111010_0;
      patterns[27538] = 25'b01101011_10010000_11111011_0;
      patterns[27539] = 25'b01101011_10010001_11111100_0;
      patterns[27540] = 25'b01101011_10010010_11111101_0;
      patterns[27541] = 25'b01101011_10010011_11111110_0;
      patterns[27542] = 25'b01101011_10010100_11111111_0;
      patterns[27543] = 25'b01101011_10010101_00000000_1;
      patterns[27544] = 25'b01101011_10010110_00000001_1;
      patterns[27545] = 25'b01101011_10010111_00000010_1;
      patterns[27546] = 25'b01101011_10011000_00000011_1;
      patterns[27547] = 25'b01101011_10011001_00000100_1;
      patterns[27548] = 25'b01101011_10011010_00000101_1;
      patterns[27549] = 25'b01101011_10011011_00000110_1;
      patterns[27550] = 25'b01101011_10011100_00000111_1;
      patterns[27551] = 25'b01101011_10011101_00001000_1;
      patterns[27552] = 25'b01101011_10011110_00001001_1;
      patterns[27553] = 25'b01101011_10011111_00001010_1;
      patterns[27554] = 25'b01101011_10100000_00001011_1;
      patterns[27555] = 25'b01101011_10100001_00001100_1;
      patterns[27556] = 25'b01101011_10100010_00001101_1;
      patterns[27557] = 25'b01101011_10100011_00001110_1;
      patterns[27558] = 25'b01101011_10100100_00001111_1;
      patterns[27559] = 25'b01101011_10100101_00010000_1;
      patterns[27560] = 25'b01101011_10100110_00010001_1;
      patterns[27561] = 25'b01101011_10100111_00010010_1;
      patterns[27562] = 25'b01101011_10101000_00010011_1;
      patterns[27563] = 25'b01101011_10101001_00010100_1;
      patterns[27564] = 25'b01101011_10101010_00010101_1;
      patterns[27565] = 25'b01101011_10101011_00010110_1;
      patterns[27566] = 25'b01101011_10101100_00010111_1;
      patterns[27567] = 25'b01101011_10101101_00011000_1;
      patterns[27568] = 25'b01101011_10101110_00011001_1;
      patterns[27569] = 25'b01101011_10101111_00011010_1;
      patterns[27570] = 25'b01101011_10110000_00011011_1;
      patterns[27571] = 25'b01101011_10110001_00011100_1;
      patterns[27572] = 25'b01101011_10110010_00011101_1;
      patterns[27573] = 25'b01101011_10110011_00011110_1;
      patterns[27574] = 25'b01101011_10110100_00011111_1;
      patterns[27575] = 25'b01101011_10110101_00100000_1;
      patterns[27576] = 25'b01101011_10110110_00100001_1;
      patterns[27577] = 25'b01101011_10110111_00100010_1;
      patterns[27578] = 25'b01101011_10111000_00100011_1;
      patterns[27579] = 25'b01101011_10111001_00100100_1;
      patterns[27580] = 25'b01101011_10111010_00100101_1;
      patterns[27581] = 25'b01101011_10111011_00100110_1;
      patterns[27582] = 25'b01101011_10111100_00100111_1;
      patterns[27583] = 25'b01101011_10111101_00101000_1;
      patterns[27584] = 25'b01101011_10111110_00101001_1;
      patterns[27585] = 25'b01101011_10111111_00101010_1;
      patterns[27586] = 25'b01101011_11000000_00101011_1;
      patterns[27587] = 25'b01101011_11000001_00101100_1;
      patterns[27588] = 25'b01101011_11000010_00101101_1;
      patterns[27589] = 25'b01101011_11000011_00101110_1;
      patterns[27590] = 25'b01101011_11000100_00101111_1;
      patterns[27591] = 25'b01101011_11000101_00110000_1;
      patterns[27592] = 25'b01101011_11000110_00110001_1;
      patterns[27593] = 25'b01101011_11000111_00110010_1;
      patterns[27594] = 25'b01101011_11001000_00110011_1;
      patterns[27595] = 25'b01101011_11001001_00110100_1;
      patterns[27596] = 25'b01101011_11001010_00110101_1;
      patterns[27597] = 25'b01101011_11001011_00110110_1;
      patterns[27598] = 25'b01101011_11001100_00110111_1;
      patterns[27599] = 25'b01101011_11001101_00111000_1;
      patterns[27600] = 25'b01101011_11001110_00111001_1;
      patterns[27601] = 25'b01101011_11001111_00111010_1;
      patterns[27602] = 25'b01101011_11010000_00111011_1;
      patterns[27603] = 25'b01101011_11010001_00111100_1;
      patterns[27604] = 25'b01101011_11010010_00111101_1;
      patterns[27605] = 25'b01101011_11010011_00111110_1;
      patterns[27606] = 25'b01101011_11010100_00111111_1;
      patterns[27607] = 25'b01101011_11010101_01000000_1;
      patterns[27608] = 25'b01101011_11010110_01000001_1;
      patterns[27609] = 25'b01101011_11010111_01000010_1;
      patterns[27610] = 25'b01101011_11011000_01000011_1;
      patterns[27611] = 25'b01101011_11011001_01000100_1;
      patterns[27612] = 25'b01101011_11011010_01000101_1;
      patterns[27613] = 25'b01101011_11011011_01000110_1;
      patterns[27614] = 25'b01101011_11011100_01000111_1;
      patterns[27615] = 25'b01101011_11011101_01001000_1;
      patterns[27616] = 25'b01101011_11011110_01001001_1;
      patterns[27617] = 25'b01101011_11011111_01001010_1;
      patterns[27618] = 25'b01101011_11100000_01001011_1;
      patterns[27619] = 25'b01101011_11100001_01001100_1;
      patterns[27620] = 25'b01101011_11100010_01001101_1;
      patterns[27621] = 25'b01101011_11100011_01001110_1;
      patterns[27622] = 25'b01101011_11100100_01001111_1;
      patterns[27623] = 25'b01101011_11100101_01010000_1;
      patterns[27624] = 25'b01101011_11100110_01010001_1;
      patterns[27625] = 25'b01101011_11100111_01010010_1;
      patterns[27626] = 25'b01101011_11101000_01010011_1;
      patterns[27627] = 25'b01101011_11101001_01010100_1;
      patterns[27628] = 25'b01101011_11101010_01010101_1;
      patterns[27629] = 25'b01101011_11101011_01010110_1;
      patterns[27630] = 25'b01101011_11101100_01010111_1;
      patterns[27631] = 25'b01101011_11101101_01011000_1;
      patterns[27632] = 25'b01101011_11101110_01011001_1;
      patterns[27633] = 25'b01101011_11101111_01011010_1;
      patterns[27634] = 25'b01101011_11110000_01011011_1;
      patterns[27635] = 25'b01101011_11110001_01011100_1;
      patterns[27636] = 25'b01101011_11110010_01011101_1;
      patterns[27637] = 25'b01101011_11110011_01011110_1;
      patterns[27638] = 25'b01101011_11110100_01011111_1;
      patterns[27639] = 25'b01101011_11110101_01100000_1;
      patterns[27640] = 25'b01101011_11110110_01100001_1;
      patterns[27641] = 25'b01101011_11110111_01100010_1;
      patterns[27642] = 25'b01101011_11111000_01100011_1;
      patterns[27643] = 25'b01101011_11111001_01100100_1;
      patterns[27644] = 25'b01101011_11111010_01100101_1;
      patterns[27645] = 25'b01101011_11111011_01100110_1;
      patterns[27646] = 25'b01101011_11111100_01100111_1;
      patterns[27647] = 25'b01101011_11111101_01101000_1;
      patterns[27648] = 25'b01101011_11111110_01101001_1;
      patterns[27649] = 25'b01101011_11111111_01101010_1;
      patterns[27650] = 25'b01101100_00000000_01101100_0;
      patterns[27651] = 25'b01101100_00000001_01101101_0;
      patterns[27652] = 25'b01101100_00000010_01101110_0;
      patterns[27653] = 25'b01101100_00000011_01101111_0;
      patterns[27654] = 25'b01101100_00000100_01110000_0;
      patterns[27655] = 25'b01101100_00000101_01110001_0;
      patterns[27656] = 25'b01101100_00000110_01110010_0;
      patterns[27657] = 25'b01101100_00000111_01110011_0;
      patterns[27658] = 25'b01101100_00001000_01110100_0;
      patterns[27659] = 25'b01101100_00001001_01110101_0;
      patterns[27660] = 25'b01101100_00001010_01110110_0;
      patterns[27661] = 25'b01101100_00001011_01110111_0;
      patterns[27662] = 25'b01101100_00001100_01111000_0;
      patterns[27663] = 25'b01101100_00001101_01111001_0;
      patterns[27664] = 25'b01101100_00001110_01111010_0;
      patterns[27665] = 25'b01101100_00001111_01111011_0;
      patterns[27666] = 25'b01101100_00010000_01111100_0;
      patterns[27667] = 25'b01101100_00010001_01111101_0;
      patterns[27668] = 25'b01101100_00010010_01111110_0;
      patterns[27669] = 25'b01101100_00010011_01111111_0;
      patterns[27670] = 25'b01101100_00010100_10000000_0;
      patterns[27671] = 25'b01101100_00010101_10000001_0;
      patterns[27672] = 25'b01101100_00010110_10000010_0;
      patterns[27673] = 25'b01101100_00010111_10000011_0;
      patterns[27674] = 25'b01101100_00011000_10000100_0;
      patterns[27675] = 25'b01101100_00011001_10000101_0;
      patterns[27676] = 25'b01101100_00011010_10000110_0;
      patterns[27677] = 25'b01101100_00011011_10000111_0;
      patterns[27678] = 25'b01101100_00011100_10001000_0;
      patterns[27679] = 25'b01101100_00011101_10001001_0;
      patterns[27680] = 25'b01101100_00011110_10001010_0;
      patterns[27681] = 25'b01101100_00011111_10001011_0;
      patterns[27682] = 25'b01101100_00100000_10001100_0;
      patterns[27683] = 25'b01101100_00100001_10001101_0;
      patterns[27684] = 25'b01101100_00100010_10001110_0;
      patterns[27685] = 25'b01101100_00100011_10001111_0;
      patterns[27686] = 25'b01101100_00100100_10010000_0;
      patterns[27687] = 25'b01101100_00100101_10010001_0;
      patterns[27688] = 25'b01101100_00100110_10010010_0;
      patterns[27689] = 25'b01101100_00100111_10010011_0;
      patterns[27690] = 25'b01101100_00101000_10010100_0;
      patterns[27691] = 25'b01101100_00101001_10010101_0;
      patterns[27692] = 25'b01101100_00101010_10010110_0;
      patterns[27693] = 25'b01101100_00101011_10010111_0;
      patterns[27694] = 25'b01101100_00101100_10011000_0;
      patterns[27695] = 25'b01101100_00101101_10011001_0;
      patterns[27696] = 25'b01101100_00101110_10011010_0;
      patterns[27697] = 25'b01101100_00101111_10011011_0;
      patterns[27698] = 25'b01101100_00110000_10011100_0;
      patterns[27699] = 25'b01101100_00110001_10011101_0;
      patterns[27700] = 25'b01101100_00110010_10011110_0;
      patterns[27701] = 25'b01101100_00110011_10011111_0;
      patterns[27702] = 25'b01101100_00110100_10100000_0;
      patterns[27703] = 25'b01101100_00110101_10100001_0;
      patterns[27704] = 25'b01101100_00110110_10100010_0;
      patterns[27705] = 25'b01101100_00110111_10100011_0;
      patterns[27706] = 25'b01101100_00111000_10100100_0;
      patterns[27707] = 25'b01101100_00111001_10100101_0;
      patterns[27708] = 25'b01101100_00111010_10100110_0;
      patterns[27709] = 25'b01101100_00111011_10100111_0;
      patterns[27710] = 25'b01101100_00111100_10101000_0;
      patterns[27711] = 25'b01101100_00111101_10101001_0;
      patterns[27712] = 25'b01101100_00111110_10101010_0;
      patterns[27713] = 25'b01101100_00111111_10101011_0;
      patterns[27714] = 25'b01101100_01000000_10101100_0;
      patterns[27715] = 25'b01101100_01000001_10101101_0;
      patterns[27716] = 25'b01101100_01000010_10101110_0;
      patterns[27717] = 25'b01101100_01000011_10101111_0;
      patterns[27718] = 25'b01101100_01000100_10110000_0;
      patterns[27719] = 25'b01101100_01000101_10110001_0;
      patterns[27720] = 25'b01101100_01000110_10110010_0;
      patterns[27721] = 25'b01101100_01000111_10110011_0;
      patterns[27722] = 25'b01101100_01001000_10110100_0;
      patterns[27723] = 25'b01101100_01001001_10110101_0;
      patterns[27724] = 25'b01101100_01001010_10110110_0;
      patterns[27725] = 25'b01101100_01001011_10110111_0;
      patterns[27726] = 25'b01101100_01001100_10111000_0;
      patterns[27727] = 25'b01101100_01001101_10111001_0;
      patterns[27728] = 25'b01101100_01001110_10111010_0;
      patterns[27729] = 25'b01101100_01001111_10111011_0;
      patterns[27730] = 25'b01101100_01010000_10111100_0;
      patterns[27731] = 25'b01101100_01010001_10111101_0;
      patterns[27732] = 25'b01101100_01010010_10111110_0;
      patterns[27733] = 25'b01101100_01010011_10111111_0;
      patterns[27734] = 25'b01101100_01010100_11000000_0;
      patterns[27735] = 25'b01101100_01010101_11000001_0;
      patterns[27736] = 25'b01101100_01010110_11000010_0;
      patterns[27737] = 25'b01101100_01010111_11000011_0;
      patterns[27738] = 25'b01101100_01011000_11000100_0;
      patterns[27739] = 25'b01101100_01011001_11000101_0;
      patterns[27740] = 25'b01101100_01011010_11000110_0;
      patterns[27741] = 25'b01101100_01011011_11000111_0;
      patterns[27742] = 25'b01101100_01011100_11001000_0;
      patterns[27743] = 25'b01101100_01011101_11001001_0;
      patterns[27744] = 25'b01101100_01011110_11001010_0;
      patterns[27745] = 25'b01101100_01011111_11001011_0;
      patterns[27746] = 25'b01101100_01100000_11001100_0;
      patterns[27747] = 25'b01101100_01100001_11001101_0;
      patterns[27748] = 25'b01101100_01100010_11001110_0;
      patterns[27749] = 25'b01101100_01100011_11001111_0;
      patterns[27750] = 25'b01101100_01100100_11010000_0;
      patterns[27751] = 25'b01101100_01100101_11010001_0;
      patterns[27752] = 25'b01101100_01100110_11010010_0;
      patterns[27753] = 25'b01101100_01100111_11010011_0;
      patterns[27754] = 25'b01101100_01101000_11010100_0;
      patterns[27755] = 25'b01101100_01101001_11010101_0;
      patterns[27756] = 25'b01101100_01101010_11010110_0;
      patterns[27757] = 25'b01101100_01101011_11010111_0;
      patterns[27758] = 25'b01101100_01101100_11011000_0;
      patterns[27759] = 25'b01101100_01101101_11011001_0;
      patterns[27760] = 25'b01101100_01101110_11011010_0;
      patterns[27761] = 25'b01101100_01101111_11011011_0;
      patterns[27762] = 25'b01101100_01110000_11011100_0;
      patterns[27763] = 25'b01101100_01110001_11011101_0;
      patterns[27764] = 25'b01101100_01110010_11011110_0;
      patterns[27765] = 25'b01101100_01110011_11011111_0;
      patterns[27766] = 25'b01101100_01110100_11100000_0;
      patterns[27767] = 25'b01101100_01110101_11100001_0;
      patterns[27768] = 25'b01101100_01110110_11100010_0;
      patterns[27769] = 25'b01101100_01110111_11100011_0;
      patterns[27770] = 25'b01101100_01111000_11100100_0;
      patterns[27771] = 25'b01101100_01111001_11100101_0;
      patterns[27772] = 25'b01101100_01111010_11100110_0;
      patterns[27773] = 25'b01101100_01111011_11100111_0;
      patterns[27774] = 25'b01101100_01111100_11101000_0;
      patterns[27775] = 25'b01101100_01111101_11101001_0;
      patterns[27776] = 25'b01101100_01111110_11101010_0;
      patterns[27777] = 25'b01101100_01111111_11101011_0;
      patterns[27778] = 25'b01101100_10000000_11101100_0;
      patterns[27779] = 25'b01101100_10000001_11101101_0;
      patterns[27780] = 25'b01101100_10000010_11101110_0;
      patterns[27781] = 25'b01101100_10000011_11101111_0;
      patterns[27782] = 25'b01101100_10000100_11110000_0;
      patterns[27783] = 25'b01101100_10000101_11110001_0;
      patterns[27784] = 25'b01101100_10000110_11110010_0;
      patterns[27785] = 25'b01101100_10000111_11110011_0;
      patterns[27786] = 25'b01101100_10001000_11110100_0;
      patterns[27787] = 25'b01101100_10001001_11110101_0;
      patterns[27788] = 25'b01101100_10001010_11110110_0;
      patterns[27789] = 25'b01101100_10001011_11110111_0;
      patterns[27790] = 25'b01101100_10001100_11111000_0;
      patterns[27791] = 25'b01101100_10001101_11111001_0;
      patterns[27792] = 25'b01101100_10001110_11111010_0;
      patterns[27793] = 25'b01101100_10001111_11111011_0;
      patterns[27794] = 25'b01101100_10010000_11111100_0;
      patterns[27795] = 25'b01101100_10010001_11111101_0;
      patterns[27796] = 25'b01101100_10010010_11111110_0;
      patterns[27797] = 25'b01101100_10010011_11111111_0;
      patterns[27798] = 25'b01101100_10010100_00000000_1;
      patterns[27799] = 25'b01101100_10010101_00000001_1;
      patterns[27800] = 25'b01101100_10010110_00000010_1;
      patterns[27801] = 25'b01101100_10010111_00000011_1;
      patterns[27802] = 25'b01101100_10011000_00000100_1;
      patterns[27803] = 25'b01101100_10011001_00000101_1;
      patterns[27804] = 25'b01101100_10011010_00000110_1;
      patterns[27805] = 25'b01101100_10011011_00000111_1;
      patterns[27806] = 25'b01101100_10011100_00001000_1;
      patterns[27807] = 25'b01101100_10011101_00001001_1;
      patterns[27808] = 25'b01101100_10011110_00001010_1;
      patterns[27809] = 25'b01101100_10011111_00001011_1;
      patterns[27810] = 25'b01101100_10100000_00001100_1;
      patterns[27811] = 25'b01101100_10100001_00001101_1;
      patterns[27812] = 25'b01101100_10100010_00001110_1;
      patterns[27813] = 25'b01101100_10100011_00001111_1;
      patterns[27814] = 25'b01101100_10100100_00010000_1;
      patterns[27815] = 25'b01101100_10100101_00010001_1;
      patterns[27816] = 25'b01101100_10100110_00010010_1;
      patterns[27817] = 25'b01101100_10100111_00010011_1;
      patterns[27818] = 25'b01101100_10101000_00010100_1;
      patterns[27819] = 25'b01101100_10101001_00010101_1;
      patterns[27820] = 25'b01101100_10101010_00010110_1;
      patterns[27821] = 25'b01101100_10101011_00010111_1;
      patterns[27822] = 25'b01101100_10101100_00011000_1;
      patterns[27823] = 25'b01101100_10101101_00011001_1;
      patterns[27824] = 25'b01101100_10101110_00011010_1;
      patterns[27825] = 25'b01101100_10101111_00011011_1;
      patterns[27826] = 25'b01101100_10110000_00011100_1;
      patterns[27827] = 25'b01101100_10110001_00011101_1;
      patterns[27828] = 25'b01101100_10110010_00011110_1;
      patterns[27829] = 25'b01101100_10110011_00011111_1;
      patterns[27830] = 25'b01101100_10110100_00100000_1;
      patterns[27831] = 25'b01101100_10110101_00100001_1;
      patterns[27832] = 25'b01101100_10110110_00100010_1;
      patterns[27833] = 25'b01101100_10110111_00100011_1;
      patterns[27834] = 25'b01101100_10111000_00100100_1;
      patterns[27835] = 25'b01101100_10111001_00100101_1;
      patterns[27836] = 25'b01101100_10111010_00100110_1;
      patterns[27837] = 25'b01101100_10111011_00100111_1;
      patterns[27838] = 25'b01101100_10111100_00101000_1;
      patterns[27839] = 25'b01101100_10111101_00101001_1;
      patterns[27840] = 25'b01101100_10111110_00101010_1;
      patterns[27841] = 25'b01101100_10111111_00101011_1;
      patterns[27842] = 25'b01101100_11000000_00101100_1;
      patterns[27843] = 25'b01101100_11000001_00101101_1;
      patterns[27844] = 25'b01101100_11000010_00101110_1;
      patterns[27845] = 25'b01101100_11000011_00101111_1;
      patterns[27846] = 25'b01101100_11000100_00110000_1;
      patterns[27847] = 25'b01101100_11000101_00110001_1;
      patterns[27848] = 25'b01101100_11000110_00110010_1;
      patterns[27849] = 25'b01101100_11000111_00110011_1;
      patterns[27850] = 25'b01101100_11001000_00110100_1;
      patterns[27851] = 25'b01101100_11001001_00110101_1;
      patterns[27852] = 25'b01101100_11001010_00110110_1;
      patterns[27853] = 25'b01101100_11001011_00110111_1;
      patterns[27854] = 25'b01101100_11001100_00111000_1;
      patterns[27855] = 25'b01101100_11001101_00111001_1;
      patterns[27856] = 25'b01101100_11001110_00111010_1;
      patterns[27857] = 25'b01101100_11001111_00111011_1;
      patterns[27858] = 25'b01101100_11010000_00111100_1;
      patterns[27859] = 25'b01101100_11010001_00111101_1;
      patterns[27860] = 25'b01101100_11010010_00111110_1;
      patterns[27861] = 25'b01101100_11010011_00111111_1;
      patterns[27862] = 25'b01101100_11010100_01000000_1;
      patterns[27863] = 25'b01101100_11010101_01000001_1;
      patterns[27864] = 25'b01101100_11010110_01000010_1;
      patterns[27865] = 25'b01101100_11010111_01000011_1;
      patterns[27866] = 25'b01101100_11011000_01000100_1;
      patterns[27867] = 25'b01101100_11011001_01000101_1;
      patterns[27868] = 25'b01101100_11011010_01000110_1;
      patterns[27869] = 25'b01101100_11011011_01000111_1;
      patterns[27870] = 25'b01101100_11011100_01001000_1;
      patterns[27871] = 25'b01101100_11011101_01001001_1;
      patterns[27872] = 25'b01101100_11011110_01001010_1;
      patterns[27873] = 25'b01101100_11011111_01001011_1;
      patterns[27874] = 25'b01101100_11100000_01001100_1;
      patterns[27875] = 25'b01101100_11100001_01001101_1;
      patterns[27876] = 25'b01101100_11100010_01001110_1;
      patterns[27877] = 25'b01101100_11100011_01001111_1;
      patterns[27878] = 25'b01101100_11100100_01010000_1;
      patterns[27879] = 25'b01101100_11100101_01010001_1;
      patterns[27880] = 25'b01101100_11100110_01010010_1;
      patterns[27881] = 25'b01101100_11100111_01010011_1;
      patterns[27882] = 25'b01101100_11101000_01010100_1;
      patterns[27883] = 25'b01101100_11101001_01010101_1;
      patterns[27884] = 25'b01101100_11101010_01010110_1;
      patterns[27885] = 25'b01101100_11101011_01010111_1;
      patterns[27886] = 25'b01101100_11101100_01011000_1;
      patterns[27887] = 25'b01101100_11101101_01011001_1;
      patterns[27888] = 25'b01101100_11101110_01011010_1;
      patterns[27889] = 25'b01101100_11101111_01011011_1;
      patterns[27890] = 25'b01101100_11110000_01011100_1;
      patterns[27891] = 25'b01101100_11110001_01011101_1;
      patterns[27892] = 25'b01101100_11110010_01011110_1;
      patterns[27893] = 25'b01101100_11110011_01011111_1;
      patterns[27894] = 25'b01101100_11110100_01100000_1;
      patterns[27895] = 25'b01101100_11110101_01100001_1;
      patterns[27896] = 25'b01101100_11110110_01100010_1;
      patterns[27897] = 25'b01101100_11110111_01100011_1;
      patterns[27898] = 25'b01101100_11111000_01100100_1;
      patterns[27899] = 25'b01101100_11111001_01100101_1;
      patterns[27900] = 25'b01101100_11111010_01100110_1;
      patterns[27901] = 25'b01101100_11111011_01100111_1;
      patterns[27902] = 25'b01101100_11111100_01101000_1;
      patterns[27903] = 25'b01101100_11111101_01101001_1;
      patterns[27904] = 25'b01101100_11111110_01101010_1;
      patterns[27905] = 25'b01101100_11111111_01101011_1;
      patterns[27906] = 25'b01101101_00000000_01101101_0;
      patterns[27907] = 25'b01101101_00000001_01101110_0;
      patterns[27908] = 25'b01101101_00000010_01101111_0;
      patterns[27909] = 25'b01101101_00000011_01110000_0;
      patterns[27910] = 25'b01101101_00000100_01110001_0;
      patterns[27911] = 25'b01101101_00000101_01110010_0;
      patterns[27912] = 25'b01101101_00000110_01110011_0;
      patterns[27913] = 25'b01101101_00000111_01110100_0;
      patterns[27914] = 25'b01101101_00001000_01110101_0;
      patterns[27915] = 25'b01101101_00001001_01110110_0;
      patterns[27916] = 25'b01101101_00001010_01110111_0;
      patterns[27917] = 25'b01101101_00001011_01111000_0;
      patterns[27918] = 25'b01101101_00001100_01111001_0;
      patterns[27919] = 25'b01101101_00001101_01111010_0;
      patterns[27920] = 25'b01101101_00001110_01111011_0;
      patterns[27921] = 25'b01101101_00001111_01111100_0;
      patterns[27922] = 25'b01101101_00010000_01111101_0;
      patterns[27923] = 25'b01101101_00010001_01111110_0;
      patterns[27924] = 25'b01101101_00010010_01111111_0;
      patterns[27925] = 25'b01101101_00010011_10000000_0;
      patterns[27926] = 25'b01101101_00010100_10000001_0;
      patterns[27927] = 25'b01101101_00010101_10000010_0;
      patterns[27928] = 25'b01101101_00010110_10000011_0;
      patterns[27929] = 25'b01101101_00010111_10000100_0;
      patterns[27930] = 25'b01101101_00011000_10000101_0;
      patterns[27931] = 25'b01101101_00011001_10000110_0;
      patterns[27932] = 25'b01101101_00011010_10000111_0;
      patterns[27933] = 25'b01101101_00011011_10001000_0;
      patterns[27934] = 25'b01101101_00011100_10001001_0;
      patterns[27935] = 25'b01101101_00011101_10001010_0;
      patterns[27936] = 25'b01101101_00011110_10001011_0;
      patterns[27937] = 25'b01101101_00011111_10001100_0;
      patterns[27938] = 25'b01101101_00100000_10001101_0;
      patterns[27939] = 25'b01101101_00100001_10001110_0;
      patterns[27940] = 25'b01101101_00100010_10001111_0;
      patterns[27941] = 25'b01101101_00100011_10010000_0;
      patterns[27942] = 25'b01101101_00100100_10010001_0;
      patterns[27943] = 25'b01101101_00100101_10010010_0;
      patterns[27944] = 25'b01101101_00100110_10010011_0;
      patterns[27945] = 25'b01101101_00100111_10010100_0;
      patterns[27946] = 25'b01101101_00101000_10010101_0;
      patterns[27947] = 25'b01101101_00101001_10010110_0;
      patterns[27948] = 25'b01101101_00101010_10010111_0;
      patterns[27949] = 25'b01101101_00101011_10011000_0;
      patterns[27950] = 25'b01101101_00101100_10011001_0;
      patterns[27951] = 25'b01101101_00101101_10011010_0;
      patterns[27952] = 25'b01101101_00101110_10011011_0;
      patterns[27953] = 25'b01101101_00101111_10011100_0;
      patterns[27954] = 25'b01101101_00110000_10011101_0;
      patterns[27955] = 25'b01101101_00110001_10011110_0;
      patterns[27956] = 25'b01101101_00110010_10011111_0;
      patterns[27957] = 25'b01101101_00110011_10100000_0;
      patterns[27958] = 25'b01101101_00110100_10100001_0;
      patterns[27959] = 25'b01101101_00110101_10100010_0;
      patterns[27960] = 25'b01101101_00110110_10100011_0;
      patterns[27961] = 25'b01101101_00110111_10100100_0;
      patterns[27962] = 25'b01101101_00111000_10100101_0;
      patterns[27963] = 25'b01101101_00111001_10100110_0;
      patterns[27964] = 25'b01101101_00111010_10100111_0;
      patterns[27965] = 25'b01101101_00111011_10101000_0;
      patterns[27966] = 25'b01101101_00111100_10101001_0;
      patterns[27967] = 25'b01101101_00111101_10101010_0;
      patterns[27968] = 25'b01101101_00111110_10101011_0;
      patterns[27969] = 25'b01101101_00111111_10101100_0;
      patterns[27970] = 25'b01101101_01000000_10101101_0;
      patterns[27971] = 25'b01101101_01000001_10101110_0;
      patterns[27972] = 25'b01101101_01000010_10101111_0;
      patterns[27973] = 25'b01101101_01000011_10110000_0;
      patterns[27974] = 25'b01101101_01000100_10110001_0;
      patterns[27975] = 25'b01101101_01000101_10110010_0;
      patterns[27976] = 25'b01101101_01000110_10110011_0;
      patterns[27977] = 25'b01101101_01000111_10110100_0;
      patterns[27978] = 25'b01101101_01001000_10110101_0;
      patterns[27979] = 25'b01101101_01001001_10110110_0;
      patterns[27980] = 25'b01101101_01001010_10110111_0;
      patterns[27981] = 25'b01101101_01001011_10111000_0;
      patterns[27982] = 25'b01101101_01001100_10111001_0;
      patterns[27983] = 25'b01101101_01001101_10111010_0;
      patterns[27984] = 25'b01101101_01001110_10111011_0;
      patterns[27985] = 25'b01101101_01001111_10111100_0;
      patterns[27986] = 25'b01101101_01010000_10111101_0;
      patterns[27987] = 25'b01101101_01010001_10111110_0;
      patterns[27988] = 25'b01101101_01010010_10111111_0;
      patterns[27989] = 25'b01101101_01010011_11000000_0;
      patterns[27990] = 25'b01101101_01010100_11000001_0;
      patterns[27991] = 25'b01101101_01010101_11000010_0;
      patterns[27992] = 25'b01101101_01010110_11000011_0;
      patterns[27993] = 25'b01101101_01010111_11000100_0;
      patterns[27994] = 25'b01101101_01011000_11000101_0;
      patterns[27995] = 25'b01101101_01011001_11000110_0;
      patterns[27996] = 25'b01101101_01011010_11000111_0;
      patterns[27997] = 25'b01101101_01011011_11001000_0;
      patterns[27998] = 25'b01101101_01011100_11001001_0;
      patterns[27999] = 25'b01101101_01011101_11001010_0;
      patterns[28000] = 25'b01101101_01011110_11001011_0;
      patterns[28001] = 25'b01101101_01011111_11001100_0;
      patterns[28002] = 25'b01101101_01100000_11001101_0;
      patterns[28003] = 25'b01101101_01100001_11001110_0;
      patterns[28004] = 25'b01101101_01100010_11001111_0;
      patterns[28005] = 25'b01101101_01100011_11010000_0;
      patterns[28006] = 25'b01101101_01100100_11010001_0;
      patterns[28007] = 25'b01101101_01100101_11010010_0;
      patterns[28008] = 25'b01101101_01100110_11010011_0;
      patterns[28009] = 25'b01101101_01100111_11010100_0;
      patterns[28010] = 25'b01101101_01101000_11010101_0;
      patterns[28011] = 25'b01101101_01101001_11010110_0;
      patterns[28012] = 25'b01101101_01101010_11010111_0;
      patterns[28013] = 25'b01101101_01101011_11011000_0;
      patterns[28014] = 25'b01101101_01101100_11011001_0;
      patterns[28015] = 25'b01101101_01101101_11011010_0;
      patterns[28016] = 25'b01101101_01101110_11011011_0;
      patterns[28017] = 25'b01101101_01101111_11011100_0;
      patterns[28018] = 25'b01101101_01110000_11011101_0;
      patterns[28019] = 25'b01101101_01110001_11011110_0;
      patterns[28020] = 25'b01101101_01110010_11011111_0;
      patterns[28021] = 25'b01101101_01110011_11100000_0;
      patterns[28022] = 25'b01101101_01110100_11100001_0;
      patterns[28023] = 25'b01101101_01110101_11100010_0;
      patterns[28024] = 25'b01101101_01110110_11100011_0;
      patterns[28025] = 25'b01101101_01110111_11100100_0;
      patterns[28026] = 25'b01101101_01111000_11100101_0;
      patterns[28027] = 25'b01101101_01111001_11100110_0;
      patterns[28028] = 25'b01101101_01111010_11100111_0;
      patterns[28029] = 25'b01101101_01111011_11101000_0;
      patterns[28030] = 25'b01101101_01111100_11101001_0;
      patterns[28031] = 25'b01101101_01111101_11101010_0;
      patterns[28032] = 25'b01101101_01111110_11101011_0;
      patterns[28033] = 25'b01101101_01111111_11101100_0;
      patterns[28034] = 25'b01101101_10000000_11101101_0;
      patterns[28035] = 25'b01101101_10000001_11101110_0;
      patterns[28036] = 25'b01101101_10000010_11101111_0;
      patterns[28037] = 25'b01101101_10000011_11110000_0;
      patterns[28038] = 25'b01101101_10000100_11110001_0;
      patterns[28039] = 25'b01101101_10000101_11110010_0;
      patterns[28040] = 25'b01101101_10000110_11110011_0;
      patterns[28041] = 25'b01101101_10000111_11110100_0;
      patterns[28042] = 25'b01101101_10001000_11110101_0;
      patterns[28043] = 25'b01101101_10001001_11110110_0;
      patterns[28044] = 25'b01101101_10001010_11110111_0;
      patterns[28045] = 25'b01101101_10001011_11111000_0;
      patterns[28046] = 25'b01101101_10001100_11111001_0;
      patterns[28047] = 25'b01101101_10001101_11111010_0;
      patterns[28048] = 25'b01101101_10001110_11111011_0;
      patterns[28049] = 25'b01101101_10001111_11111100_0;
      patterns[28050] = 25'b01101101_10010000_11111101_0;
      patterns[28051] = 25'b01101101_10010001_11111110_0;
      patterns[28052] = 25'b01101101_10010010_11111111_0;
      patterns[28053] = 25'b01101101_10010011_00000000_1;
      patterns[28054] = 25'b01101101_10010100_00000001_1;
      patterns[28055] = 25'b01101101_10010101_00000010_1;
      patterns[28056] = 25'b01101101_10010110_00000011_1;
      patterns[28057] = 25'b01101101_10010111_00000100_1;
      patterns[28058] = 25'b01101101_10011000_00000101_1;
      patterns[28059] = 25'b01101101_10011001_00000110_1;
      patterns[28060] = 25'b01101101_10011010_00000111_1;
      patterns[28061] = 25'b01101101_10011011_00001000_1;
      patterns[28062] = 25'b01101101_10011100_00001001_1;
      patterns[28063] = 25'b01101101_10011101_00001010_1;
      patterns[28064] = 25'b01101101_10011110_00001011_1;
      patterns[28065] = 25'b01101101_10011111_00001100_1;
      patterns[28066] = 25'b01101101_10100000_00001101_1;
      patterns[28067] = 25'b01101101_10100001_00001110_1;
      patterns[28068] = 25'b01101101_10100010_00001111_1;
      patterns[28069] = 25'b01101101_10100011_00010000_1;
      patterns[28070] = 25'b01101101_10100100_00010001_1;
      patterns[28071] = 25'b01101101_10100101_00010010_1;
      patterns[28072] = 25'b01101101_10100110_00010011_1;
      patterns[28073] = 25'b01101101_10100111_00010100_1;
      patterns[28074] = 25'b01101101_10101000_00010101_1;
      patterns[28075] = 25'b01101101_10101001_00010110_1;
      patterns[28076] = 25'b01101101_10101010_00010111_1;
      patterns[28077] = 25'b01101101_10101011_00011000_1;
      patterns[28078] = 25'b01101101_10101100_00011001_1;
      patterns[28079] = 25'b01101101_10101101_00011010_1;
      patterns[28080] = 25'b01101101_10101110_00011011_1;
      patterns[28081] = 25'b01101101_10101111_00011100_1;
      patterns[28082] = 25'b01101101_10110000_00011101_1;
      patterns[28083] = 25'b01101101_10110001_00011110_1;
      patterns[28084] = 25'b01101101_10110010_00011111_1;
      patterns[28085] = 25'b01101101_10110011_00100000_1;
      patterns[28086] = 25'b01101101_10110100_00100001_1;
      patterns[28087] = 25'b01101101_10110101_00100010_1;
      patterns[28088] = 25'b01101101_10110110_00100011_1;
      patterns[28089] = 25'b01101101_10110111_00100100_1;
      patterns[28090] = 25'b01101101_10111000_00100101_1;
      patterns[28091] = 25'b01101101_10111001_00100110_1;
      patterns[28092] = 25'b01101101_10111010_00100111_1;
      patterns[28093] = 25'b01101101_10111011_00101000_1;
      patterns[28094] = 25'b01101101_10111100_00101001_1;
      patterns[28095] = 25'b01101101_10111101_00101010_1;
      patterns[28096] = 25'b01101101_10111110_00101011_1;
      patterns[28097] = 25'b01101101_10111111_00101100_1;
      patterns[28098] = 25'b01101101_11000000_00101101_1;
      patterns[28099] = 25'b01101101_11000001_00101110_1;
      patterns[28100] = 25'b01101101_11000010_00101111_1;
      patterns[28101] = 25'b01101101_11000011_00110000_1;
      patterns[28102] = 25'b01101101_11000100_00110001_1;
      patterns[28103] = 25'b01101101_11000101_00110010_1;
      patterns[28104] = 25'b01101101_11000110_00110011_1;
      patterns[28105] = 25'b01101101_11000111_00110100_1;
      patterns[28106] = 25'b01101101_11001000_00110101_1;
      patterns[28107] = 25'b01101101_11001001_00110110_1;
      patterns[28108] = 25'b01101101_11001010_00110111_1;
      patterns[28109] = 25'b01101101_11001011_00111000_1;
      patterns[28110] = 25'b01101101_11001100_00111001_1;
      patterns[28111] = 25'b01101101_11001101_00111010_1;
      patterns[28112] = 25'b01101101_11001110_00111011_1;
      patterns[28113] = 25'b01101101_11001111_00111100_1;
      patterns[28114] = 25'b01101101_11010000_00111101_1;
      patterns[28115] = 25'b01101101_11010001_00111110_1;
      patterns[28116] = 25'b01101101_11010010_00111111_1;
      patterns[28117] = 25'b01101101_11010011_01000000_1;
      patterns[28118] = 25'b01101101_11010100_01000001_1;
      patterns[28119] = 25'b01101101_11010101_01000010_1;
      patterns[28120] = 25'b01101101_11010110_01000011_1;
      patterns[28121] = 25'b01101101_11010111_01000100_1;
      patterns[28122] = 25'b01101101_11011000_01000101_1;
      patterns[28123] = 25'b01101101_11011001_01000110_1;
      patterns[28124] = 25'b01101101_11011010_01000111_1;
      patterns[28125] = 25'b01101101_11011011_01001000_1;
      patterns[28126] = 25'b01101101_11011100_01001001_1;
      patterns[28127] = 25'b01101101_11011101_01001010_1;
      patterns[28128] = 25'b01101101_11011110_01001011_1;
      patterns[28129] = 25'b01101101_11011111_01001100_1;
      patterns[28130] = 25'b01101101_11100000_01001101_1;
      patterns[28131] = 25'b01101101_11100001_01001110_1;
      patterns[28132] = 25'b01101101_11100010_01001111_1;
      patterns[28133] = 25'b01101101_11100011_01010000_1;
      patterns[28134] = 25'b01101101_11100100_01010001_1;
      patterns[28135] = 25'b01101101_11100101_01010010_1;
      patterns[28136] = 25'b01101101_11100110_01010011_1;
      patterns[28137] = 25'b01101101_11100111_01010100_1;
      patterns[28138] = 25'b01101101_11101000_01010101_1;
      patterns[28139] = 25'b01101101_11101001_01010110_1;
      patterns[28140] = 25'b01101101_11101010_01010111_1;
      patterns[28141] = 25'b01101101_11101011_01011000_1;
      patterns[28142] = 25'b01101101_11101100_01011001_1;
      patterns[28143] = 25'b01101101_11101101_01011010_1;
      patterns[28144] = 25'b01101101_11101110_01011011_1;
      patterns[28145] = 25'b01101101_11101111_01011100_1;
      patterns[28146] = 25'b01101101_11110000_01011101_1;
      patterns[28147] = 25'b01101101_11110001_01011110_1;
      patterns[28148] = 25'b01101101_11110010_01011111_1;
      patterns[28149] = 25'b01101101_11110011_01100000_1;
      patterns[28150] = 25'b01101101_11110100_01100001_1;
      patterns[28151] = 25'b01101101_11110101_01100010_1;
      patterns[28152] = 25'b01101101_11110110_01100011_1;
      patterns[28153] = 25'b01101101_11110111_01100100_1;
      patterns[28154] = 25'b01101101_11111000_01100101_1;
      patterns[28155] = 25'b01101101_11111001_01100110_1;
      patterns[28156] = 25'b01101101_11111010_01100111_1;
      patterns[28157] = 25'b01101101_11111011_01101000_1;
      patterns[28158] = 25'b01101101_11111100_01101001_1;
      patterns[28159] = 25'b01101101_11111101_01101010_1;
      patterns[28160] = 25'b01101101_11111110_01101011_1;
      patterns[28161] = 25'b01101101_11111111_01101100_1;
      patterns[28162] = 25'b01101110_00000000_01101110_0;
      patterns[28163] = 25'b01101110_00000001_01101111_0;
      patterns[28164] = 25'b01101110_00000010_01110000_0;
      patterns[28165] = 25'b01101110_00000011_01110001_0;
      patterns[28166] = 25'b01101110_00000100_01110010_0;
      patterns[28167] = 25'b01101110_00000101_01110011_0;
      patterns[28168] = 25'b01101110_00000110_01110100_0;
      patterns[28169] = 25'b01101110_00000111_01110101_0;
      patterns[28170] = 25'b01101110_00001000_01110110_0;
      patterns[28171] = 25'b01101110_00001001_01110111_0;
      patterns[28172] = 25'b01101110_00001010_01111000_0;
      patterns[28173] = 25'b01101110_00001011_01111001_0;
      patterns[28174] = 25'b01101110_00001100_01111010_0;
      patterns[28175] = 25'b01101110_00001101_01111011_0;
      patterns[28176] = 25'b01101110_00001110_01111100_0;
      patterns[28177] = 25'b01101110_00001111_01111101_0;
      patterns[28178] = 25'b01101110_00010000_01111110_0;
      patterns[28179] = 25'b01101110_00010001_01111111_0;
      patterns[28180] = 25'b01101110_00010010_10000000_0;
      patterns[28181] = 25'b01101110_00010011_10000001_0;
      patterns[28182] = 25'b01101110_00010100_10000010_0;
      patterns[28183] = 25'b01101110_00010101_10000011_0;
      patterns[28184] = 25'b01101110_00010110_10000100_0;
      patterns[28185] = 25'b01101110_00010111_10000101_0;
      patterns[28186] = 25'b01101110_00011000_10000110_0;
      patterns[28187] = 25'b01101110_00011001_10000111_0;
      patterns[28188] = 25'b01101110_00011010_10001000_0;
      patterns[28189] = 25'b01101110_00011011_10001001_0;
      patterns[28190] = 25'b01101110_00011100_10001010_0;
      patterns[28191] = 25'b01101110_00011101_10001011_0;
      patterns[28192] = 25'b01101110_00011110_10001100_0;
      patterns[28193] = 25'b01101110_00011111_10001101_0;
      patterns[28194] = 25'b01101110_00100000_10001110_0;
      patterns[28195] = 25'b01101110_00100001_10001111_0;
      patterns[28196] = 25'b01101110_00100010_10010000_0;
      patterns[28197] = 25'b01101110_00100011_10010001_0;
      patterns[28198] = 25'b01101110_00100100_10010010_0;
      patterns[28199] = 25'b01101110_00100101_10010011_0;
      patterns[28200] = 25'b01101110_00100110_10010100_0;
      patterns[28201] = 25'b01101110_00100111_10010101_0;
      patterns[28202] = 25'b01101110_00101000_10010110_0;
      patterns[28203] = 25'b01101110_00101001_10010111_0;
      patterns[28204] = 25'b01101110_00101010_10011000_0;
      patterns[28205] = 25'b01101110_00101011_10011001_0;
      patterns[28206] = 25'b01101110_00101100_10011010_0;
      patterns[28207] = 25'b01101110_00101101_10011011_0;
      patterns[28208] = 25'b01101110_00101110_10011100_0;
      patterns[28209] = 25'b01101110_00101111_10011101_0;
      patterns[28210] = 25'b01101110_00110000_10011110_0;
      patterns[28211] = 25'b01101110_00110001_10011111_0;
      patterns[28212] = 25'b01101110_00110010_10100000_0;
      patterns[28213] = 25'b01101110_00110011_10100001_0;
      patterns[28214] = 25'b01101110_00110100_10100010_0;
      patterns[28215] = 25'b01101110_00110101_10100011_0;
      patterns[28216] = 25'b01101110_00110110_10100100_0;
      patterns[28217] = 25'b01101110_00110111_10100101_0;
      patterns[28218] = 25'b01101110_00111000_10100110_0;
      patterns[28219] = 25'b01101110_00111001_10100111_0;
      patterns[28220] = 25'b01101110_00111010_10101000_0;
      patterns[28221] = 25'b01101110_00111011_10101001_0;
      patterns[28222] = 25'b01101110_00111100_10101010_0;
      patterns[28223] = 25'b01101110_00111101_10101011_0;
      patterns[28224] = 25'b01101110_00111110_10101100_0;
      patterns[28225] = 25'b01101110_00111111_10101101_0;
      patterns[28226] = 25'b01101110_01000000_10101110_0;
      patterns[28227] = 25'b01101110_01000001_10101111_0;
      patterns[28228] = 25'b01101110_01000010_10110000_0;
      patterns[28229] = 25'b01101110_01000011_10110001_0;
      patterns[28230] = 25'b01101110_01000100_10110010_0;
      patterns[28231] = 25'b01101110_01000101_10110011_0;
      patterns[28232] = 25'b01101110_01000110_10110100_0;
      patterns[28233] = 25'b01101110_01000111_10110101_0;
      patterns[28234] = 25'b01101110_01001000_10110110_0;
      patterns[28235] = 25'b01101110_01001001_10110111_0;
      patterns[28236] = 25'b01101110_01001010_10111000_0;
      patterns[28237] = 25'b01101110_01001011_10111001_0;
      patterns[28238] = 25'b01101110_01001100_10111010_0;
      patterns[28239] = 25'b01101110_01001101_10111011_0;
      patterns[28240] = 25'b01101110_01001110_10111100_0;
      patterns[28241] = 25'b01101110_01001111_10111101_0;
      patterns[28242] = 25'b01101110_01010000_10111110_0;
      patterns[28243] = 25'b01101110_01010001_10111111_0;
      patterns[28244] = 25'b01101110_01010010_11000000_0;
      patterns[28245] = 25'b01101110_01010011_11000001_0;
      patterns[28246] = 25'b01101110_01010100_11000010_0;
      patterns[28247] = 25'b01101110_01010101_11000011_0;
      patterns[28248] = 25'b01101110_01010110_11000100_0;
      patterns[28249] = 25'b01101110_01010111_11000101_0;
      patterns[28250] = 25'b01101110_01011000_11000110_0;
      patterns[28251] = 25'b01101110_01011001_11000111_0;
      patterns[28252] = 25'b01101110_01011010_11001000_0;
      patterns[28253] = 25'b01101110_01011011_11001001_0;
      patterns[28254] = 25'b01101110_01011100_11001010_0;
      patterns[28255] = 25'b01101110_01011101_11001011_0;
      patterns[28256] = 25'b01101110_01011110_11001100_0;
      patterns[28257] = 25'b01101110_01011111_11001101_0;
      patterns[28258] = 25'b01101110_01100000_11001110_0;
      patterns[28259] = 25'b01101110_01100001_11001111_0;
      patterns[28260] = 25'b01101110_01100010_11010000_0;
      patterns[28261] = 25'b01101110_01100011_11010001_0;
      patterns[28262] = 25'b01101110_01100100_11010010_0;
      patterns[28263] = 25'b01101110_01100101_11010011_0;
      patterns[28264] = 25'b01101110_01100110_11010100_0;
      patterns[28265] = 25'b01101110_01100111_11010101_0;
      patterns[28266] = 25'b01101110_01101000_11010110_0;
      patterns[28267] = 25'b01101110_01101001_11010111_0;
      patterns[28268] = 25'b01101110_01101010_11011000_0;
      patterns[28269] = 25'b01101110_01101011_11011001_0;
      patterns[28270] = 25'b01101110_01101100_11011010_0;
      patterns[28271] = 25'b01101110_01101101_11011011_0;
      patterns[28272] = 25'b01101110_01101110_11011100_0;
      patterns[28273] = 25'b01101110_01101111_11011101_0;
      patterns[28274] = 25'b01101110_01110000_11011110_0;
      patterns[28275] = 25'b01101110_01110001_11011111_0;
      patterns[28276] = 25'b01101110_01110010_11100000_0;
      patterns[28277] = 25'b01101110_01110011_11100001_0;
      patterns[28278] = 25'b01101110_01110100_11100010_0;
      patterns[28279] = 25'b01101110_01110101_11100011_0;
      patterns[28280] = 25'b01101110_01110110_11100100_0;
      patterns[28281] = 25'b01101110_01110111_11100101_0;
      patterns[28282] = 25'b01101110_01111000_11100110_0;
      patterns[28283] = 25'b01101110_01111001_11100111_0;
      patterns[28284] = 25'b01101110_01111010_11101000_0;
      patterns[28285] = 25'b01101110_01111011_11101001_0;
      patterns[28286] = 25'b01101110_01111100_11101010_0;
      patterns[28287] = 25'b01101110_01111101_11101011_0;
      patterns[28288] = 25'b01101110_01111110_11101100_0;
      patterns[28289] = 25'b01101110_01111111_11101101_0;
      patterns[28290] = 25'b01101110_10000000_11101110_0;
      patterns[28291] = 25'b01101110_10000001_11101111_0;
      patterns[28292] = 25'b01101110_10000010_11110000_0;
      patterns[28293] = 25'b01101110_10000011_11110001_0;
      patterns[28294] = 25'b01101110_10000100_11110010_0;
      patterns[28295] = 25'b01101110_10000101_11110011_0;
      patterns[28296] = 25'b01101110_10000110_11110100_0;
      patterns[28297] = 25'b01101110_10000111_11110101_0;
      patterns[28298] = 25'b01101110_10001000_11110110_0;
      patterns[28299] = 25'b01101110_10001001_11110111_0;
      patterns[28300] = 25'b01101110_10001010_11111000_0;
      patterns[28301] = 25'b01101110_10001011_11111001_0;
      patterns[28302] = 25'b01101110_10001100_11111010_0;
      patterns[28303] = 25'b01101110_10001101_11111011_0;
      patterns[28304] = 25'b01101110_10001110_11111100_0;
      patterns[28305] = 25'b01101110_10001111_11111101_0;
      patterns[28306] = 25'b01101110_10010000_11111110_0;
      patterns[28307] = 25'b01101110_10010001_11111111_0;
      patterns[28308] = 25'b01101110_10010010_00000000_1;
      patterns[28309] = 25'b01101110_10010011_00000001_1;
      patterns[28310] = 25'b01101110_10010100_00000010_1;
      patterns[28311] = 25'b01101110_10010101_00000011_1;
      patterns[28312] = 25'b01101110_10010110_00000100_1;
      patterns[28313] = 25'b01101110_10010111_00000101_1;
      patterns[28314] = 25'b01101110_10011000_00000110_1;
      patterns[28315] = 25'b01101110_10011001_00000111_1;
      patterns[28316] = 25'b01101110_10011010_00001000_1;
      patterns[28317] = 25'b01101110_10011011_00001001_1;
      patterns[28318] = 25'b01101110_10011100_00001010_1;
      patterns[28319] = 25'b01101110_10011101_00001011_1;
      patterns[28320] = 25'b01101110_10011110_00001100_1;
      patterns[28321] = 25'b01101110_10011111_00001101_1;
      patterns[28322] = 25'b01101110_10100000_00001110_1;
      patterns[28323] = 25'b01101110_10100001_00001111_1;
      patterns[28324] = 25'b01101110_10100010_00010000_1;
      patterns[28325] = 25'b01101110_10100011_00010001_1;
      patterns[28326] = 25'b01101110_10100100_00010010_1;
      patterns[28327] = 25'b01101110_10100101_00010011_1;
      patterns[28328] = 25'b01101110_10100110_00010100_1;
      patterns[28329] = 25'b01101110_10100111_00010101_1;
      patterns[28330] = 25'b01101110_10101000_00010110_1;
      patterns[28331] = 25'b01101110_10101001_00010111_1;
      patterns[28332] = 25'b01101110_10101010_00011000_1;
      patterns[28333] = 25'b01101110_10101011_00011001_1;
      patterns[28334] = 25'b01101110_10101100_00011010_1;
      patterns[28335] = 25'b01101110_10101101_00011011_1;
      patterns[28336] = 25'b01101110_10101110_00011100_1;
      patterns[28337] = 25'b01101110_10101111_00011101_1;
      patterns[28338] = 25'b01101110_10110000_00011110_1;
      patterns[28339] = 25'b01101110_10110001_00011111_1;
      patterns[28340] = 25'b01101110_10110010_00100000_1;
      patterns[28341] = 25'b01101110_10110011_00100001_1;
      patterns[28342] = 25'b01101110_10110100_00100010_1;
      patterns[28343] = 25'b01101110_10110101_00100011_1;
      patterns[28344] = 25'b01101110_10110110_00100100_1;
      patterns[28345] = 25'b01101110_10110111_00100101_1;
      patterns[28346] = 25'b01101110_10111000_00100110_1;
      patterns[28347] = 25'b01101110_10111001_00100111_1;
      patterns[28348] = 25'b01101110_10111010_00101000_1;
      patterns[28349] = 25'b01101110_10111011_00101001_1;
      patterns[28350] = 25'b01101110_10111100_00101010_1;
      patterns[28351] = 25'b01101110_10111101_00101011_1;
      patterns[28352] = 25'b01101110_10111110_00101100_1;
      patterns[28353] = 25'b01101110_10111111_00101101_1;
      patterns[28354] = 25'b01101110_11000000_00101110_1;
      patterns[28355] = 25'b01101110_11000001_00101111_1;
      patterns[28356] = 25'b01101110_11000010_00110000_1;
      patterns[28357] = 25'b01101110_11000011_00110001_1;
      patterns[28358] = 25'b01101110_11000100_00110010_1;
      patterns[28359] = 25'b01101110_11000101_00110011_1;
      patterns[28360] = 25'b01101110_11000110_00110100_1;
      patterns[28361] = 25'b01101110_11000111_00110101_1;
      patterns[28362] = 25'b01101110_11001000_00110110_1;
      patterns[28363] = 25'b01101110_11001001_00110111_1;
      patterns[28364] = 25'b01101110_11001010_00111000_1;
      patterns[28365] = 25'b01101110_11001011_00111001_1;
      patterns[28366] = 25'b01101110_11001100_00111010_1;
      patterns[28367] = 25'b01101110_11001101_00111011_1;
      patterns[28368] = 25'b01101110_11001110_00111100_1;
      patterns[28369] = 25'b01101110_11001111_00111101_1;
      patterns[28370] = 25'b01101110_11010000_00111110_1;
      patterns[28371] = 25'b01101110_11010001_00111111_1;
      patterns[28372] = 25'b01101110_11010010_01000000_1;
      patterns[28373] = 25'b01101110_11010011_01000001_1;
      patterns[28374] = 25'b01101110_11010100_01000010_1;
      patterns[28375] = 25'b01101110_11010101_01000011_1;
      patterns[28376] = 25'b01101110_11010110_01000100_1;
      patterns[28377] = 25'b01101110_11010111_01000101_1;
      patterns[28378] = 25'b01101110_11011000_01000110_1;
      patterns[28379] = 25'b01101110_11011001_01000111_1;
      patterns[28380] = 25'b01101110_11011010_01001000_1;
      patterns[28381] = 25'b01101110_11011011_01001001_1;
      patterns[28382] = 25'b01101110_11011100_01001010_1;
      patterns[28383] = 25'b01101110_11011101_01001011_1;
      patterns[28384] = 25'b01101110_11011110_01001100_1;
      patterns[28385] = 25'b01101110_11011111_01001101_1;
      patterns[28386] = 25'b01101110_11100000_01001110_1;
      patterns[28387] = 25'b01101110_11100001_01001111_1;
      patterns[28388] = 25'b01101110_11100010_01010000_1;
      patterns[28389] = 25'b01101110_11100011_01010001_1;
      patterns[28390] = 25'b01101110_11100100_01010010_1;
      patterns[28391] = 25'b01101110_11100101_01010011_1;
      patterns[28392] = 25'b01101110_11100110_01010100_1;
      patterns[28393] = 25'b01101110_11100111_01010101_1;
      patterns[28394] = 25'b01101110_11101000_01010110_1;
      patterns[28395] = 25'b01101110_11101001_01010111_1;
      patterns[28396] = 25'b01101110_11101010_01011000_1;
      patterns[28397] = 25'b01101110_11101011_01011001_1;
      patterns[28398] = 25'b01101110_11101100_01011010_1;
      patterns[28399] = 25'b01101110_11101101_01011011_1;
      patterns[28400] = 25'b01101110_11101110_01011100_1;
      patterns[28401] = 25'b01101110_11101111_01011101_1;
      patterns[28402] = 25'b01101110_11110000_01011110_1;
      patterns[28403] = 25'b01101110_11110001_01011111_1;
      patterns[28404] = 25'b01101110_11110010_01100000_1;
      patterns[28405] = 25'b01101110_11110011_01100001_1;
      patterns[28406] = 25'b01101110_11110100_01100010_1;
      patterns[28407] = 25'b01101110_11110101_01100011_1;
      patterns[28408] = 25'b01101110_11110110_01100100_1;
      patterns[28409] = 25'b01101110_11110111_01100101_1;
      patterns[28410] = 25'b01101110_11111000_01100110_1;
      patterns[28411] = 25'b01101110_11111001_01100111_1;
      patterns[28412] = 25'b01101110_11111010_01101000_1;
      patterns[28413] = 25'b01101110_11111011_01101001_1;
      patterns[28414] = 25'b01101110_11111100_01101010_1;
      patterns[28415] = 25'b01101110_11111101_01101011_1;
      patterns[28416] = 25'b01101110_11111110_01101100_1;
      patterns[28417] = 25'b01101110_11111111_01101101_1;
      patterns[28418] = 25'b01101111_00000000_01101111_0;
      patterns[28419] = 25'b01101111_00000001_01110000_0;
      patterns[28420] = 25'b01101111_00000010_01110001_0;
      patterns[28421] = 25'b01101111_00000011_01110010_0;
      patterns[28422] = 25'b01101111_00000100_01110011_0;
      patterns[28423] = 25'b01101111_00000101_01110100_0;
      patterns[28424] = 25'b01101111_00000110_01110101_0;
      patterns[28425] = 25'b01101111_00000111_01110110_0;
      patterns[28426] = 25'b01101111_00001000_01110111_0;
      patterns[28427] = 25'b01101111_00001001_01111000_0;
      patterns[28428] = 25'b01101111_00001010_01111001_0;
      patterns[28429] = 25'b01101111_00001011_01111010_0;
      patterns[28430] = 25'b01101111_00001100_01111011_0;
      patterns[28431] = 25'b01101111_00001101_01111100_0;
      patterns[28432] = 25'b01101111_00001110_01111101_0;
      patterns[28433] = 25'b01101111_00001111_01111110_0;
      patterns[28434] = 25'b01101111_00010000_01111111_0;
      patterns[28435] = 25'b01101111_00010001_10000000_0;
      patterns[28436] = 25'b01101111_00010010_10000001_0;
      patterns[28437] = 25'b01101111_00010011_10000010_0;
      patterns[28438] = 25'b01101111_00010100_10000011_0;
      patterns[28439] = 25'b01101111_00010101_10000100_0;
      patterns[28440] = 25'b01101111_00010110_10000101_0;
      patterns[28441] = 25'b01101111_00010111_10000110_0;
      patterns[28442] = 25'b01101111_00011000_10000111_0;
      patterns[28443] = 25'b01101111_00011001_10001000_0;
      patterns[28444] = 25'b01101111_00011010_10001001_0;
      patterns[28445] = 25'b01101111_00011011_10001010_0;
      patterns[28446] = 25'b01101111_00011100_10001011_0;
      patterns[28447] = 25'b01101111_00011101_10001100_0;
      patterns[28448] = 25'b01101111_00011110_10001101_0;
      patterns[28449] = 25'b01101111_00011111_10001110_0;
      patterns[28450] = 25'b01101111_00100000_10001111_0;
      patterns[28451] = 25'b01101111_00100001_10010000_0;
      patterns[28452] = 25'b01101111_00100010_10010001_0;
      patterns[28453] = 25'b01101111_00100011_10010010_0;
      patterns[28454] = 25'b01101111_00100100_10010011_0;
      patterns[28455] = 25'b01101111_00100101_10010100_0;
      patterns[28456] = 25'b01101111_00100110_10010101_0;
      patterns[28457] = 25'b01101111_00100111_10010110_0;
      patterns[28458] = 25'b01101111_00101000_10010111_0;
      patterns[28459] = 25'b01101111_00101001_10011000_0;
      patterns[28460] = 25'b01101111_00101010_10011001_0;
      patterns[28461] = 25'b01101111_00101011_10011010_0;
      patterns[28462] = 25'b01101111_00101100_10011011_0;
      patterns[28463] = 25'b01101111_00101101_10011100_0;
      patterns[28464] = 25'b01101111_00101110_10011101_0;
      patterns[28465] = 25'b01101111_00101111_10011110_0;
      patterns[28466] = 25'b01101111_00110000_10011111_0;
      patterns[28467] = 25'b01101111_00110001_10100000_0;
      patterns[28468] = 25'b01101111_00110010_10100001_0;
      patterns[28469] = 25'b01101111_00110011_10100010_0;
      patterns[28470] = 25'b01101111_00110100_10100011_0;
      patterns[28471] = 25'b01101111_00110101_10100100_0;
      patterns[28472] = 25'b01101111_00110110_10100101_0;
      patterns[28473] = 25'b01101111_00110111_10100110_0;
      patterns[28474] = 25'b01101111_00111000_10100111_0;
      patterns[28475] = 25'b01101111_00111001_10101000_0;
      patterns[28476] = 25'b01101111_00111010_10101001_0;
      patterns[28477] = 25'b01101111_00111011_10101010_0;
      patterns[28478] = 25'b01101111_00111100_10101011_0;
      patterns[28479] = 25'b01101111_00111101_10101100_0;
      patterns[28480] = 25'b01101111_00111110_10101101_0;
      patterns[28481] = 25'b01101111_00111111_10101110_0;
      patterns[28482] = 25'b01101111_01000000_10101111_0;
      patterns[28483] = 25'b01101111_01000001_10110000_0;
      patterns[28484] = 25'b01101111_01000010_10110001_0;
      patterns[28485] = 25'b01101111_01000011_10110010_0;
      patterns[28486] = 25'b01101111_01000100_10110011_0;
      patterns[28487] = 25'b01101111_01000101_10110100_0;
      patterns[28488] = 25'b01101111_01000110_10110101_0;
      patterns[28489] = 25'b01101111_01000111_10110110_0;
      patterns[28490] = 25'b01101111_01001000_10110111_0;
      patterns[28491] = 25'b01101111_01001001_10111000_0;
      patterns[28492] = 25'b01101111_01001010_10111001_0;
      patterns[28493] = 25'b01101111_01001011_10111010_0;
      patterns[28494] = 25'b01101111_01001100_10111011_0;
      patterns[28495] = 25'b01101111_01001101_10111100_0;
      patterns[28496] = 25'b01101111_01001110_10111101_0;
      patterns[28497] = 25'b01101111_01001111_10111110_0;
      patterns[28498] = 25'b01101111_01010000_10111111_0;
      patterns[28499] = 25'b01101111_01010001_11000000_0;
      patterns[28500] = 25'b01101111_01010010_11000001_0;
      patterns[28501] = 25'b01101111_01010011_11000010_0;
      patterns[28502] = 25'b01101111_01010100_11000011_0;
      patterns[28503] = 25'b01101111_01010101_11000100_0;
      patterns[28504] = 25'b01101111_01010110_11000101_0;
      patterns[28505] = 25'b01101111_01010111_11000110_0;
      patterns[28506] = 25'b01101111_01011000_11000111_0;
      patterns[28507] = 25'b01101111_01011001_11001000_0;
      patterns[28508] = 25'b01101111_01011010_11001001_0;
      patterns[28509] = 25'b01101111_01011011_11001010_0;
      patterns[28510] = 25'b01101111_01011100_11001011_0;
      patterns[28511] = 25'b01101111_01011101_11001100_0;
      patterns[28512] = 25'b01101111_01011110_11001101_0;
      patterns[28513] = 25'b01101111_01011111_11001110_0;
      patterns[28514] = 25'b01101111_01100000_11001111_0;
      patterns[28515] = 25'b01101111_01100001_11010000_0;
      patterns[28516] = 25'b01101111_01100010_11010001_0;
      patterns[28517] = 25'b01101111_01100011_11010010_0;
      patterns[28518] = 25'b01101111_01100100_11010011_0;
      patterns[28519] = 25'b01101111_01100101_11010100_0;
      patterns[28520] = 25'b01101111_01100110_11010101_0;
      patterns[28521] = 25'b01101111_01100111_11010110_0;
      patterns[28522] = 25'b01101111_01101000_11010111_0;
      patterns[28523] = 25'b01101111_01101001_11011000_0;
      patterns[28524] = 25'b01101111_01101010_11011001_0;
      patterns[28525] = 25'b01101111_01101011_11011010_0;
      patterns[28526] = 25'b01101111_01101100_11011011_0;
      patterns[28527] = 25'b01101111_01101101_11011100_0;
      patterns[28528] = 25'b01101111_01101110_11011101_0;
      patterns[28529] = 25'b01101111_01101111_11011110_0;
      patterns[28530] = 25'b01101111_01110000_11011111_0;
      patterns[28531] = 25'b01101111_01110001_11100000_0;
      patterns[28532] = 25'b01101111_01110010_11100001_0;
      patterns[28533] = 25'b01101111_01110011_11100010_0;
      patterns[28534] = 25'b01101111_01110100_11100011_0;
      patterns[28535] = 25'b01101111_01110101_11100100_0;
      patterns[28536] = 25'b01101111_01110110_11100101_0;
      patterns[28537] = 25'b01101111_01110111_11100110_0;
      patterns[28538] = 25'b01101111_01111000_11100111_0;
      patterns[28539] = 25'b01101111_01111001_11101000_0;
      patterns[28540] = 25'b01101111_01111010_11101001_0;
      patterns[28541] = 25'b01101111_01111011_11101010_0;
      patterns[28542] = 25'b01101111_01111100_11101011_0;
      patterns[28543] = 25'b01101111_01111101_11101100_0;
      patterns[28544] = 25'b01101111_01111110_11101101_0;
      patterns[28545] = 25'b01101111_01111111_11101110_0;
      patterns[28546] = 25'b01101111_10000000_11101111_0;
      patterns[28547] = 25'b01101111_10000001_11110000_0;
      patterns[28548] = 25'b01101111_10000010_11110001_0;
      patterns[28549] = 25'b01101111_10000011_11110010_0;
      patterns[28550] = 25'b01101111_10000100_11110011_0;
      patterns[28551] = 25'b01101111_10000101_11110100_0;
      patterns[28552] = 25'b01101111_10000110_11110101_0;
      patterns[28553] = 25'b01101111_10000111_11110110_0;
      patterns[28554] = 25'b01101111_10001000_11110111_0;
      patterns[28555] = 25'b01101111_10001001_11111000_0;
      patterns[28556] = 25'b01101111_10001010_11111001_0;
      patterns[28557] = 25'b01101111_10001011_11111010_0;
      patterns[28558] = 25'b01101111_10001100_11111011_0;
      patterns[28559] = 25'b01101111_10001101_11111100_0;
      patterns[28560] = 25'b01101111_10001110_11111101_0;
      patterns[28561] = 25'b01101111_10001111_11111110_0;
      patterns[28562] = 25'b01101111_10010000_11111111_0;
      patterns[28563] = 25'b01101111_10010001_00000000_1;
      patterns[28564] = 25'b01101111_10010010_00000001_1;
      patterns[28565] = 25'b01101111_10010011_00000010_1;
      patterns[28566] = 25'b01101111_10010100_00000011_1;
      patterns[28567] = 25'b01101111_10010101_00000100_1;
      patterns[28568] = 25'b01101111_10010110_00000101_1;
      patterns[28569] = 25'b01101111_10010111_00000110_1;
      patterns[28570] = 25'b01101111_10011000_00000111_1;
      patterns[28571] = 25'b01101111_10011001_00001000_1;
      patterns[28572] = 25'b01101111_10011010_00001001_1;
      patterns[28573] = 25'b01101111_10011011_00001010_1;
      patterns[28574] = 25'b01101111_10011100_00001011_1;
      patterns[28575] = 25'b01101111_10011101_00001100_1;
      patterns[28576] = 25'b01101111_10011110_00001101_1;
      patterns[28577] = 25'b01101111_10011111_00001110_1;
      patterns[28578] = 25'b01101111_10100000_00001111_1;
      patterns[28579] = 25'b01101111_10100001_00010000_1;
      patterns[28580] = 25'b01101111_10100010_00010001_1;
      patterns[28581] = 25'b01101111_10100011_00010010_1;
      patterns[28582] = 25'b01101111_10100100_00010011_1;
      patterns[28583] = 25'b01101111_10100101_00010100_1;
      patterns[28584] = 25'b01101111_10100110_00010101_1;
      patterns[28585] = 25'b01101111_10100111_00010110_1;
      patterns[28586] = 25'b01101111_10101000_00010111_1;
      patterns[28587] = 25'b01101111_10101001_00011000_1;
      patterns[28588] = 25'b01101111_10101010_00011001_1;
      patterns[28589] = 25'b01101111_10101011_00011010_1;
      patterns[28590] = 25'b01101111_10101100_00011011_1;
      patterns[28591] = 25'b01101111_10101101_00011100_1;
      patterns[28592] = 25'b01101111_10101110_00011101_1;
      patterns[28593] = 25'b01101111_10101111_00011110_1;
      patterns[28594] = 25'b01101111_10110000_00011111_1;
      patterns[28595] = 25'b01101111_10110001_00100000_1;
      patterns[28596] = 25'b01101111_10110010_00100001_1;
      patterns[28597] = 25'b01101111_10110011_00100010_1;
      patterns[28598] = 25'b01101111_10110100_00100011_1;
      patterns[28599] = 25'b01101111_10110101_00100100_1;
      patterns[28600] = 25'b01101111_10110110_00100101_1;
      patterns[28601] = 25'b01101111_10110111_00100110_1;
      patterns[28602] = 25'b01101111_10111000_00100111_1;
      patterns[28603] = 25'b01101111_10111001_00101000_1;
      patterns[28604] = 25'b01101111_10111010_00101001_1;
      patterns[28605] = 25'b01101111_10111011_00101010_1;
      patterns[28606] = 25'b01101111_10111100_00101011_1;
      patterns[28607] = 25'b01101111_10111101_00101100_1;
      patterns[28608] = 25'b01101111_10111110_00101101_1;
      patterns[28609] = 25'b01101111_10111111_00101110_1;
      patterns[28610] = 25'b01101111_11000000_00101111_1;
      patterns[28611] = 25'b01101111_11000001_00110000_1;
      patterns[28612] = 25'b01101111_11000010_00110001_1;
      patterns[28613] = 25'b01101111_11000011_00110010_1;
      patterns[28614] = 25'b01101111_11000100_00110011_1;
      patterns[28615] = 25'b01101111_11000101_00110100_1;
      patterns[28616] = 25'b01101111_11000110_00110101_1;
      patterns[28617] = 25'b01101111_11000111_00110110_1;
      patterns[28618] = 25'b01101111_11001000_00110111_1;
      patterns[28619] = 25'b01101111_11001001_00111000_1;
      patterns[28620] = 25'b01101111_11001010_00111001_1;
      patterns[28621] = 25'b01101111_11001011_00111010_1;
      patterns[28622] = 25'b01101111_11001100_00111011_1;
      patterns[28623] = 25'b01101111_11001101_00111100_1;
      patterns[28624] = 25'b01101111_11001110_00111101_1;
      patterns[28625] = 25'b01101111_11001111_00111110_1;
      patterns[28626] = 25'b01101111_11010000_00111111_1;
      patterns[28627] = 25'b01101111_11010001_01000000_1;
      patterns[28628] = 25'b01101111_11010010_01000001_1;
      patterns[28629] = 25'b01101111_11010011_01000010_1;
      patterns[28630] = 25'b01101111_11010100_01000011_1;
      patterns[28631] = 25'b01101111_11010101_01000100_1;
      patterns[28632] = 25'b01101111_11010110_01000101_1;
      patterns[28633] = 25'b01101111_11010111_01000110_1;
      patterns[28634] = 25'b01101111_11011000_01000111_1;
      patterns[28635] = 25'b01101111_11011001_01001000_1;
      patterns[28636] = 25'b01101111_11011010_01001001_1;
      patterns[28637] = 25'b01101111_11011011_01001010_1;
      patterns[28638] = 25'b01101111_11011100_01001011_1;
      patterns[28639] = 25'b01101111_11011101_01001100_1;
      patterns[28640] = 25'b01101111_11011110_01001101_1;
      patterns[28641] = 25'b01101111_11011111_01001110_1;
      patterns[28642] = 25'b01101111_11100000_01001111_1;
      patterns[28643] = 25'b01101111_11100001_01010000_1;
      patterns[28644] = 25'b01101111_11100010_01010001_1;
      patterns[28645] = 25'b01101111_11100011_01010010_1;
      patterns[28646] = 25'b01101111_11100100_01010011_1;
      patterns[28647] = 25'b01101111_11100101_01010100_1;
      patterns[28648] = 25'b01101111_11100110_01010101_1;
      patterns[28649] = 25'b01101111_11100111_01010110_1;
      patterns[28650] = 25'b01101111_11101000_01010111_1;
      patterns[28651] = 25'b01101111_11101001_01011000_1;
      patterns[28652] = 25'b01101111_11101010_01011001_1;
      patterns[28653] = 25'b01101111_11101011_01011010_1;
      patterns[28654] = 25'b01101111_11101100_01011011_1;
      patterns[28655] = 25'b01101111_11101101_01011100_1;
      patterns[28656] = 25'b01101111_11101110_01011101_1;
      patterns[28657] = 25'b01101111_11101111_01011110_1;
      patterns[28658] = 25'b01101111_11110000_01011111_1;
      patterns[28659] = 25'b01101111_11110001_01100000_1;
      patterns[28660] = 25'b01101111_11110010_01100001_1;
      patterns[28661] = 25'b01101111_11110011_01100010_1;
      patterns[28662] = 25'b01101111_11110100_01100011_1;
      patterns[28663] = 25'b01101111_11110101_01100100_1;
      patterns[28664] = 25'b01101111_11110110_01100101_1;
      patterns[28665] = 25'b01101111_11110111_01100110_1;
      patterns[28666] = 25'b01101111_11111000_01100111_1;
      patterns[28667] = 25'b01101111_11111001_01101000_1;
      patterns[28668] = 25'b01101111_11111010_01101001_1;
      patterns[28669] = 25'b01101111_11111011_01101010_1;
      patterns[28670] = 25'b01101111_11111100_01101011_1;
      patterns[28671] = 25'b01101111_11111101_01101100_1;
      patterns[28672] = 25'b01101111_11111110_01101101_1;
      patterns[28673] = 25'b01101111_11111111_01101110_1;
      patterns[28674] = 25'b01110000_00000000_01110000_0;
      patterns[28675] = 25'b01110000_00000001_01110001_0;
      patterns[28676] = 25'b01110000_00000010_01110010_0;
      patterns[28677] = 25'b01110000_00000011_01110011_0;
      patterns[28678] = 25'b01110000_00000100_01110100_0;
      patterns[28679] = 25'b01110000_00000101_01110101_0;
      patterns[28680] = 25'b01110000_00000110_01110110_0;
      patterns[28681] = 25'b01110000_00000111_01110111_0;
      patterns[28682] = 25'b01110000_00001000_01111000_0;
      patterns[28683] = 25'b01110000_00001001_01111001_0;
      patterns[28684] = 25'b01110000_00001010_01111010_0;
      patterns[28685] = 25'b01110000_00001011_01111011_0;
      patterns[28686] = 25'b01110000_00001100_01111100_0;
      patterns[28687] = 25'b01110000_00001101_01111101_0;
      patterns[28688] = 25'b01110000_00001110_01111110_0;
      patterns[28689] = 25'b01110000_00001111_01111111_0;
      patterns[28690] = 25'b01110000_00010000_10000000_0;
      patterns[28691] = 25'b01110000_00010001_10000001_0;
      patterns[28692] = 25'b01110000_00010010_10000010_0;
      patterns[28693] = 25'b01110000_00010011_10000011_0;
      patterns[28694] = 25'b01110000_00010100_10000100_0;
      patterns[28695] = 25'b01110000_00010101_10000101_0;
      patterns[28696] = 25'b01110000_00010110_10000110_0;
      patterns[28697] = 25'b01110000_00010111_10000111_0;
      patterns[28698] = 25'b01110000_00011000_10001000_0;
      patterns[28699] = 25'b01110000_00011001_10001001_0;
      patterns[28700] = 25'b01110000_00011010_10001010_0;
      patterns[28701] = 25'b01110000_00011011_10001011_0;
      patterns[28702] = 25'b01110000_00011100_10001100_0;
      patterns[28703] = 25'b01110000_00011101_10001101_0;
      patterns[28704] = 25'b01110000_00011110_10001110_0;
      patterns[28705] = 25'b01110000_00011111_10001111_0;
      patterns[28706] = 25'b01110000_00100000_10010000_0;
      patterns[28707] = 25'b01110000_00100001_10010001_0;
      patterns[28708] = 25'b01110000_00100010_10010010_0;
      patterns[28709] = 25'b01110000_00100011_10010011_0;
      patterns[28710] = 25'b01110000_00100100_10010100_0;
      patterns[28711] = 25'b01110000_00100101_10010101_0;
      patterns[28712] = 25'b01110000_00100110_10010110_0;
      patterns[28713] = 25'b01110000_00100111_10010111_0;
      patterns[28714] = 25'b01110000_00101000_10011000_0;
      patterns[28715] = 25'b01110000_00101001_10011001_0;
      patterns[28716] = 25'b01110000_00101010_10011010_0;
      patterns[28717] = 25'b01110000_00101011_10011011_0;
      patterns[28718] = 25'b01110000_00101100_10011100_0;
      patterns[28719] = 25'b01110000_00101101_10011101_0;
      patterns[28720] = 25'b01110000_00101110_10011110_0;
      patterns[28721] = 25'b01110000_00101111_10011111_0;
      patterns[28722] = 25'b01110000_00110000_10100000_0;
      patterns[28723] = 25'b01110000_00110001_10100001_0;
      patterns[28724] = 25'b01110000_00110010_10100010_0;
      patterns[28725] = 25'b01110000_00110011_10100011_0;
      patterns[28726] = 25'b01110000_00110100_10100100_0;
      patterns[28727] = 25'b01110000_00110101_10100101_0;
      patterns[28728] = 25'b01110000_00110110_10100110_0;
      patterns[28729] = 25'b01110000_00110111_10100111_0;
      patterns[28730] = 25'b01110000_00111000_10101000_0;
      patterns[28731] = 25'b01110000_00111001_10101001_0;
      patterns[28732] = 25'b01110000_00111010_10101010_0;
      patterns[28733] = 25'b01110000_00111011_10101011_0;
      patterns[28734] = 25'b01110000_00111100_10101100_0;
      patterns[28735] = 25'b01110000_00111101_10101101_0;
      patterns[28736] = 25'b01110000_00111110_10101110_0;
      patterns[28737] = 25'b01110000_00111111_10101111_0;
      patterns[28738] = 25'b01110000_01000000_10110000_0;
      patterns[28739] = 25'b01110000_01000001_10110001_0;
      patterns[28740] = 25'b01110000_01000010_10110010_0;
      patterns[28741] = 25'b01110000_01000011_10110011_0;
      patterns[28742] = 25'b01110000_01000100_10110100_0;
      patterns[28743] = 25'b01110000_01000101_10110101_0;
      patterns[28744] = 25'b01110000_01000110_10110110_0;
      patterns[28745] = 25'b01110000_01000111_10110111_0;
      patterns[28746] = 25'b01110000_01001000_10111000_0;
      patterns[28747] = 25'b01110000_01001001_10111001_0;
      patterns[28748] = 25'b01110000_01001010_10111010_0;
      patterns[28749] = 25'b01110000_01001011_10111011_0;
      patterns[28750] = 25'b01110000_01001100_10111100_0;
      patterns[28751] = 25'b01110000_01001101_10111101_0;
      patterns[28752] = 25'b01110000_01001110_10111110_0;
      patterns[28753] = 25'b01110000_01001111_10111111_0;
      patterns[28754] = 25'b01110000_01010000_11000000_0;
      patterns[28755] = 25'b01110000_01010001_11000001_0;
      patterns[28756] = 25'b01110000_01010010_11000010_0;
      patterns[28757] = 25'b01110000_01010011_11000011_0;
      patterns[28758] = 25'b01110000_01010100_11000100_0;
      patterns[28759] = 25'b01110000_01010101_11000101_0;
      patterns[28760] = 25'b01110000_01010110_11000110_0;
      patterns[28761] = 25'b01110000_01010111_11000111_0;
      patterns[28762] = 25'b01110000_01011000_11001000_0;
      patterns[28763] = 25'b01110000_01011001_11001001_0;
      patterns[28764] = 25'b01110000_01011010_11001010_0;
      patterns[28765] = 25'b01110000_01011011_11001011_0;
      patterns[28766] = 25'b01110000_01011100_11001100_0;
      patterns[28767] = 25'b01110000_01011101_11001101_0;
      patterns[28768] = 25'b01110000_01011110_11001110_0;
      patterns[28769] = 25'b01110000_01011111_11001111_0;
      patterns[28770] = 25'b01110000_01100000_11010000_0;
      patterns[28771] = 25'b01110000_01100001_11010001_0;
      patterns[28772] = 25'b01110000_01100010_11010010_0;
      patterns[28773] = 25'b01110000_01100011_11010011_0;
      patterns[28774] = 25'b01110000_01100100_11010100_0;
      patterns[28775] = 25'b01110000_01100101_11010101_0;
      patterns[28776] = 25'b01110000_01100110_11010110_0;
      patterns[28777] = 25'b01110000_01100111_11010111_0;
      patterns[28778] = 25'b01110000_01101000_11011000_0;
      patterns[28779] = 25'b01110000_01101001_11011001_0;
      patterns[28780] = 25'b01110000_01101010_11011010_0;
      patterns[28781] = 25'b01110000_01101011_11011011_0;
      patterns[28782] = 25'b01110000_01101100_11011100_0;
      patterns[28783] = 25'b01110000_01101101_11011101_0;
      patterns[28784] = 25'b01110000_01101110_11011110_0;
      patterns[28785] = 25'b01110000_01101111_11011111_0;
      patterns[28786] = 25'b01110000_01110000_11100000_0;
      patterns[28787] = 25'b01110000_01110001_11100001_0;
      patterns[28788] = 25'b01110000_01110010_11100010_0;
      patterns[28789] = 25'b01110000_01110011_11100011_0;
      patterns[28790] = 25'b01110000_01110100_11100100_0;
      patterns[28791] = 25'b01110000_01110101_11100101_0;
      patterns[28792] = 25'b01110000_01110110_11100110_0;
      patterns[28793] = 25'b01110000_01110111_11100111_0;
      patterns[28794] = 25'b01110000_01111000_11101000_0;
      patterns[28795] = 25'b01110000_01111001_11101001_0;
      patterns[28796] = 25'b01110000_01111010_11101010_0;
      patterns[28797] = 25'b01110000_01111011_11101011_0;
      patterns[28798] = 25'b01110000_01111100_11101100_0;
      patterns[28799] = 25'b01110000_01111101_11101101_0;
      patterns[28800] = 25'b01110000_01111110_11101110_0;
      patterns[28801] = 25'b01110000_01111111_11101111_0;
      patterns[28802] = 25'b01110000_10000000_11110000_0;
      patterns[28803] = 25'b01110000_10000001_11110001_0;
      patterns[28804] = 25'b01110000_10000010_11110010_0;
      patterns[28805] = 25'b01110000_10000011_11110011_0;
      patterns[28806] = 25'b01110000_10000100_11110100_0;
      patterns[28807] = 25'b01110000_10000101_11110101_0;
      patterns[28808] = 25'b01110000_10000110_11110110_0;
      patterns[28809] = 25'b01110000_10000111_11110111_0;
      patterns[28810] = 25'b01110000_10001000_11111000_0;
      patterns[28811] = 25'b01110000_10001001_11111001_0;
      patterns[28812] = 25'b01110000_10001010_11111010_0;
      patterns[28813] = 25'b01110000_10001011_11111011_0;
      patterns[28814] = 25'b01110000_10001100_11111100_0;
      patterns[28815] = 25'b01110000_10001101_11111101_0;
      patterns[28816] = 25'b01110000_10001110_11111110_0;
      patterns[28817] = 25'b01110000_10001111_11111111_0;
      patterns[28818] = 25'b01110000_10010000_00000000_1;
      patterns[28819] = 25'b01110000_10010001_00000001_1;
      patterns[28820] = 25'b01110000_10010010_00000010_1;
      patterns[28821] = 25'b01110000_10010011_00000011_1;
      patterns[28822] = 25'b01110000_10010100_00000100_1;
      patterns[28823] = 25'b01110000_10010101_00000101_1;
      patterns[28824] = 25'b01110000_10010110_00000110_1;
      patterns[28825] = 25'b01110000_10010111_00000111_1;
      patterns[28826] = 25'b01110000_10011000_00001000_1;
      patterns[28827] = 25'b01110000_10011001_00001001_1;
      patterns[28828] = 25'b01110000_10011010_00001010_1;
      patterns[28829] = 25'b01110000_10011011_00001011_1;
      patterns[28830] = 25'b01110000_10011100_00001100_1;
      patterns[28831] = 25'b01110000_10011101_00001101_1;
      patterns[28832] = 25'b01110000_10011110_00001110_1;
      patterns[28833] = 25'b01110000_10011111_00001111_1;
      patterns[28834] = 25'b01110000_10100000_00010000_1;
      patterns[28835] = 25'b01110000_10100001_00010001_1;
      patterns[28836] = 25'b01110000_10100010_00010010_1;
      patterns[28837] = 25'b01110000_10100011_00010011_1;
      patterns[28838] = 25'b01110000_10100100_00010100_1;
      patterns[28839] = 25'b01110000_10100101_00010101_1;
      patterns[28840] = 25'b01110000_10100110_00010110_1;
      patterns[28841] = 25'b01110000_10100111_00010111_1;
      patterns[28842] = 25'b01110000_10101000_00011000_1;
      patterns[28843] = 25'b01110000_10101001_00011001_1;
      patterns[28844] = 25'b01110000_10101010_00011010_1;
      patterns[28845] = 25'b01110000_10101011_00011011_1;
      patterns[28846] = 25'b01110000_10101100_00011100_1;
      patterns[28847] = 25'b01110000_10101101_00011101_1;
      patterns[28848] = 25'b01110000_10101110_00011110_1;
      patterns[28849] = 25'b01110000_10101111_00011111_1;
      patterns[28850] = 25'b01110000_10110000_00100000_1;
      patterns[28851] = 25'b01110000_10110001_00100001_1;
      patterns[28852] = 25'b01110000_10110010_00100010_1;
      patterns[28853] = 25'b01110000_10110011_00100011_1;
      patterns[28854] = 25'b01110000_10110100_00100100_1;
      patterns[28855] = 25'b01110000_10110101_00100101_1;
      patterns[28856] = 25'b01110000_10110110_00100110_1;
      patterns[28857] = 25'b01110000_10110111_00100111_1;
      patterns[28858] = 25'b01110000_10111000_00101000_1;
      patterns[28859] = 25'b01110000_10111001_00101001_1;
      patterns[28860] = 25'b01110000_10111010_00101010_1;
      patterns[28861] = 25'b01110000_10111011_00101011_1;
      patterns[28862] = 25'b01110000_10111100_00101100_1;
      patterns[28863] = 25'b01110000_10111101_00101101_1;
      patterns[28864] = 25'b01110000_10111110_00101110_1;
      patterns[28865] = 25'b01110000_10111111_00101111_1;
      patterns[28866] = 25'b01110000_11000000_00110000_1;
      patterns[28867] = 25'b01110000_11000001_00110001_1;
      patterns[28868] = 25'b01110000_11000010_00110010_1;
      patterns[28869] = 25'b01110000_11000011_00110011_1;
      patterns[28870] = 25'b01110000_11000100_00110100_1;
      patterns[28871] = 25'b01110000_11000101_00110101_1;
      patterns[28872] = 25'b01110000_11000110_00110110_1;
      patterns[28873] = 25'b01110000_11000111_00110111_1;
      patterns[28874] = 25'b01110000_11001000_00111000_1;
      patterns[28875] = 25'b01110000_11001001_00111001_1;
      patterns[28876] = 25'b01110000_11001010_00111010_1;
      patterns[28877] = 25'b01110000_11001011_00111011_1;
      patterns[28878] = 25'b01110000_11001100_00111100_1;
      patterns[28879] = 25'b01110000_11001101_00111101_1;
      patterns[28880] = 25'b01110000_11001110_00111110_1;
      patterns[28881] = 25'b01110000_11001111_00111111_1;
      patterns[28882] = 25'b01110000_11010000_01000000_1;
      patterns[28883] = 25'b01110000_11010001_01000001_1;
      patterns[28884] = 25'b01110000_11010010_01000010_1;
      patterns[28885] = 25'b01110000_11010011_01000011_1;
      patterns[28886] = 25'b01110000_11010100_01000100_1;
      patterns[28887] = 25'b01110000_11010101_01000101_1;
      patterns[28888] = 25'b01110000_11010110_01000110_1;
      patterns[28889] = 25'b01110000_11010111_01000111_1;
      patterns[28890] = 25'b01110000_11011000_01001000_1;
      patterns[28891] = 25'b01110000_11011001_01001001_1;
      patterns[28892] = 25'b01110000_11011010_01001010_1;
      patterns[28893] = 25'b01110000_11011011_01001011_1;
      patterns[28894] = 25'b01110000_11011100_01001100_1;
      patterns[28895] = 25'b01110000_11011101_01001101_1;
      patterns[28896] = 25'b01110000_11011110_01001110_1;
      patterns[28897] = 25'b01110000_11011111_01001111_1;
      patterns[28898] = 25'b01110000_11100000_01010000_1;
      patterns[28899] = 25'b01110000_11100001_01010001_1;
      patterns[28900] = 25'b01110000_11100010_01010010_1;
      patterns[28901] = 25'b01110000_11100011_01010011_1;
      patterns[28902] = 25'b01110000_11100100_01010100_1;
      patterns[28903] = 25'b01110000_11100101_01010101_1;
      patterns[28904] = 25'b01110000_11100110_01010110_1;
      patterns[28905] = 25'b01110000_11100111_01010111_1;
      patterns[28906] = 25'b01110000_11101000_01011000_1;
      patterns[28907] = 25'b01110000_11101001_01011001_1;
      patterns[28908] = 25'b01110000_11101010_01011010_1;
      patterns[28909] = 25'b01110000_11101011_01011011_1;
      patterns[28910] = 25'b01110000_11101100_01011100_1;
      patterns[28911] = 25'b01110000_11101101_01011101_1;
      patterns[28912] = 25'b01110000_11101110_01011110_1;
      patterns[28913] = 25'b01110000_11101111_01011111_1;
      patterns[28914] = 25'b01110000_11110000_01100000_1;
      patterns[28915] = 25'b01110000_11110001_01100001_1;
      patterns[28916] = 25'b01110000_11110010_01100010_1;
      patterns[28917] = 25'b01110000_11110011_01100011_1;
      patterns[28918] = 25'b01110000_11110100_01100100_1;
      patterns[28919] = 25'b01110000_11110101_01100101_1;
      patterns[28920] = 25'b01110000_11110110_01100110_1;
      patterns[28921] = 25'b01110000_11110111_01100111_1;
      patterns[28922] = 25'b01110000_11111000_01101000_1;
      patterns[28923] = 25'b01110000_11111001_01101001_1;
      patterns[28924] = 25'b01110000_11111010_01101010_1;
      patterns[28925] = 25'b01110000_11111011_01101011_1;
      patterns[28926] = 25'b01110000_11111100_01101100_1;
      patterns[28927] = 25'b01110000_11111101_01101101_1;
      patterns[28928] = 25'b01110000_11111110_01101110_1;
      patterns[28929] = 25'b01110000_11111111_01101111_1;
      patterns[28930] = 25'b01110001_00000000_01110001_0;
      patterns[28931] = 25'b01110001_00000001_01110010_0;
      patterns[28932] = 25'b01110001_00000010_01110011_0;
      patterns[28933] = 25'b01110001_00000011_01110100_0;
      patterns[28934] = 25'b01110001_00000100_01110101_0;
      patterns[28935] = 25'b01110001_00000101_01110110_0;
      patterns[28936] = 25'b01110001_00000110_01110111_0;
      patterns[28937] = 25'b01110001_00000111_01111000_0;
      patterns[28938] = 25'b01110001_00001000_01111001_0;
      patterns[28939] = 25'b01110001_00001001_01111010_0;
      patterns[28940] = 25'b01110001_00001010_01111011_0;
      patterns[28941] = 25'b01110001_00001011_01111100_0;
      patterns[28942] = 25'b01110001_00001100_01111101_0;
      patterns[28943] = 25'b01110001_00001101_01111110_0;
      patterns[28944] = 25'b01110001_00001110_01111111_0;
      patterns[28945] = 25'b01110001_00001111_10000000_0;
      patterns[28946] = 25'b01110001_00010000_10000001_0;
      patterns[28947] = 25'b01110001_00010001_10000010_0;
      patterns[28948] = 25'b01110001_00010010_10000011_0;
      patterns[28949] = 25'b01110001_00010011_10000100_0;
      patterns[28950] = 25'b01110001_00010100_10000101_0;
      patterns[28951] = 25'b01110001_00010101_10000110_0;
      patterns[28952] = 25'b01110001_00010110_10000111_0;
      patterns[28953] = 25'b01110001_00010111_10001000_0;
      patterns[28954] = 25'b01110001_00011000_10001001_0;
      patterns[28955] = 25'b01110001_00011001_10001010_0;
      patterns[28956] = 25'b01110001_00011010_10001011_0;
      patterns[28957] = 25'b01110001_00011011_10001100_0;
      patterns[28958] = 25'b01110001_00011100_10001101_0;
      patterns[28959] = 25'b01110001_00011101_10001110_0;
      patterns[28960] = 25'b01110001_00011110_10001111_0;
      patterns[28961] = 25'b01110001_00011111_10010000_0;
      patterns[28962] = 25'b01110001_00100000_10010001_0;
      patterns[28963] = 25'b01110001_00100001_10010010_0;
      patterns[28964] = 25'b01110001_00100010_10010011_0;
      patterns[28965] = 25'b01110001_00100011_10010100_0;
      patterns[28966] = 25'b01110001_00100100_10010101_0;
      patterns[28967] = 25'b01110001_00100101_10010110_0;
      patterns[28968] = 25'b01110001_00100110_10010111_0;
      patterns[28969] = 25'b01110001_00100111_10011000_0;
      patterns[28970] = 25'b01110001_00101000_10011001_0;
      patterns[28971] = 25'b01110001_00101001_10011010_0;
      patterns[28972] = 25'b01110001_00101010_10011011_0;
      patterns[28973] = 25'b01110001_00101011_10011100_0;
      patterns[28974] = 25'b01110001_00101100_10011101_0;
      patterns[28975] = 25'b01110001_00101101_10011110_0;
      patterns[28976] = 25'b01110001_00101110_10011111_0;
      patterns[28977] = 25'b01110001_00101111_10100000_0;
      patterns[28978] = 25'b01110001_00110000_10100001_0;
      patterns[28979] = 25'b01110001_00110001_10100010_0;
      patterns[28980] = 25'b01110001_00110010_10100011_0;
      patterns[28981] = 25'b01110001_00110011_10100100_0;
      patterns[28982] = 25'b01110001_00110100_10100101_0;
      patterns[28983] = 25'b01110001_00110101_10100110_0;
      patterns[28984] = 25'b01110001_00110110_10100111_0;
      patterns[28985] = 25'b01110001_00110111_10101000_0;
      patterns[28986] = 25'b01110001_00111000_10101001_0;
      patterns[28987] = 25'b01110001_00111001_10101010_0;
      patterns[28988] = 25'b01110001_00111010_10101011_0;
      patterns[28989] = 25'b01110001_00111011_10101100_0;
      patterns[28990] = 25'b01110001_00111100_10101101_0;
      patterns[28991] = 25'b01110001_00111101_10101110_0;
      patterns[28992] = 25'b01110001_00111110_10101111_0;
      patterns[28993] = 25'b01110001_00111111_10110000_0;
      patterns[28994] = 25'b01110001_01000000_10110001_0;
      patterns[28995] = 25'b01110001_01000001_10110010_0;
      patterns[28996] = 25'b01110001_01000010_10110011_0;
      patterns[28997] = 25'b01110001_01000011_10110100_0;
      patterns[28998] = 25'b01110001_01000100_10110101_0;
      patterns[28999] = 25'b01110001_01000101_10110110_0;
      patterns[29000] = 25'b01110001_01000110_10110111_0;
      patterns[29001] = 25'b01110001_01000111_10111000_0;
      patterns[29002] = 25'b01110001_01001000_10111001_0;
      patterns[29003] = 25'b01110001_01001001_10111010_0;
      patterns[29004] = 25'b01110001_01001010_10111011_0;
      patterns[29005] = 25'b01110001_01001011_10111100_0;
      patterns[29006] = 25'b01110001_01001100_10111101_0;
      patterns[29007] = 25'b01110001_01001101_10111110_0;
      patterns[29008] = 25'b01110001_01001110_10111111_0;
      patterns[29009] = 25'b01110001_01001111_11000000_0;
      patterns[29010] = 25'b01110001_01010000_11000001_0;
      patterns[29011] = 25'b01110001_01010001_11000010_0;
      patterns[29012] = 25'b01110001_01010010_11000011_0;
      patterns[29013] = 25'b01110001_01010011_11000100_0;
      patterns[29014] = 25'b01110001_01010100_11000101_0;
      patterns[29015] = 25'b01110001_01010101_11000110_0;
      patterns[29016] = 25'b01110001_01010110_11000111_0;
      patterns[29017] = 25'b01110001_01010111_11001000_0;
      patterns[29018] = 25'b01110001_01011000_11001001_0;
      patterns[29019] = 25'b01110001_01011001_11001010_0;
      patterns[29020] = 25'b01110001_01011010_11001011_0;
      patterns[29021] = 25'b01110001_01011011_11001100_0;
      patterns[29022] = 25'b01110001_01011100_11001101_0;
      patterns[29023] = 25'b01110001_01011101_11001110_0;
      patterns[29024] = 25'b01110001_01011110_11001111_0;
      patterns[29025] = 25'b01110001_01011111_11010000_0;
      patterns[29026] = 25'b01110001_01100000_11010001_0;
      patterns[29027] = 25'b01110001_01100001_11010010_0;
      patterns[29028] = 25'b01110001_01100010_11010011_0;
      patterns[29029] = 25'b01110001_01100011_11010100_0;
      patterns[29030] = 25'b01110001_01100100_11010101_0;
      patterns[29031] = 25'b01110001_01100101_11010110_0;
      patterns[29032] = 25'b01110001_01100110_11010111_0;
      patterns[29033] = 25'b01110001_01100111_11011000_0;
      patterns[29034] = 25'b01110001_01101000_11011001_0;
      patterns[29035] = 25'b01110001_01101001_11011010_0;
      patterns[29036] = 25'b01110001_01101010_11011011_0;
      patterns[29037] = 25'b01110001_01101011_11011100_0;
      patterns[29038] = 25'b01110001_01101100_11011101_0;
      patterns[29039] = 25'b01110001_01101101_11011110_0;
      patterns[29040] = 25'b01110001_01101110_11011111_0;
      patterns[29041] = 25'b01110001_01101111_11100000_0;
      patterns[29042] = 25'b01110001_01110000_11100001_0;
      patterns[29043] = 25'b01110001_01110001_11100010_0;
      patterns[29044] = 25'b01110001_01110010_11100011_0;
      patterns[29045] = 25'b01110001_01110011_11100100_0;
      patterns[29046] = 25'b01110001_01110100_11100101_0;
      patterns[29047] = 25'b01110001_01110101_11100110_0;
      patterns[29048] = 25'b01110001_01110110_11100111_0;
      patterns[29049] = 25'b01110001_01110111_11101000_0;
      patterns[29050] = 25'b01110001_01111000_11101001_0;
      patterns[29051] = 25'b01110001_01111001_11101010_0;
      patterns[29052] = 25'b01110001_01111010_11101011_0;
      patterns[29053] = 25'b01110001_01111011_11101100_0;
      patterns[29054] = 25'b01110001_01111100_11101101_0;
      patterns[29055] = 25'b01110001_01111101_11101110_0;
      patterns[29056] = 25'b01110001_01111110_11101111_0;
      patterns[29057] = 25'b01110001_01111111_11110000_0;
      patterns[29058] = 25'b01110001_10000000_11110001_0;
      patterns[29059] = 25'b01110001_10000001_11110010_0;
      patterns[29060] = 25'b01110001_10000010_11110011_0;
      patterns[29061] = 25'b01110001_10000011_11110100_0;
      patterns[29062] = 25'b01110001_10000100_11110101_0;
      patterns[29063] = 25'b01110001_10000101_11110110_0;
      patterns[29064] = 25'b01110001_10000110_11110111_0;
      patterns[29065] = 25'b01110001_10000111_11111000_0;
      patterns[29066] = 25'b01110001_10001000_11111001_0;
      patterns[29067] = 25'b01110001_10001001_11111010_0;
      patterns[29068] = 25'b01110001_10001010_11111011_0;
      patterns[29069] = 25'b01110001_10001011_11111100_0;
      patterns[29070] = 25'b01110001_10001100_11111101_0;
      patterns[29071] = 25'b01110001_10001101_11111110_0;
      patterns[29072] = 25'b01110001_10001110_11111111_0;
      patterns[29073] = 25'b01110001_10001111_00000000_1;
      patterns[29074] = 25'b01110001_10010000_00000001_1;
      patterns[29075] = 25'b01110001_10010001_00000010_1;
      patterns[29076] = 25'b01110001_10010010_00000011_1;
      patterns[29077] = 25'b01110001_10010011_00000100_1;
      patterns[29078] = 25'b01110001_10010100_00000101_1;
      patterns[29079] = 25'b01110001_10010101_00000110_1;
      patterns[29080] = 25'b01110001_10010110_00000111_1;
      patterns[29081] = 25'b01110001_10010111_00001000_1;
      patterns[29082] = 25'b01110001_10011000_00001001_1;
      patterns[29083] = 25'b01110001_10011001_00001010_1;
      patterns[29084] = 25'b01110001_10011010_00001011_1;
      patterns[29085] = 25'b01110001_10011011_00001100_1;
      patterns[29086] = 25'b01110001_10011100_00001101_1;
      patterns[29087] = 25'b01110001_10011101_00001110_1;
      patterns[29088] = 25'b01110001_10011110_00001111_1;
      patterns[29089] = 25'b01110001_10011111_00010000_1;
      patterns[29090] = 25'b01110001_10100000_00010001_1;
      patterns[29091] = 25'b01110001_10100001_00010010_1;
      patterns[29092] = 25'b01110001_10100010_00010011_1;
      patterns[29093] = 25'b01110001_10100011_00010100_1;
      patterns[29094] = 25'b01110001_10100100_00010101_1;
      patterns[29095] = 25'b01110001_10100101_00010110_1;
      patterns[29096] = 25'b01110001_10100110_00010111_1;
      patterns[29097] = 25'b01110001_10100111_00011000_1;
      patterns[29098] = 25'b01110001_10101000_00011001_1;
      patterns[29099] = 25'b01110001_10101001_00011010_1;
      patterns[29100] = 25'b01110001_10101010_00011011_1;
      patterns[29101] = 25'b01110001_10101011_00011100_1;
      patterns[29102] = 25'b01110001_10101100_00011101_1;
      patterns[29103] = 25'b01110001_10101101_00011110_1;
      patterns[29104] = 25'b01110001_10101110_00011111_1;
      patterns[29105] = 25'b01110001_10101111_00100000_1;
      patterns[29106] = 25'b01110001_10110000_00100001_1;
      patterns[29107] = 25'b01110001_10110001_00100010_1;
      patterns[29108] = 25'b01110001_10110010_00100011_1;
      patterns[29109] = 25'b01110001_10110011_00100100_1;
      patterns[29110] = 25'b01110001_10110100_00100101_1;
      patterns[29111] = 25'b01110001_10110101_00100110_1;
      patterns[29112] = 25'b01110001_10110110_00100111_1;
      patterns[29113] = 25'b01110001_10110111_00101000_1;
      patterns[29114] = 25'b01110001_10111000_00101001_1;
      patterns[29115] = 25'b01110001_10111001_00101010_1;
      patterns[29116] = 25'b01110001_10111010_00101011_1;
      patterns[29117] = 25'b01110001_10111011_00101100_1;
      patterns[29118] = 25'b01110001_10111100_00101101_1;
      patterns[29119] = 25'b01110001_10111101_00101110_1;
      patterns[29120] = 25'b01110001_10111110_00101111_1;
      patterns[29121] = 25'b01110001_10111111_00110000_1;
      patterns[29122] = 25'b01110001_11000000_00110001_1;
      patterns[29123] = 25'b01110001_11000001_00110010_1;
      patterns[29124] = 25'b01110001_11000010_00110011_1;
      patterns[29125] = 25'b01110001_11000011_00110100_1;
      patterns[29126] = 25'b01110001_11000100_00110101_1;
      patterns[29127] = 25'b01110001_11000101_00110110_1;
      patterns[29128] = 25'b01110001_11000110_00110111_1;
      patterns[29129] = 25'b01110001_11000111_00111000_1;
      patterns[29130] = 25'b01110001_11001000_00111001_1;
      patterns[29131] = 25'b01110001_11001001_00111010_1;
      patterns[29132] = 25'b01110001_11001010_00111011_1;
      patterns[29133] = 25'b01110001_11001011_00111100_1;
      patterns[29134] = 25'b01110001_11001100_00111101_1;
      patterns[29135] = 25'b01110001_11001101_00111110_1;
      patterns[29136] = 25'b01110001_11001110_00111111_1;
      patterns[29137] = 25'b01110001_11001111_01000000_1;
      patterns[29138] = 25'b01110001_11010000_01000001_1;
      patterns[29139] = 25'b01110001_11010001_01000010_1;
      patterns[29140] = 25'b01110001_11010010_01000011_1;
      patterns[29141] = 25'b01110001_11010011_01000100_1;
      patterns[29142] = 25'b01110001_11010100_01000101_1;
      patterns[29143] = 25'b01110001_11010101_01000110_1;
      patterns[29144] = 25'b01110001_11010110_01000111_1;
      patterns[29145] = 25'b01110001_11010111_01001000_1;
      patterns[29146] = 25'b01110001_11011000_01001001_1;
      patterns[29147] = 25'b01110001_11011001_01001010_1;
      patterns[29148] = 25'b01110001_11011010_01001011_1;
      patterns[29149] = 25'b01110001_11011011_01001100_1;
      patterns[29150] = 25'b01110001_11011100_01001101_1;
      patterns[29151] = 25'b01110001_11011101_01001110_1;
      patterns[29152] = 25'b01110001_11011110_01001111_1;
      patterns[29153] = 25'b01110001_11011111_01010000_1;
      patterns[29154] = 25'b01110001_11100000_01010001_1;
      patterns[29155] = 25'b01110001_11100001_01010010_1;
      patterns[29156] = 25'b01110001_11100010_01010011_1;
      patterns[29157] = 25'b01110001_11100011_01010100_1;
      patterns[29158] = 25'b01110001_11100100_01010101_1;
      patterns[29159] = 25'b01110001_11100101_01010110_1;
      patterns[29160] = 25'b01110001_11100110_01010111_1;
      patterns[29161] = 25'b01110001_11100111_01011000_1;
      patterns[29162] = 25'b01110001_11101000_01011001_1;
      patterns[29163] = 25'b01110001_11101001_01011010_1;
      patterns[29164] = 25'b01110001_11101010_01011011_1;
      patterns[29165] = 25'b01110001_11101011_01011100_1;
      patterns[29166] = 25'b01110001_11101100_01011101_1;
      patterns[29167] = 25'b01110001_11101101_01011110_1;
      patterns[29168] = 25'b01110001_11101110_01011111_1;
      patterns[29169] = 25'b01110001_11101111_01100000_1;
      patterns[29170] = 25'b01110001_11110000_01100001_1;
      patterns[29171] = 25'b01110001_11110001_01100010_1;
      patterns[29172] = 25'b01110001_11110010_01100011_1;
      patterns[29173] = 25'b01110001_11110011_01100100_1;
      patterns[29174] = 25'b01110001_11110100_01100101_1;
      patterns[29175] = 25'b01110001_11110101_01100110_1;
      patterns[29176] = 25'b01110001_11110110_01100111_1;
      patterns[29177] = 25'b01110001_11110111_01101000_1;
      patterns[29178] = 25'b01110001_11111000_01101001_1;
      patterns[29179] = 25'b01110001_11111001_01101010_1;
      patterns[29180] = 25'b01110001_11111010_01101011_1;
      patterns[29181] = 25'b01110001_11111011_01101100_1;
      patterns[29182] = 25'b01110001_11111100_01101101_1;
      patterns[29183] = 25'b01110001_11111101_01101110_1;
      patterns[29184] = 25'b01110001_11111110_01101111_1;
      patterns[29185] = 25'b01110001_11111111_01110000_1;
      patterns[29186] = 25'b01110010_00000000_01110010_0;
      patterns[29187] = 25'b01110010_00000001_01110011_0;
      patterns[29188] = 25'b01110010_00000010_01110100_0;
      patterns[29189] = 25'b01110010_00000011_01110101_0;
      patterns[29190] = 25'b01110010_00000100_01110110_0;
      patterns[29191] = 25'b01110010_00000101_01110111_0;
      patterns[29192] = 25'b01110010_00000110_01111000_0;
      patterns[29193] = 25'b01110010_00000111_01111001_0;
      patterns[29194] = 25'b01110010_00001000_01111010_0;
      patterns[29195] = 25'b01110010_00001001_01111011_0;
      patterns[29196] = 25'b01110010_00001010_01111100_0;
      patterns[29197] = 25'b01110010_00001011_01111101_0;
      patterns[29198] = 25'b01110010_00001100_01111110_0;
      patterns[29199] = 25'b01110010_00001101_01111111_0;
      patterns[29200] = 25'b01110010_00001110_10000000_0;
      patterns[29201] = 25'b01110010_00001111_10000001_0;
      patterns[29202] = 25'b01110010_00010000_10000010_0;
      patterns[29203] = 25'b01110010_00010001_10000011_0;
      patterns[29204] = 25'b01110010_00010010_10000100_0;
      patterns[29205] = 25'b01110010_00010011_10000101_0;
      patterns[29206] = 25'b01110010_00010100_10000110_0;
      patterns[29207] = 25'b01110010_00010101_10000111_0;
      patterns[29208] = 25'b01110010_00010110_10001000_0;
      patterns[29209] = 25'b01110010_00010111_10001001_0;
      patterns[29210] = 25'b01110010_00011000_10001010_0;
      patterns[29211] = 25'b01110010_00011001_10001011_0;
      patterns[29212] = 25'b01110010_00011010_10001100_0;
      patterns[29213] = 25'b01110010_00011011_10001101_0;
      patterns[29214] = 25'b01110010_00011100_10001110_0;
      patterns[29215] = 25'b01110010_00011101_10001111_0;
      patterns[29216] = 25'b01110010_00011110_10010000_0;
      patterns[29217] = 25'b01110010_00011111_10010001_0;
      patterns[29218] = 25'b01110010_00100000_10010010_0;
      patterns[29219] = 25'b01110010_00100001_10010011_0;
      patterns[29220] = 25'b01110010_00100010_10010100_0;
      patterns[29221] = 25'b01110010_00100011_10010101_0;
      patterns[29222] = 25'b01110010_00100100_10010110_0;
      patterns[29223] = 25'b01110010_00100101_10010111_0;
      patterns[29224] = 25'b01110010_00100110_10011000_0;
      patterns[29225] = 25'b01110010_00100111_10011001_0;
      patterns[29226] = 25'b01110010_00101000_10011010_0;
      patterns[29227] = 25'b01110010_00101001_10011011_0;
      patterns[29228] = 25'b01110010_00101010_10011100_0;
      patterns[29229] = 25'b01110010_00101011_10011101_0;
      patterns[29230] = 25'b01110010_00101100_10011110_0;
      patterns[29231] = 25'b01110010_00101101_10011111_0;
      patterns[29232] = 25'b01110010_00101110_10100000_0;
      patterns[29233] = 25'b01110010_00101111_10100001_0;
      patterns[29234] = 25'b01110010_00110000_10100010_0;
      patterns[29235] = 25'b01110010_00110001_10100011_0;
      patterns[29236] = 25'b01110010_00110010_10100100_0;
      patterns[29237] = 25'b01110010_00110011_10100101_0;
      patterns[29238] = 25'b01110010_00110100_10100110_0;
      patterns[29239] = 25'b01110010_00110101_10100111_0;
      patterns[29240] = 25'b01110010_00110110_10101000_0;
      patterns[29241] = 25'b01110010_00110111_10101001_0;
      patterns[29242] = 25'b01110010_00111000_10101010_0;
      patterns[29243] = 25'b01110010_00111001_10101011_0;
      patterns[29244] = 25'b01110010_00111010_10101100_0;
      patterns[29245] = 25'b01110010_00111011_10101101_0;
      patterns[29246] = 25'b01110010_00111100_10101110_0;
      patterns[29247] = 25'b01110010_00111101_10101111_0;
      patterns[29248] = 25'b01110010_00111110_10110000_0;
      patterns[29249] = 25'b01110010_00111111_10110001_0;
      patterns[29250] = 25'b01110010_01000000_10110010_0;
      patterns[29251] = 25'b01110010_01000001_10110011_0;
      patterns[29252] = 25'b01110010_01000010_10110100_0;
      patterns[29253] = 25'b01110010_01000011_10110101_0;
      patterns[29254] = 25'b01110010_01000100_10110110_0;
      patterns[29255] = 25'b01110010_01000101_10110111_0;
      patterns[29256] = 25'b01110010_01000110_10111000_0;
      patterns[29257] = 25'b01110010_01000111_10111001_0;
      patterns[29258] = 25'b01110010_01001000_10111010_0;
      patterns[29259] = 25'b01110010_01001001_10111011_0;
      patterns[29260] = 25'b01110010_01001010_10111100_0;
      patterns[29261] = 25'b01110010_01001011_10111101_0;
      patterns[29262] = 25'b01110010_01001100_10111110_0;
      patterns[29263] = 25'b01110010_01001101_10111111_0;
      patterns[29264] = 25'b01110010_01001110_11000000_0;
      patterns[29265] = 25'b01110010_01001111_11000001_0;
      patterns[29266] = 25'b01110010_01010000_11000010_0;
      patterns[29267] = 25'b01110010_01010001_11000011_0;
      patterns[29268] = 25'b01110010_01010010_11000100_0;
      patterns[29269] = 25'b01110010_01010011_11000101_0;
      patterns[29270] = 25'b01110010_01010100_11000110_0;
      patterns[29271] = 25'b01110010_01010101_11000111_0;
      patterns[29272] = 25'b01110010_01010110_11001000_0;
      patterns[29273] = 25'b01110010_01010111_11001001_0;
      patterns[29274] = 25'b01110010_01011000_11001010_0;
      patterns[29275] = 25'b01110010_01011001_11001011_0;
      patterns[29276] = 25'b01110010_01011010_11001100_0;
      patterns[29277] = 25'b01110010_01011011_11001101_0;
      patterns[29278] = 25'b01110010_01011100_11001110_0;
      patterns[29279] = 25'b01110010_01011101_11001111_0;
      patterns[29280] = 25'b01110010_01011110_11010000_0;
      patterns[29281] = 25'b01110010_01011111_11010001_0;
      patterns[29282] = 25'b01110010_01100000_11010010_0;
      patterns[29283] = 25'b01110010_01100001_11010011_0;
      patterns[29284] = 25'b01110010_01100010_11010100_0;
      patterns[29285] = 25'b01110010_01100011_11010101_0;
      patterns[29286] = 25'b01110010_01100100_11010110_0;
      patterns[29287] = 25'b01110010_01100101_11010111_0;
      patterns[29288] = 25'b01110010_01100110_11011000_0;
      patterns[29289] = 25'b01110010_01100111_11011001_0;
      patterns[29290] = 25'b01110010_01101000_11011010_0;
      patterns[29291] = 25'b01110010_01101001_11011011_0;
      patterns[29292] = 25'b01110010_01101010_11011100_0;
      patterns[29293] = 25'b01110010_01101011_11011101_0;
      patterns[29294] = 25'b01110010_01101100_11011110_0;
      patterns[29295] = 25'b01110010_01101101_11011111_0;
      patterns[29296] = 25'b01110010_01101110_11100000_0;
      patterns[29297] = 25'b01110010_01101111_11100001_0;
      patterns[29298] = 25'b01110010_01110000_11100010_0;
      patterns[29299] = 25'b01110010_01110001_11100011_0;
      patterns[29300] = 25'b01110010_01110010_11100100_0;
      patterns[29301] = 25'b01110010_01110011_11100101_0;
      patterns[29302] = 25'b01110010_01110100_11100110_0;
      patterns[29303] = 25'b01110010_01110101_11100111_0;
      patterns[29304] = 25'b01110010_01110110_11101000_0;
      patterns[29305] = 25'b01110010_01110111_11101001_0;
      patterns[29306] = 25'b01110010_01111000_11101010_0;
      patterns[29307] = 25'b01110010_01111001_11101011_0;
      patterns[29308] = 25'b01110010_01111010_11101100_0;
      patterns[29309] = 25'b01110010_01111011_11101101_0;
      patterns[29310] = 25'b01110010_01111100_11101110_0;
      patterns[29311] = 25'b01110010_01111101_11101111_0;
      patterns[29312] = 25'b01110010_01111110_11110000_0;
      patterns[29313] = 25'b01110010_01111111_11110001_0;
      patterns[29314] = 25'b01110010_10000000_11110010_0;
      patterns[29315] = 25'b01110010_10000001_11110011_0;
      patterns[29316] = 25'b01110010_10000010_11110100_0;
      patterns[29317] = 25'b01110010_10000011_11110101_0;
      patterns[29318] = 25'b01110010_10000100_11110110_0;
      patterns[29319] = 25'b01110010_10000101_11110111_0;
      patterns[29320] = 25'b01110010_10000110_11111000_0;
      patterns[29321] = 25'b01110010_10000111_11111001_0;
      patterns[29322] = 25'b01110010_10001000_11111010_0;
      patterns[29323] = 25'b01110010_10001001_11111011_0;
      patterns[29324] = 25'b01110010_10001010_11111100_0;
      patterns[29325] = 25'b01110010_10001011_11111101_0;
      patterns[29326] = 25'b01110010_10001100_11111110_0;
      patterns[29327] = 25'b01110010_10001101_11111111_0;
      patterns[29328] = 25'b01110010_10001110_00000000_1;
      patterns[29329] = 25'b01110010_10001111_00000001_1;
      patterns[29330] = 25'b01110010_10010000_00000010_1;
      patterns[29331] = 25'b01110010_10010001_00000011_1;
      patterns[29332] = 25'b01110010_10010010_00000100_1;
      patterns[29333] = 25'b01110010_10010011_00000101_1;
      patterns[29334] = 25'b01110010_10010100_00000110_1;
      patterns[29335] = 25'b01110010_10010101_00000111_1;
      patterns[29336] = 25'b01110010_10010110_00001000_1;
      patterns[29337] = 25'b01110010_10010111_00001001_1;
      patterns[29338] = 25'b01110010_10011000_00001010_1;
      patterns[29339] = 25'b01110010_10011001_00001011_1;
      patterns[29340] = 25'b01110010_10011010_00001100_1;
      patterns[29341] = 25'b01110010_10011011_00001101_1;
      patterns[29342] = 25'b01110010_10011100_00001110_1;
      patterns[29343] = 25'b01110010_10011101_00001111_1;
      patterns[29344] = 25'b01110010_10011110_00010000_1;
      patterns[29345] = 25'b01110010_10011111_00010001_1;
      patterns[29346] = 25'b01110010_10100000_00010010_1;
      patterns[29347] = 25'b01110010_10100001_00010011_1;
      patterns[29348] = 25'b01110010_10100010_00010100_1;
      patterns[29349] = 25'b01110010_10100011_00010101_1;
      patterns[29350] = 25'b01110010_10100100_00010110_1;
      patterns[29351] = 25'b01110010_10100101_00010111_1;
      patterns[29352] = 25'b01110010_10100110_00011000_1;
      patterns[29353] = 25'b01110010_10100111_00011001_1;
      patterns[29354] = 25'b01110010_10101000_00011010_1;
      patterns[29355] = 25'b01110010_10101001_00011011_1;
      patterns[29356] = 25'b01110010_10101010_00011100_1;
      patterns[29357] = 25'b01110010_10101011_00011101_1;
      patterns[29358] = 25'b01110010_10101100_00011110_1;
      patterns[29359] = 25'b01110010_10101101_00011111_1;
      patterns[29360] = 25'b01110010_10101110_00100000_1;
      patterns[29361] = 25'b01110010_10101111_00100001_1;
      patterns[29362] = 25'b01110010_10110000_00100010_1;
      patterns[29363] = 25'b01110010_10110001_00100011_1;
      patterns[29364] = 25'b01110010_10110010_00100100_1;
      patterns[29365] = 25'b01110010_10110011_00100101_1;
      patterns[29366] = 25'b01110010_10110100_00100110_1;
      patterns[29367] = 25'b01110010_10110101_00100111_1;
      patterns[29368] = 25'b01110010_10110110_00101000_1;
      patterns[29369] = 25'b01110010_10110111_00101001_1;
      patterns[29370] = 25'b01110010_10111000_00101010_1;
      patterns[29371] = 25'b01110010_10111001_00101011_1;
      patterns[29372] = 25'b01110010_10111010_00101100_1;
      patterns[29373] = 25'b01110010_10111011_00101101_1;
      patterns[29374] = 25'b01110010_10111100_00101110_1;
      patterns[29375] = 25'b01110010_10111101_00101111_1;
      patterns[29376] = 25'b01110010_10111110_00110000_1;
      patterns[29377] = 25'b01110010_10111111_00110001_1;
      patterns[29378] = 25'b01110010_11000000_00110010_1;
      patterns[29379] = 25'b01110010_11000001_00110011_1;
      patterns[29380] = 25'b01110010_11000010_00110100_1;
      patterns[29381] = 25'b01110010_11000011_00110101_1;
      patterns[29382] = 25'b01110010_11000100_00110110_1;
      patterns[29383] = 25'b01110010_11000101_00110111_1;
      patterns[29384] = 25'b01110010_11000110_00111000_1;
      patterns[29385] = 25'b01110010_11000111_00111001_1;
      patterns[29386] = 25'b01110010_11001000_00111010_1;
      patterns[29387] = 25'b01110010_11001001_00111011_1;
      patterns[29388] = 25'b01110010_11001010_00111100_1;
      patterns[29389] = 25'b01110010_11001011_00111101_1;
      patterns[29390] = 25'b01110010_11001100_00111110_1;
      patterns[29391] = 25'b01110010_11001101_00111111_1;
      patterns[29392] = 25'b01110010_11001110_01000000_1;
      patterns[29393] = 25'b01110010_11001111_01000001_1;
      patterns[29394] = 25'b01110010_11010000_01000010_1;
      patterns[29395] = 25'b01110010_11010001_01000011_1;
      patterns[29396] = 25'b01110010_11010010_01000100_1;
      patterns[29397] = 25'b01110010_11010011_01000101_1;
      patterns[29398] = 25'b01110010_11010100_01000110_1;
      patterns[29399] = 25'b01110010_11010101_01000111_1;
      patterns[29400] = 25'b01110010_11010110_01001000_1;
      patterns[29401] = 25'b01110010_11010111_01001001_1;
      patterns[29402] = 25'b01110010_11011000_01001010_1;
      patterns[29403] = 25'b01110010_11011001_01001011_1;
      patterns[29404] = 25'b01110010_11011010_01001100_1;
      patterns[29405] = 25'b01110010_11011011_01001101_1;
      patterns[29406] = 25'b01110010_11011100_01001110_1;
      patterns[29407] = 25'b01110010_11011101_01001111_1;
      patterns[29408] = 25'b01110010_11011110_01010000_1;
      patterns[29409] = 25'b01110010_11011111_01010001_1;
      patterns[29410] = 25'b01110010_11100000_01010010_1;
      patterns[29411] = 25'b01110010_11100001_01010011_1;
      patterns[29412] = 25'b01110010_11100010_01010100_1;
      patterns[29413] = 25'b01110010_11100011_01010101_1;
      patterns[29414] = 25'b01110010_11100100_01010110_1;
      patterns[29415] = 25'b01110010_11100101_01010111_1;
      patterns[29416] = 25'b01110010_11100110_01011000_1;
      patterns[29417] = 25'b01110010_11100111_01011001_1;
      patterns[29418] = 25'b01110010_11101000_01011010_1;
      patterns[29419] = 25'b01110010_11101001_01011011_1;
      patterns[29420] = 25'b01110010_11101010_01011100_1;
      patterns[29421] = 25'b01110010_11101011_01011101_1;
      patterns[29422] = 25'b01110010_11101100_01011110_1;
      patterns[29423] = 25'b01110010_11101101_01011111_1;
      patterns[29424] = 25'b01110010_11101110_01100000_1;
      patterns[29425] = 25'b01110010_11101111_01100001_1;
      patterns[29426] = 25'b01110010_11110000_01100010_1;
      patterns[29427] = 25'b01110010_11110001_01100011_1;
      patterns[29428] = 25'b01110010_11110010_01100100_1;
      patterns[29429] = 25'b01110010_11110011_01100101_1;
      patterns[29430] = 25'b01110010_11110100_01100110_1;
      patterns[29431] = 25'b01110010_11110101_01100111_1;
      patterns[29432] = 25'b01110010_11110110_01101000_1;
      patterns[29433] = 25'b01110010_11110111_01101001_1;
      patterns[29434] = 25'b01110010_11111000_01101010_1;
      patterns[29435] = 25'b01110010_11111001_01101011_1;
      patterns[29436] = 25'b01110010_11111010_01101100_1;
      patterns[29437] = 25'b01110010_11111011_01101101_1;
      patterns[29438] = 25'b01110010_11111100_01101110_1;
      patterns[29439] = 25'b01110010_11111101_01101111_1;
      patterns[29440] = 25'b01110010_11111110_01110000_1;
      patterns[29441] = 25'b01110010_11111111_01110001_1;
      patterns[29442] = 25'b01110011_00000000_01110011_0;
      patterns[29443] = 25'b01110011_00000001_01110100_0;
      patterns[29444] = 25'b01110011_00000010_01110101_0;
      patterns[29445] = 25'b01110011_00000011_01110110_0;
      patterns[29446] = 25'b01110011_00000100_01110111_0;
      patterns[29447] = 25'b01110011_00000101_01111000_0;
      patterns[29448] = 25'b01110011_00000110_01111001_0;
      patterns[29449] = 25'b01110011_00000111_01111010_0;
      patterns[29450] = 25'b01110011_00001000_01111011_0;
      patterns[29451] = 25'b01110011_00001001_01111100_0;
      patterns[29452] = 25'b01110011_00001010_01111101_0;
      patterns[29453] = 25'b01110011_00001011_01111110_0;
      patterns[29454] = 25'b01110011_00001100_01111111_0;
      patterns[29455] = 25'b01110011_00001101_10000000_0;
      patterns[29456] = 25'b01110011_00001110_10000001_0;
      patterns[29457] = 25'b01110011_00001111_10000010_0;
      patterns[29458] = 25'b01110011_00010000_10000011_0;
      patterns[29459] = 25'b01110011_00010001_10000100_0;
      patterns[29460] = 25'b01110011_00010010_10000101_0;
      patterns[29461] = 25'b01110011_00010011_10000110_0;
      patterns[29462] = 25'b01110011_00010100_10000111_0;
      patterns[29463] = 25'b01110011_00010101_10001000_0;
      patterns[29464] = 25'b01110011_00010110_10001001_0;
      patterns[29465] = 25'b01110011_00010111_10001010_0;
      patterns[29466] = 25'b01110011_00011000_10001011_0;
      patterns[29467] = 25'b01110011_00011001_10001100_0;
      patterns[29468] = 25'b01110011_00011010_10001101_0;
      patterns[29469] = 25'b01110011_00011011_10001110_0;
      patterns[29470] = 25'b01110011_00011100_10001111_0;
      patterns[29471] = 25'b01110011_00011101_10010000_0;
      patterns[29472] = 25'b01110011_00011110_10010001_0;
      patterns[29473] = 25'b01110011_00011111_10010010_0;
      patterns[29474] = 25'b01110011_00100000_10010011_0;
      patterns[29475] = 25'b01110011_00100001_10010100_0;
      patterns[29476] = 25'b01110011_00100010_10010101_0;
      patterns[29477] = 25'b01110011_00100011_10010110_0;
      patterns[29478] = 25'b01110011_00100100_10010111_0;
      patterns[29479] = 25'b01110011_00100101_10011000_0;
      patterns[29480] = 25'b01110011_00100110_10011001_0;
      patterns[29481] = 25'b01110011_00100111_10011010_0;
      patterns[29482] = 25'b01110011_00101000_10011011_0;
      patterns[29483] = 25'b01110011_00101001_10011100_0;
      patterns[29484] = 25'b01110011_00101010_10011101_0;
      patterns[29485] = 25'b01110011_00101011_10011110_0;
      patterns[29486] = 25'b01110011_00101100_10011111_0;
      patterns[29487] = 25'b01110011_00101101_10100000_0;
      patterns[29488] = 25'b01110011_00101110_10100001_0;
      patterns[29489] = 25'b01110011_00101111_10100010_0;
      patterns[29490] = 25'b01110011_00110000_10100011_0;
      patterns[29491] = 25'b01110011_00110001_10100100_0;
      patterns[29492] = 25'b01110011_00110010_10100101_0;
      patterns[29493] = 25'b01110011_00110011_10100110_0;
      patterns[29494] = 25'b01110011_00110100_10100111_0;
      patterns[29495] = 25'b01110011_00110101_10101000_0;
      patterns[29496] = 25'b01110011_00110110_10101001_0;
      patterns[29497] = 25'b01110011_00110111_10101010_0;
      patterns[29498] = 25'b01110011_00111000_10101011_0;
      patterns[29499] = 25'b01110011_00111001_10101100_0;
      patterns[29500] = 25'b01110011_00111010_10101101_0;
      patterns[29501] = 25'b01110011_00111011_10101110_0;
      patterns[29502] = 25'b01110011_00111100_10101111_0;
      patterns[29503] = 25'b01110011_00111101_10110000_0;
      patterns[29504] = 25'b01110011_00111110_10110001_0;
      patterns[29505] = 25'b01110011_00111111_10110010_0;
      patterns[29506] = 25'b01110011_01000000_10110011_0;
      patterns[29507] = 25'b01110011_01000001_10110100_0;
      patterns[29508] = 25'b01110011_01000010_10110101_0;
      patterns[29509] = 25'b01110011_01000011_10110110_0;
      patterns[29510] = 25'b01110011_01000100_10110111_0;
      patterns[29511] = 25'b01110011_01000101_10111000_0;
      patterns[29512] = 25'b01110011_01000110_10111001_0;
      patterns[29513] = 25'b01110011_01000111_10111010_0;
      patterns[29514] = 25'b01110011_01001000_10111011_0;
      patterns[29515] = 25'b01110011_01001001_10111100_0;
      patterns[29516] = 25'b01110011_01001010_10111101_0;
      patterns[29517] = 25'b01110011_01001011_10111110_0;
      patterns[29518] = 25'b01110011_01001100_10111111_0;
      patterns[29519] = 25'b01110011_01001101_11000000_0;
      patterns[29520] = 25'b01110011_01001110_11000001_0;
      patterns[29521] = 25'b01110011_01001111_11000010_0;
      patterns[29522] = 25'b01110011_01010000_11000011_0;
      patterns[29523] = 25'b01110011_01010001_11000100_0;
      patterns[29524] = 25'b01110011_01010010_11000101_0;
      patterns[29525] = 25'b01110011_01010011_11000110_0;
      patterns[29526] = 25'b01110011_01010100_11000111_0;
      patterns[29527] = 25'b01110011_01010101_11001000_0;
      patterns[29528] = 25'b01110011_01010110_11001001_0;
      patterns[29529] = 25'b01110011_01010111_11001010_0;
      patterns[29530] = 25'b01110011_01011000_11001011_0;
      patterns[29531] = 25'b01110011_01011001_11001100_0;
      patterns[29532] = 25'b01110011_01011010_11001101_0;
      patterns[29533] = 25'b01110011_01011011_11001110_0;
      patterns[29534] = 25'b01110011_01011100_11001111_0;
      patterns[29535] = 25'b01110011_01011101_11010000_0;
      patterns[29536] = 25'b01110011_01011110_11010001_0;
      patterns[29537] = 25'b01110011_01011111_11010010_0;
      patterns[29538] = 25'b01110011_01100000_11010011_0;
      patterns[29539] = 25'b01110011_01100001_11010100_0;
      patterns[29540] = 25'b01110011_01100010_11010101_0;
      patterns[29541] = 25'b01110011_01100011_11010110_0;
      patterns[29542] = 25'b01110011_01100100_11010111_0;
      patterns[29543] = 25'b01110011_01100101_11011000_0;
      patterns[29544] = 25'b01110011_01100110_11011001_0;
      patterns[29545] = 25'b01110011_01100111_11011010_0;
      patterns[29546] = 25'b01110011_01101000_11011011_0;
      patterns[29547] = 25'b01110011_01101001_11011100_0;
      patterns[29548] = 25'b01110011_01101010_11011101_0;
      patterns[29549] = 25'b01110011_01101011_11011110_0;
      patterns[29550] = 25'b01110011_01101100_11011111_0;
      patterns[29551] = 25'b01110011_01101101_11100000_0;
      patterns[29552] = 25'b01110011_01101110_11100001_0;
      patterns[29553] = 25'b01110011_01101111_11100010_0;
      patterns[29554] = 25'b01110011_01110000_11100011_0;
      patterns[29555] = 25'b01110011_01110001_11100100_0;
      patterns[29556] = 25'b01110011_01110010_11100101_0;
      patterns[29557] = 25'b01110011_01110011_11100110_0;
      patterns[29558] = 25'b01110011_01110100_11100111_0;
      patterns[29559] = 25'b01110011_01110101_11101000_0;
      patterns[29560] = 25'b01110011_01110110_11101001_0;
      patterns[29561] = 25'b01110011_01110111_11101010_0;
      patterns[29562] = 25'b01110011_01111000_11101011_0;
      patterns[29563] = 25'b01110011_01111001_11101100_0;
      patterns[29564] = 25'b01110011_01111010_11101101_0;
      patterns[29565] = 25'b01110011_01111011_11101110_0;
      patterns[29566] = 25'b01110011_01111100_11101111_0;
      patterns[29567] = 25'b01110011_01111101_11110000_0;
      patterns[29568] = 25'b01110011_01111110_11110001_0;
      patterns[29569] = 25'b01110011_01111111_11110010_0;
      patterns[29570] = 25'b01110011_10000000_11110011_0;
      patterns[29571] = 25'b01110011_10000001_11110100_0;
      patterns[29572] = 25'b01110011_10000010_11110101_0;
      patterns[29573] = 25'b01110011_10000011_11110110_0;
      patterns[29574] = 25'b01110011_10000100_11110111_0;
      patterns[29575] = 25'b01110011_10000101_11111000_0;
      patterns[29576] = 25'b01110011_10000110_11111001_0;
      patterns[29577] = 25'b01110011_10000111_11111010_0;
      patterns[29578] = 25'b01110011_10001000_11111011_0;
      patterns[29579] = 25'b01110011_10001001_11111100_0;
      patterns[29580] = 25'b01110011_10001010_11111101_0;
      patterns[29581] = 25'b01110011_10001011_11111110_0;
      patterns[29582] = 25'b01110011_10001100_11111111_0;
      patterns[29583] = 25'b01110011_10001101_00000000_1;
      patterns[29584] = 25'b01110011_10001110_00000001_1;
      patterns[29585] = 25'b01110011_10001111_00000010_1;
      patterns[29586] = 25'b01110011_10010000_00000011_1;
      patterns[29587] = 25'b01110011_10010001_00000100_1;
      patterns[29588] = 25'b01110011_10010010_00000101_1;
      patterns[29589] = 25'b01110011_10010011_00000110_1;
      patterns[29590] = 25'b01110011_10010100_00000111_1;
      patterns[29591] = 25'b01110011_10010101_00001000_1;
      patterns[29592] = 25'b01110011_10010110_00001001_1;
      patterns[29593] = 25'b01110011_10010111_00001010_1;
      patterns[29594] = 25'b01110011_10011000_00001011_1;
      patterns[29595] = 25'b01110011_10011001_00001100_1;
      patterns[29596] = 25'b01110011_10011010_00001101_1;
      patterns[29597] = 25'b01110011_10011011_00001110_1;
      patterns[29598] = 25'b01110011_10011100_00001111_1;
      patterns[29599] = 25'b01110011_10011101_00010000_1;
      patterns[29600] = 25'b01110011_10011110_00010001_1;
      patterns[29601] = 25'b01110011_10011111_00010010_1;
      patterns[29602] = 25'b01110011_10100000_00010011_1;
      patterns[29603] = 25'b01110011_10100001_00010100_1;
      patterns[29604] = 25'b01110011_10100010_00010101_1;
      patterns[29605] = 25'b01110011_10100011_00010110_1;
      patterns[29606] = 25'b01110011_10100100_00010111_1;
      patterns[29607] = 25'b01110011_10100101_00011000_1;
      patterns[29608] = 25'b01110011_10100110_00011001_1;
      patterns[29609] = 25'b01110011_10100111_00011010_1;
      patterns[29610] = 25'b01110011_10101000_00011011_1;
      patterns[29611] = 25'b01110011_10101001_00011100_1;
      patterns[29612] = 25'b01110011_10101010_00011101_1;
      patterns[29613] = 25'b01110011_10101011_00011110_1;
      patterns[29614] = 25'b01110011_10101100_00011111_1;
      patterns[29615] = 25'b01110011_10101101_00100000_1;
      patterns[29616] = 25'b01110011_10101110_00100001_1;
      patterns[29617] = 25'b01110011_10101111_00100010_1;
      patterns[29618] = 25'b01110011_10110000_00100011_1;
      patterns[29619] = 25'b01110011_10110001_00100100_1;
      patterns[29620] = 25'b01110011_10110010_00100101_1;
      patterns[29621] = 25'b01110011_10110011_00100110_1;
      patterns[29622] = 25'b01110011_10110100_00100111_1;
      patterns[29623] = 25'b01110011_10110101_00101000_1;
      patterns[29624] = 25'b01110011_10110110_00101001_1;
      patterns[29625] = 25'b01110011_10110111_00101010_1;
      patterns[29626] = 25'b01110011_10111000_00101011_1;
      patterns[29627] = 25'b01110011_10111001_00101100_1;
      patterns[29628] = 25'b01110011_10111010_00101101_1;
      patterns[29629] = 25'b01110011_10111011_00101110_1;
      patterns[29630] = 25'b01110011_10111100_00101111_1;
      patterns[29631] = 25'b01110011_10111101_00110000_1;
      patterns[29632] = 25'b01110011_10111110_00110001_1;
      patterns[29633] = 25'b01110011_10111111_00110010_1;
      patterns[29634] = 25'b01110011_11000000_00110011_1;
      patterns[29635] = 25'b01110011_11000001_00110100_1;
      patterns[29636] = 25'b01110011_11000010_00110101_1;
      patterns[29637] = 25'b01110011_11000011_00110110_1;
      patterns[29638] = 25'b01110011_11000100_00110111_1;
      patterns[29639] = 25'b01110011_11000101_00111000_1;
      patterns[29640] = 25'b01110011_11000110_00111001_1;
      patterns[29641] = 25'b01110011_11000111_00111010_1;
      patterns[29642] = 25'b01110011_11001000_00111011_1;
      patterns[29643] = 25'b01110011_11001001_00111100_1;
      patterns[29644] = 25'b01110011_11001010_00111101_1;
      patterns[29645] = 25'b01110011_11001011_00111110_1;
      patterns[29646] = 25'b01110011_11001100_00111111_1;
      patterns[29647] = 25'b01110011_11001101_01000000_1;
      patterns[29648] = 25'b01110011_11001110_01000001_1;
      patterns[29649] = 25'b01110011_11001111_01000010_1;
      patterns[29650] = 25'b01110011_11010000_01000011_1;
      patterns[29651] = 25'b01110011_11010001_01000100_1;
      patterns[29652] = 25'b01110011_11010010_01000101_1;
      patterns[29653] = 25'b01110011_11010011_01000110_1;
      patterns[29654] = 25'b01110011_11010100_01000111_1;
      patterns[29655] = 25'b01110011_11010101_01001000_1;
      patterns[29656] = 25'b01110011_11010110_01001001_1;
      patterns[29657] = 25'b01110011_11010111_01001010_1;
      patterns[29658] = 25'b01110011_11011000_01001011_1;
      patterns[29659] = 25'b01110011_11011001_01001100_1;
      patterns[29660] = 25'b01110011_11011010_01001101_1;
      patterns[29661] = 25'b01110011_11011011_01001110_1;
      patterns[29662] = 25'b01110011_11011100_01001111_1;
      patterns[29663] = 25'b01110011_11011101_01010000_1;
      patterns[29664] = 25'b01110011_11011110_01010001_1;
      patterns[29665] = 25'b01110011_11011111_01010010_1;
      patterns[29666] = 25'b01110011_11100000_01010011_1;
      patterns[29667] = 25'b01110011_11100001_01010100_1;
      patterns[29668] = 25'b01110011_11100010_01010101_1;
      patterns[29669] = 25'b01110011_11100011_01010110_1;
      patterns[29670] = 25'b01110011_11100100_01010111_1;
      patterns[29671] = 25'b01110011_11100101_01011000_1;
      patterns[29672] = 25'b01110011_11100110_01011001_1;
      patterns[29673] = 25'b01110011_11100111_01011010_1;
      patterns[29674] = 25'b01110011_11101000_01011011_1;
      patterns[29675] = 25'b01110011_11101001_01011100_1;
      patterns[29676] = 25'b01110011_11101010_01011101_1;
      patterns[29677] = 25'b01110011_11101011_01011110_1;
      patterns[29678] = 25'b01110011_11101100_01011111_1;
      patterns[29679] = 25'b01110011_11101101_01100000_1;
      patterns[29680] = 25'b01110011_11101110_01100001_1;
      patterns[29681] = 25'b01110011_11101111_01100010_1;
      patterns[29682] = 25'b01110011_11110000_01100011_1;
      patterns[29683] = 25'b01110011_11110001_01100100_1;
      patterns[29684] = 25'b01110011_11110010_01100101_1;
      patterns[29685] = 25'b01110011_11110011_01100110_1;
      patterns[29686] = 25'b01110011_11110100_01100111_1;
      patterns[29687] = 25'b01110011_11110101_01101000_1;
      patterns[29688] = 25'b01110011_11110110_01101001_1;
      patterns[29689] = 25'b01110011_11110111_01101010_1;
      patterns[29690] = 25'b01110011_11111000_01101011_1;
      patterns[29691] = 25'b01110011_11111001_01101100_1;
      patterns[29692] = 25'b01110011_11111010_01101101_1;
      patterns[29693] = 25'b01110011_11111011_01101110_1;
      patterns[29694] = 25'b01110011_11111100_01101111_1;
      patterns[29695] = 25'b01110011_11111101_01110000_1;
      patterns[29696] = 25'b01110011_11111110_01110001_1;
      patterns[29697] = 25'b01110011_11111111_01110010_1;
      patterns[29698] = 25'b01110100_00000000_01110100_0;
      patterns[29699] = 25'b01110100_00000001_01110101_0;
      patterns[29700] = 25'b01110100_00000010_01110110_0;
      patterns[29701] = 25'b01110100_00000011_01110111_0;
      patterns[29702] = 25'b01110100_00000100_01111000_0;
      patterns[29703] = 25'b01110100_00000101_01111001_0;
      patterns[29704] = 25'b01110100_00000110_01111010_0;
      patterns[29705] = 25'b01110100_00000111_01111011_0;
      patterns[29706] = 25'b01110100_00001000_01111100_0;
      patterns[29707] = 25'b01110100_00001001_01111101_0;
      patterns[29708] = 25'b01110100_00001010_01111110_0;
      patterns[29709] = 25'b01110100_00001011_01111111_0;
      patterns[29710] = 25'b01110100_00001100_10000000_0;
      patterns[29711] = 25'b01110100_00001101_10000001_0;
      patterns[29712] = 25'b01110100_00001110_10000010_0;
      patterns[29713] = 25'b01110100_00001111_10000011_0;
      patterns[29714] = 25'b01110100_00010000_10000100_0;
      patterns[29715] = 25'b01110100_00010001_10000101_0;
      patterns[29716] = 25'b01110100_00010010_10000110_0;
      patterns[29717] = 25'b01110100_00010011_10000111_0;
      patterns[29718] = 25'b01110100_00010100_10001000_0;
      patterns[29719] = 25'b01110100_00010101_10001001_0;
      patterns[29720] = 25'b01110100_00010110_10001010_0;
      patterns[29721] = 25'b01110100_00010111_10001011_0;
      patterns[29722] = 25'b01110100_00011000_10001100_0;
      patterns[29723] = 25'b01110100_00011001_10001101_0;
      patterns[29724] = 25'b01110100_00011010_10001110_0;
      patterns[29725] = 25'b01110100_00011011_10001111_0;
      patterns[29726] = 25'b01110100_00011100_10010000_0;
      patterns[29727] = 25'b01110100_00011101_10010001_0;
      patterns[29728] = 25'b01110100_00011110_10010010_0;
      patterns[29729] = 25'b01110100_00011111_10010011_0;
      patterns[29730] = 25'b01110100_00100000_10010100_0;
      patterns[29731] = 25'b01110100_00100001_10010101_0;
      patterns[29732] = 25'b01110100_00100010_10010110_0;
      patterns[29733] = 25'b01110100_00100011_10010111_0;
      patterns[29734] = 25'b01110100_00100100_10011000_0;
      patterns[29735] = 25'b01110100_00100101_10011001_0;
      patterns[29736] = 25'b01110100_00100110_10011010_0;
      patterns[29737] = 25'b01110100_00100111_10011011_0;
      patterns[29738] = 25'b01110100_00101000_10011100_0;
      patterns[29739] = 25'b01110100_00101001_10011101_0;
      patterns[29740] = 25'b01110100_00101010_10011110_0;
      patterns[29741] = 25'b01110100_00101011_10011111_0;
      patterns[29742] = 25'b01110100_00101100_10100000_0;
      patterns[29743] = 25'b01110100_00101101_10100001_0;
      patterns[29744] = 25'b01110100_00101110_10100010_0;
      patterns[29745] = 25'b01110100_00101111_10100011_0;
      patterns[29746] = 25'b01110100_00110000_10100100_0;
      patterns[29747] = 25'b01110100_00110001_10100101_0;
      patterns[29748] = 25'b01110100_00110010_10100110_0;
      patterns[29749] = 25'b01110100_00110011_10100111_0;
      patterns[29750] = 25'b01110100_00110100_10101000_0;
      patterns[29751] = 25'b01110100_00110101_10101001_0;
      patterns[29752] = 25'b01110100_00110110_10101010_0;
      patterns[29753] = 25'b01110100_00110111_10101011_0;
      patterns[29754] = 25'b01110100_00111000_10101100_0;
      patterns[29755] = 25'b01110100_00111001_10101101_0;
      patterns[29756] = 25'b01110100_00111010_10101110_0;
      patterns[29757] = 25'b01110100_00111011_10101111_0;
      patterns[29758] = 25'b01110100_00111100_10110000_0;
      patterns[29759] = 25'b01110100_00111101_10110001_0;
      patterns[29760] = 25'b01110100_00111110_10110010_0;
      patterns[29761] = 25'b01110100_00111111_10110011_0;
      patterns[29762] = 25'b01110100_01000000_10110100_0;
      patterns[29763] = 25'b01110100_01000001_10110101_0;
      patterns[29764] = 25'b01110100_01000010_10110110_0;
      patterns[29765] = 25'b01110100_01000011_10110111_0;
      patterns[29766] = 25'b01110100_01000100_10111000_0;
      patterns[29767] = 25'b01110100_01000101_10111001_0;
      patterns[29768] = 25'b01110100_01000110_10111010_0;
      patterns[29769] = 25'b01110100_01000111_10111011_0;
      patterns[29770] = 25'b01110100_01001000_10111100_0;
      patterns[29771] = 25'b01110100_01001001_10111101_0;
      patterns[29772] = 25'b01110100_01001010_10111110_0;
      patterns[29773] = 25'b01110100_01001011_10111111_0;
      patterns[29774] = 25'b01110100_01001100_11000000_0;
      patterns[29775] = 25'b01110100_01001101_11000001_0;
      patterns[29776] = 25'b01110100_01001110_11000010_0;
      patterns[29777] = 25'b01110100_01001111_11000011_0;
      patterns[29778] = 25'b01110100_01010000_11000100_0;
      patterns[29779] = 25'b01110100_01010001_11000101_0;
      patterns[29780] = 25'b01110100_01010010_11000110_0;
      patterns[29781] = 25'b01110100_01010011_11000111_0;
      patterns[29782] = 25'b01110100_01010100_11001000_0;
      patterns[29783] = 25'b01110100_01010101_11001001_0;
      patterns[29784] = 25'b01110100_01010110_11001010_0;
      patterns[29785] = 25'b01110100_01010111_11001011_0;
      patterns[29786] = 25'b01110100_01011000_11001100_0;
      patterns[29787] = 25'b01110100_01011001_11001101_0;
      patterns[29788] = 25'b01110100_01011010_11001110_0;
      patterns[29789] = 25'b01110100_01011011_11001111_0;
      patterns[29790] = 25'b01110100_01011100_11010000_0;
      patterns[29791] = 25'b01110100_01011101_11010001_0;
      patterns[29792] = 25'b01110100_01011110_11010010_0;
      patterns[29793] = 25'b01110100_01011111_11010011_0;
      patterns[29794] = 25'b01110100_01100000_11010100_0;
      patterns[29795] = 25'b01110100_01100001_11010101_0;
      patterns[29796] = 25'b01110100_01100010_11010110_0;
      patterns[29797] = 25'b01110100_01100011_11010111_0;
      patterns[29798] = 25'b01110100_01100100_11011000_0;
      patterns[29799] = 25'b01110100_01100101_11011001_0;
      patterns[29800] = 25'b01110100_01100110_11011010_0;
      patterns[29801] = 25'b01110100_01100111_11011011_0;
      patterns[29802] = 25'b01110100_01101000_11011100_0;
      patterns[29803] = 25'b01110100_01101001_11011101_0;
      patterns[29804] = 25'b01110100_01101010_11011110_0;
      patterns[29805] = 25'b01110100_01101011_11011111_0;
      patterns[29806] = 25'b01110100_01101100_11100000_0;
      patterns[29807] = 25'b01110100_01101101_11100001_0;
      patterns[29808] = 25'b01110100_01101110_11100010_0;
      patterns[29809] = 25'b01110100_01101111_11100011_0;
      patterns[29810] = 25'b01110100_01110000_11100100_0;
      patterns[29811] = 25'b01110100_01110001_11100101_0;
      patterns[29812] = 25'b01110100_01110010_11100110_0;
      patterns[29813] = 25'b01110100_01110011_11100111_0;
      patterns[29814] = 25'b01110100_01110100_11101000_0;
      patterns[29815] = 25'b01110100_01110101_11101001_0;
      patterns[29816] = 25'b01110100_01110110_11101010_0;
      patterns[29817] = 25'b01110100_01110111_11101011_0;
      patterns[29818] = 25'b01110100_01111000_11101100_0;
      patterns[29819] = 25'b01110100_01111001_11101101_0;
      patterns[29820] = 25'b01110100_01111010_11101110_0;
      patterns[29821] = 25'b01110100_01111011_11101111_0;
      patterns[29822] = 25'b01110100_01111100_11110000_0;
      patterns[29823] = 25'b01110100_01111101_11110001_0;
      patterns[29824] = 25'b01110100_01111110_11110010_0;
      patterns[29825] = 25'b01110100_01111111_11110011_0;
      patterns[29826] = 25'b01110100_10000000_11110100_0;
      patterns[29827] = 25'b01110100_10000001_11110101_0;
      patterns[29828] = 25'b01110100_10000010_11110110_0;
      patterns[29829] = 25'b01110100_10000011_11110111_0;
      patterns[29830] = 25'b01110100_10000100_11111000_0;
      patterns[29831] = 25'b01110100_10000101_11111001_0;
      patterns[29832] = 25'b01110100_10000110_11111010_0;
      patterns[29833] = 25'b01110100_10000111_11111011_0;
      patterns[29834] = 25'b01110100_10001000_11111100_0;
      patterns[29835] = 25'b01110100_10001001_11111101_0;
      patterns[29836] = 25'b01110100_10001010_11111110_0;
      patterns[29837] = 25'b01110100_10001011_11111111_0;
      patterns[29838] = 25'b01110100_10001100_00000000_1;
      patterns[29839] = 25'b01110100_10001101_00000001_1;
      patterns[29840] = 25'b01110100_10001110_00000010_1;
      patterns[29841] = 25'b01110100_10001111_00000011_1;
      patterns[29842] = 25'b01110100_10010000_00000100_1;
      patterns[29843] = 25'b01110100_10010001_00000101_1;
      patterns[29844] = 25'b01110100_10010010_00000110_1;
      patterns[29845] = 25'b01110100_10010011_00000111_1;
      patterns[29846] = 25'b01110100_10010100_00001000_1;
      patterns[29847] = 25'b01110100_10010101_00001001_1;
      patterns[29848] = 25'b01110100_10010110_00001010_1;
      patterns[29849] = 25'b01110100_10010111_00001011_1;
      patterns[29850] = 25'b01110100_10011000_00001100_1;
      patterns[29851] = 25'b01110100_10011001_00001101_1;
      patterns[29852] = 25'b01110100_10011010_00001110_1;
      patterns[29853] = 25'b01110100_10011011_00001111_1;
      patterns[29854] = 25'b01110100_10011100_00010000_1;
      patterns[29855] = 25'b01110100_10011101_00010001_1;
      patterns[29856] = 25'b01110100_10011110_00010010_1;
      patterns[29857] = 25'b01110100_10011111_00010011_1;
      patterns[29858] = 25'b01110100_10100000_00010100_1;
      patterns[29859] = 25'b01110100_10100001_00010101_1;
      patterns[29860] = 25'b01110100_10100010_00010110_1;
      patterns[29861] = 25'b01110100_10100011_00010111_1;
      patterns[29862] = 25'b01110100_10100100_00011000_1;
      patterns[29863] = 25'b01110100_10100101_00011001_1;
      patterns[29864] = 25'b01110100_10100110_00011010_1;
      patterns[29865] = 25'b01110100_10100111_00011011_1;
      patterns[29866] = 25'b01110100_10101000_00011100_1;
      patterns[29867] = 25'b01110100_10101001_00011101_1;
      patterns[29868] = 25'b01110100_10101010_00011110_1;
      patterns[29869] = 25'b01110100_10101011_00011111_1;
      patterns[29870] = 25'b01110100_10101100_00100000_1;
      patterns[29871] = 25'b01110100_10101101_00100001_1;
      patterns[29872] = 25'b01110100_10101110_00100010_1;
      patterns[29873] = 25'b01110100_10101111_00100011_1;
      patterns[29874] = 25'b01110100_10110000_00100100_1;
      patterns[29875] = 25'b01110100_10110001_00100101_1;
      patterns[29876] = 25'b01110100_10110010_00100110_1;
      patterns[29877] = 25'b01110100_10110011_00100111_1;
      patterns[29878] = 25'b01110100_10110100_00101000_1;
      patterns[29879] = 25'b01110100_10110101_00101001_1;
      patterns[29880] = 25'b01110100_10110110_00101010_1;
      patterns[29881] = 25'b01110100_10110111_00101011_1;
      patterns[29882] = 25'b01110100_10111000_00101100_1;
      patterns[29883] = 25'b01110100_10111001_00101101_1;
      patterns[29884] = 25'b01110100_10111010_00101110_1;
      patterns[29885] = 25'b01110100_10111011_00101111_1;
      patterns[29886] = 25'b01110100_10111100_00110000_1;
      patterns[29887] = 25'b01110100_10111101_00110001_1;
      patterns[29888] = 25'b01110100_10111110_00110010_1;
      patterns[29889] = 25'b01110100_10111111_00110011_1;
      patterns[29890] = 25'b01110100_11000000_00110100_1;
      patterns[29891] = 25'b01110100_11000001_00110101_1;
      patterns[29892] = 25'b01110100_11000010_00110110_1;
      patterns[29893] = 25'b01110100_11000011_00110111_1;
      patterns[29894] = 25'b01110100_11000100_00111000_1;
      patterns[29895] = 25'b01110100_11000101_00111001_1;
      patterns[29896] = 25'b01110100_11000110_00111010_1;
      patterns[29897] = 25'b01110100_11000111_00111011_1;
      patterns[29898] = 25'b01110100_11001000_00111100_1;
      patterns[29899] = 25'b01110100_11001001_00111101_1;
      patterns[29900] = 25'b01110100_11001010_00111110_1;
      patterns[29901] = 25'b01110100_11001011_00111111_1;
      patterns[29902] = 25'b01110100_11001100_01000000_1;
      patterns[29903] = 25'b01110100_11001101_01000001_1;
      patterns[29904] = 25'b01110100_11001110_01000010_1;
      patterns[29905] = 25'b01110100_11001111_01000011_1;
      patterns[29906] = 25'b01110100_11010000_01000100_1;
      patterns[29907] = 25'b01110100_11010001_01000101_1;
      patterns[29908] = 25'b01110100_11010010_01000110_1;
      patterns[29909] = 25'b01110100_11010011_01000111_1;
      patterns[29910] = 25'b01110100_11010100_01001000_1;
      patterns[29911] = 25'b01110100_11010101_01001001_1;
      patterns[29912] = 25'b01110100_11010110_01001010_1;
      patterns[29913] = 25'b01110100_11010111_01001011_1;
      patterns[29914] = 25'b01110100_11011000_01001100_1;
      patterns[29915] = 25'b01110100_11011001_01001101_1;
      patterns[29916] = 25'b01110100_11011010_01001110_1;
      patterns[29917] = 25'b01110100_11011011_01001111_1;
      patterns[29918] = 25'b01110100_11011100_01010000_1;
      patterns[29919] = 25'b01110100_11011101_01010001_1;
      patterns[29920] = 25'b01110100_11011110_01010010_1;
      patterns[29921] = 25'b01110100_11011111_01010011_1;
      patterns[29922] = 25'b01110100_11100000_01010100_1;
      patterns[29923] = 25'b01110100_11100001_01010101_1;
      patterns[29924] = 25'b01110100_11100010_01010110_1;
      patterns[29925] = 25'b01110100_11100011_01010111_1;
      patterns[29926] = 25'b01110100_11100100_01011000_1;
      patterns[29927] = 25'b01110100_11100101_01011001_1;
      patterns[29928] = 25'b01110100_11100110_01011010_1;
      patterns[29929] = 25'b01110100_11100111_01011011_1;
      patterns[29930] = 25'b01110100_11101000_01011100_1;
      patterns[29931] = 25'b01110100_11101001_01011101_1;
      patterns[29932] = 25'b01110100_11101010_01011110_1;
      patterns[29933] = 25'b01110100_11101011_01011111_1;
      patterns[29934] = 25'b01110100_11101100_01100000_1;
      patterns[29935] = 25'b01110100_11101101_01100001_1;
      patterns[29936] = 25'b01110100_11101110_01100010_1;
      patterns[29937] = 25'b01110100_11101111_01100011_1;
      patterns[29938] = 25'b01110100_11110000_01100100_1;
      patterns[29939] = 25'b01110100_11110001_01100101_1;
      patterns[29940] = 25'b01110100_11110010_01100110_1;
      patterns[29941] = 25'b01110100_11110011_01100111_1;
      patterns[29942] = 25'b01110100_11110100_01101000_1;
      patterns[29943] = 25'b01110100_11110101_01101001_1;
      patterns[29944] = 25'b01110100_11110110_01101010_1;
      patterns[29945] = 25'b01110100_11110111_01101011_1;
      patterns[29946] = 25'b01110100_11111000_01101100_1;
      patterns[29947] = 25'b01110100_11111001_01101101_1;
      patterns[29948] = 25'b01110100_11111010_01101110_1;
      patterns[29949] = 25'b01110100_11111011_01101111_1;
      patterns[29950] = 25'b01110100_11111100_01110000_1;
      patterns[29951] = 25'b01110100_11111101_01110001_1;
      patterns[29952] = 25'b01110100_11111110_01110010_1;
      patterns[29953] = 25'b01110100_11111111_01110011_1;
      patterns[29954] = 25'b01110101_00000000_01110101_0;
      patterns[29955] = 25'b01110101_00000001_01110110_0;
      patterns[29956] = 25'b01110101_00000010_01110111_0;
      patterns[29957] = 25'b01110101_00000011_01111000_0;
      patterns[29958] = 25'b01110101_00000100_01111001_0;
      patterns[29959] = 25'b01110101_00000101_01111010_0;
      patterns[29960] = 25'b01110101_00000110_01111011_0;
      patterns[29961] = 25'b01110101_00000111_01111100_0;
      patterns[29962] = 25'b01110101_00001000_01111101_0;
      patterns[29963] = 25'b01110101_00001001_01111110_0;
      patterns[29964] = 25'b01110101_00001010_01111111_0;
      patterns[29965] = 25'b01110101_00001011_10000000_0;
      patterns[29966] = 25'b01110101_00001100_10000001_0;
      patterns[29967] = 25'b01110101_00001101_10000010_0;
      patterns[29968] = 25'b01110101_00001110_10000011_0;
      patterns[29969] = 25'b01110101_00001111_10000100_0;
      patterns[29970] = 25'b01110101_00010000_10000101_0;
      patterns[29971] = 25'b01110101_00010001_10000110_0;
      patterns[29972] = 25'b01110101_00010010_10000111_0;
      patterns[29973] = 25'b01110101_00010011_10001000_0;
      patterns[29974] = 25'b01110101_00010100_10001001_0;
      patterns[29975] = 25'b01110101_00010101_10001010_0;
      patterns[29976] = 25'b01110101_00010110_10001011_0;
      patterns[29977] = 25'b01110101_00010111_10001100_0;
      patterns[29978] = 25'b01110101_00011000_10001101_0;
      patterns[29979] = 25'b01110101_00011001_10001110_0;
      patterns[29980] = 25'b01110101_00011010_10001111_0;
      patterns[29981] = 25'b01110101_00011011_10010000_0;
      patterns[29982] = 25'b01110101_00011100_10010001_0;
      patterns[29983] = 25'b01110101_00011101_10010010_0;
      patterns[29984] = 25'b01110101_00011110_10010011_0;
      patterns[29985] = 25'b01110101_00011111_10010100_0;
      patterns[29986] = 25'b01110101_00100000_10010101_0;
      patterns[29987] = 25'b01110101_00100001_10010110_0;
      patterns[29988] = 25'b01110101_00100010_10010111_0;
      patterns[29989] = 25'b01110101_00100011_10011000_0;
      patterns[29990] = 25'b01110101_00100100_10011001_0;
      patterns[29991] = 25'b01110101_00100101_10011010_0;
      patterns[29992] = 25'b01110101_00100110_10011011_0;
      patterns[29993] = 25'b01110101_00100111_10011100_0;
      patterns[29994] = 25'b01110101_00101000_10011101_0;
      patterns[29995] = 25'b01110101_00101001_10011110_0;
      patterns[29996] = 25'b01110101_00101010_10011111_0;
      patterns[29997] = 25'b01110101_00101011_10100000_0;
      patterns[29998] = 25'b01110101_00101100_10100001_0;
      patterns[29999] = 25'b01110101_00101101_10100010_0;
      patterns[30000] = 25'b01110101_00101110_10100011_0;
      patterns[30001] = 25'b01110101_00101111_10100100_0;
      patterns[30002] = 25'b01110101_00110000_10100101_0;
      patterns[30003] = 25'b01110101_00110001_10100110_0;
      patterns[30004] = 25'b01110101_00110010_10100111_0;
      patterns[30005] = 25'b01110101_00110011_10101000_0;
      patterns[30006] = 25'b01110101_00110100_10101001_0;
      patterns[30007] = 25'b01110101_00110101_10101010_0;
      patterns[30008] = 25'b01110101_00110110_10101011_0;
      patterns[30009] = 25'b01110101_00110111_10101100_0;
      patterns[30010] = 25'b01110101_00111000_10101101_0;
      patterns[30011] = 25'b01110101_00111001_10101110_0;
      patterns[30012] = 25'b01110101_00111010_10101111_0;
      patterns[30013] = 25'b01110101_00111011_10110000_0;
      patterns[30014] = 25'b01110101_00111100_10110001_0;
      patterns[30015] = 25'b01110101_00111101_10110010_0;
      patterns[30016] = 25'b01110101_00111110_10110011_0;
      patterns[30017] = 25'b01110101_00111111_10110100_0;
      patterns[30018] = 25'b01110101_01000000_10110101_0;
      patterns[30019] = 25'b01110101_01000001_10110110_0;
      patterns[30020] = 25'b01110101_01000010_10110111_0;
      patterns[30021] = 25'b01110101_01000011_10111000_0;
      patterns[30022] = 25'b01110101_01000100_10111001_0;
      patterns[30023] = 25'b01110101_01000101_10111010_0;
      patterns[30024] = 25'b01110101_01000110_10111011_0;
      patterns[30025] = 25'b01110101_01000111_10111100_0;
      patterns[30026] = 25'b01110101_01001000_10111101_0;
      patterns[30027] = 25'b01110101_01001001_10111110_0;
      patterns[30028] = 25'b01110101_01001010_10111111_0;
      patterns[30029] = 25'b01110101_01001011_11000000_0;
      patterns[30030] = 25'b01110101_01001100_11000001_0;
      patterns[30031] = 25'b01110101_01001101_11000010_0;
      patterns[30032] = 25'b01110101_01001110_11000011_0;
      patterns[30033] = 25'b01110101_01001111_11000100_0;
      patterns[30034] = 25'b01110101_01010000_11000101_0;
      patterns[30035] = 25'b01110101_01010001_11000110_0;
      patterns[30036] = 25'b01110101_01010010_11000111_0;
      patterns[30037] = 25'b01110101_01010011_11001000_0;
      patterns[30038] = 25'b01110101_01010100_11001001_0;
      patterns[30039] = 25'b01110101_01010101_11001010_0;
      patterns[30040] = 25'b01110101_01010110_11001011_0;
      patterns[30041] = 25'b01110101_01010111_11001100_0;
      patterns[30042] = 25'b01110101_01011000_11001101_0;
      patterns[30043] = 25'b01110101_01011001_11001110_0;
      patterns[30044] = 25'b01110101_01011010_11001111_0;
      patterns[30045] = 25'b01110101_01011011_11010000_0;
      patterns[30046] = 25'b01110101_01011100_11010001_0;
      patterns[30047] = 25'b01110101_01011101_11010010_0;
      patterns[30048] = 25'b01110101_01011110_11010011_0;
      patterns[30049] = 25'b01110101_01011111_11010100_0;
      patterns[30050] = 25'b01110101_01100000_11010101_0;
      patterns[30051] = 25'b01110101_01100001_11010110_0;
      patterns[30052] = 25'b01110101_01100010_11010111_0;
      patterns[30053] = 25'b01110101_01100011_11011000_0;
      patterns[30054] = 25'b01110101_01100100_11011001_0;
      patterns[30055] = 25'b01110101_01100101_11011010_0;
      patterns[30056] = 25'b01110101_01100110_11011011_0;
      patterns[30057] = 25'b01110101_01100111_11011100_0;
      patterns[30058] = 25'b01110101_01101000_11011101_0;
      patterns[30059] = 25'b01110101_01101001_11011110_0;
      patterns[30060] = 25'b01110101_01101010_11011111_0;
      patterns[30061] = 25'b01110101_01101011_11100000_0;
      patterns[30062] = 25'b01110101_01101100_11100001_0;
      patterns[30063] = 25'b01110101_01101101_11100010_0;
      patterns[30064] = 25'b01110101_01101110_11100011_0;
      patterns[30065] = 25'b01110101_01101111_11100100_0;
      patterns[30066] = 25'b01110101_01110000_11100101_0;
      patterns[30067] = 25'b01110101_01110001_11100110_0;
      patterns[30068] = 25'b01110101_01110010_11100111_0;
      patterns[30069] = 25'b01110101_01110011_11101000_0;
      patterns[30070] = 25'b01110101_01110100_11101001_0;
      patterns[30071] = 25'b01110101_01110101_11101010_0;
      patterns[30072] = 25'b01110101_01110110_11101011_0;
      patterns[30073] = 25'b01110101_01110111_11101100_0;
      patterns[30074] = 25'b01110101_01111000_11101101_0;
      patterns[30075] = 25'b01110101_01111001_11101110_0;
      patterns[30076] = 25'b01110101_01111010_11101111_0;
      patterns[30077] = 25'b01110101_01111011_11110000_0;
      patterns[30078] = 25'b01110101_01111100_11110001_0;
      patterns[30079] = 25'b01110101_01111101_11110010_0;
      patterns[30080] = 25'b01110101_01111110_11110011_0;
      patterns[30081] = 25'b01110101_01111111_11110100_0;
      patterns[30082] = 25'b01110101_10000000_11110101_0;
      patterns[30083] = 25'b01110101_10000001_11110110_0;
      patterns[30084] = 25'b01110101_10000010_11110111_0;
      patterns[30085] = 25'b01110101_10000011_11111000_0;
      patterns[30086] = 25'b01110101_10000100_11111001_0;
      patterns[30087] = 25'b01110101_10000101_11111010_0;
      patterns[30088] = 25'b01110101_10000110_11111011_0;
      patterns[30089] = 25'b01110101_10000111_11111100_0;
      patterns[30090] = 25'b01110101_10001000_11111101_0;
      patterns[30091] = 25'b01110101_10001001_11111110_0;
      patterns[30092] = 25'b01110101_10001010_11111111_0;
      patterns[30093] = 25'b01110101_10001011_00000000_1;
      patterns[30094] = 25'b01110101_10001100_00000001_1;
      patterns[30095] = 25'b01110101_10001101_00000010_1;
      patterns[30096] = 25'b01110101_10001110_00000011_1;
      patterns[30097] = 25'b01110101_10001111_00000100_1;
      patterns[30098] = 25'b01110101_10010000_00000101_1;
      patterns[30099] = 25'b01110101_10010001_00000110_1;
      patterns[30100] = 25'b01110101_10010010_00000111_1;
      patterns[30101] = 25'b01110101_10010011_00001000_1;
      patterns[30102] = 25'b01110101_10010100_00001001_1;
      patterns[30103] = 25'b01110101_10010101_00001010_1;
      patterns[30104] = 25'b01110101_10010110_00001011_1;
      patterns[30105] = 25'b01110101_10010111_00001100_1;
      patterns[30106] = 25'b01110101_10011000_00001101_1;
      patterns[30107] = 25'b01110101_10011001_00001110_1;
      patterns[30108] = 25'b01110101_10011010_00001111_1;
      patterns[30109] = 25'b01110101_10011011_00010000_1;
      patterns[30110] = 25'b01110101_10011100_00010001_1;
      patterns[30111] = 25'b01110101_10011101_00010010_1;
      patterns[30112] = 25'b01110101_10011110_00010011_1;
      patterns[30113] = 25'b01110101_10011111_00010100_1;
      patterns[30114] = 25'b01110101_10100000_00010101_1;
      patterns[30115] = 25'b01110101_10100001_00010110_1;
      patterns[30116] = 25'b01110101_10100010_00010111_1;
      patterns[30117] = 25'b01110101_10100011_00011000_1;
      patterns[30118] = 25'b01110101_10100100_00011001_1;
      patterns[30119] = 25'b01110101_10100101_00011010_1;
      patterns[30120] = 25'b01110101_10100110_00011011_1;
      patterns[30121] = 25'b01110101_10100111_00011100_1;
      patterns[30122] = 25'b01110101_10101000_00011101_1;
      patterns[30123] = 25'b01110101_10101001_00011110_1;
      patterns[30124] = 25'b01110101_10101010_00011111_1;
      patterns[30125] = 25'b01110101_10101011_00100000_1;
      patterns[30126] = 25'b01110101_10101100_00100001_1;
      patterns[30127] = 25'b01110101_10101101_00100010_1;
      patterns[30128] = 25'b01110101_10101110_00100011_1;
      patterns[30129] = 25'b01110101_10101111_00100100_1;
      patterns[30130] = 25'b01110101_10110000_00100101_1;
      patterns[30131] = 25'b01110101_10110001_00100110_1;
      patterns[30132] = 25'b01110101_10110010_00100111_1;
      patterns[30133] = 25'b01110101_10110011_00101000_1;
      patterns[30134] = 25'b01110101_10110100_00101001_1;
      patterns[30135] = 25'b01110101_10110101_00101010_1;
      patterns[30136] = 25'b01110101_10110110_00101011_1;
      patterns[30137] = 25'b01110101_10110111_00101100_1;
      patterns[30138] = 25'b01110101_10111000_00101101_1;
      patterns[30139] = 25'b01110101_10111001_00101110_1;
      patterns[30140] = 25'b01110101_10111010_00101111_1;
      patterns[30141] = 25'b01110101_10111011_00110000_1;
      patterns[30142] = 25'b01110101_10111100_00110001_1;
      patterns[30143] = 25'b01110101_10111101_00110010_1;
      patterns[30144] = 25'b01110101_10111110_00110011_1;
      patterns[30145] = 25'b01110101_10111111_00110100_1;
      patterns[30146] = 25'b01110101_11000000_00110101_1;
      patterns[30147] = 25'b01110101_11000001_00110110_1;
      patterns[30148] = 25'b01110101_11000010_00110111_1;
      patterns[30149] = 25'b01110101_11000011_00111000_1;
      patterns[30150] = 25'b01110101_11000100_00111001_1;
      patterns[30151] = 25'b01110101_11000101_00111010_1;
      patterns[30152] = 25'b01110101_11000110_00111011_1;
      patterns[30153] = 25'b01110101_11000111_00111100_1;
      patterns[30154] = 25'b01110101_11001000_00111101_1;
      patterns[30155] = 25'b01110101_11001001_00111110_1;
      patterns[30156] = 25'b01110101_11001010_00111111_1;
      patterns[30157] = 25'b01110101_11001011_01000000_1;
      patterns[30158] = 25'b01110101_11001100_01000001_1;
      patterns[30159] = 25'b01110101_11001101_01000010_1;
      patterns[30160] = 25'b01110101_11001110_01000011_1;
      patterns[30161] = 25'b01110101_11001111_01000100_1;
      patterns[30162] = 25'b01110101_11010000_01000101_1;
      patterns[30163] = 25'b01110101_11010001_01000110_1;
      patterns[30164] = 25'b01110101_11010010_01000111_1;
      patterns[30165] = 25'b01110101_11010011_01001000_1;
      patterns[30166] = 25'b01110101_11010100_01001001_1;
      patterns[30167] = 25'b01110101_11010101_01001010_1;
      patterns[30168] = 25'b01110101_11010110_01001011_1;
      patterns[30169] = 25'b01110101_11010111_01001100_1;
      patterns[30170] = 25'b01110101_11011000_01001101_1;
      patterns[30171] = 25'b01110101_11011001_01001110_1;
      patterns[30172] = 25'b01110101_11011010_01001111_1;
      patterns[30173] = 25'b01110101_11011011_01010000_1;
      patterns[30174] = 25'b01110101_11011100_01010001_1;
      patterns[30175] = 25'b01110101_11011101_01010010_1;
      patterns[30176] = 25'b01110101_11011110_01010011_1;
      patterns[30177] = 25'b01110101_11011111_01010100_1;
      patterns[30178] = 25'b01110101_11100000_01010101_1;
      patterns[30179] = 25'b01110101_11100001_01010110_1;
      patterns[30180] = 25'b01110101_11100010_01010111_1;
      patterns[30181] = 25'b01110101_11100011_01011000_1;
      patterns[30182] = 25'b01110101_11100100_01011001_1;
      patterns[30183] = 25'b01110101_11100101_01011010_1;
      patterns[30184] = 25'b01110101_11100110_01011011_1;
      patterns[30185] = 25'b01110101_11100111_01011100_1;
      patterns[30186] = 25'b01110101_11101000_01011101_1;
      patterns[30187] = 25'b01110101_11101001_01011110_1;
      patterns[30188] = 25'b01110101_11101010_01011111_1;
      patterns[30189] = 25'b01110101_11101011_01100000_1;
      patterns[30190] = 25'b01110101_11101100_01100001_1;
      patterns[30191] = 25'b01110101_11101101_01100010_1;
      patterns[30192] = 25'b01110101_11101110_01100011_1;
      patterns[30193] = 25'b01110101_11101111_01100100_1;
      patterns[30194] = 25'b01110101_11110000_01100101_1;
      patterns[30195] = 25'b01110101_11110001_01100110_1;
      patterns[30196] = 25'b01110101_11110010_01100111_1;
      patterns[30197] = 25'b01110101_11110011_01101000_1;
      patterns[30198] = 25'b01110101_11110100_01101001_1;
      patterns[30199] = 25'b01110101_11110101_01101010_1;
      patterns[30200] = 25'b01110101_11110110_01101011_1;
      patterns[30201] = 25'b01110101_11110111_01101100_1;
      patterns[30202] = 25'b01110101_11111000_01101101_1;
      patterns[30203] = 25'b01110101_11111001_01101110_1;
      patterns[30204] = 25'b01110101_11111010_01101111_1;
      patterns[30205] = 25'b01110101_11111011_01110000_1;
      patterns[30206] = 25'b01110101_11111100_01110001_1;
      patterns[30207] = 25'b01110101_11111101_01110010_1;
      patterns[30208] = 25'b01110101_11111110_01110011_1;
      patterns[30209] = 25'b01110101_11111111_01110100_1;
      patterns[30210] = 25'b01110110_00000000_01110110_0;
      patterns[30211] = 25'b01110110_00000001_01110111_0;
      patterns[30212] = 25'b01110110_00000010_01111000_0;
      patterns[30213] = 25'b01110110_00000011_01111001_0;
      patterns[30214] = 25'b01110110_00000100_01111010_0;
      patterns[30215] = 25'b01110110_00000101_01111011_0;
      patterns[30216] = 25'b01110110_00000110_01111100_0;
      patterns[30217] = 25'b01110110_00000111_01111101_0;
      patterns[30218] = 25'b01110110_00001000_01111110_0;
      patterns[30219] = 25'b01110110_00001001_01111111_0;
      patterns[30220] = 25'b01110110_00001010_10000000_0;
      patterns[30221] = 25'b01110110_00001011_10000001_0;
      patterns[30222] = 25'b01110110_00001100_10000010_0;
      patterns[30223] = 25'b01110110_00001101_10000011_0;
      patterns[30224] = 25'b01110110_00001110_10000100_0;
      patterns[30225] = 25'b01110110_00001111_10000101_0;
      patterns[30226] = 25'b01110110_00010000_10000110_0;
      patterns[30227] = 25'b01110110_00010001_10000111_0;
      patterns[30228] = 25'b01110110_00010010_10001000_0;
      patterns[30229] = 25'b01110110_00010011_10001001_0;
      patterns[30230] = 25'b01110110_00010100_10001010_0;
      patterns[30231] = 25'b01110110_00010101_10001011_0;
      patterns[30232] = 25'b01110110_00010110_10001100_0;
      patterns[30233] = 25'b01110110_00010111_10001101_0;
      patterns[30234] = 25'b01110110_00011000_10001110_0;
      patterns[30235] = 25'b01110110_00011001_10001111_0;
      patterns[30236] = 25'b01110110_00011010_10010000_0;
      patterns[30237] = 25'b01110110_00011011_10010001_0;
      patterns[30238] = 25'b01110110_00011100_10010010_0;
      patterns[30239] = 25'b01110110_00011101_10010011_0;
      patterns[30240] = 25'b01110110_00011110_10010100_0;
      patterns[30241] = 25'b01110110_00011111_10010101_0;
      patterns[30242] = 25'b01110110_00100000_10010110_0;
      patterns[30243] = 25'b01110110_00100001_10010111_0;
      patterns[30244] = 25'b01110110_00100010_10011000_0;
      patterns[30245] = 25'b01110110_00100011_10011001_0;
      patterns[30246] = 25'b01110110_00100100_10011010_0;
      patterns[30247] = 25'b01110110_00100101_10011011_0;
      patterns[30248] = 25'b01110110_00100110_10011100_0;
      patterns[30249] = 25'b01110110_00100111_10011101_0;
      patterns[30250] = 25'b01110110_00101000_10011110_0;
      patterns[30251] = 25'b01110110_00101001_10011111_0;
      patterns[30252] = 25'b01110110_00101010_10100000_0;
      patterns[30253] = 25'b01110110_00101011_10100001_0;
      patterns[30254] = 25'b01110110_00101100_10100010_0;
      patterns[30255] = 25'b01110110_00101101_10100011_0;
      patterns[30256] = 25'b01110110_00101110_10100100_0;
      patterns[30257] = 25'b01110110_00101111_10100101_0;
      patterns[30258] = 25'b01110110_00110000_10100110_0;
      patterns[30259] = 25'b01110110_00110001_10100111_0;
      patterns[30260] = 25'b01110110_00110010_10101000_0;
      patterns[30261] = 25'b01110110_00110011_10101001_0;
      patterns[30262] = 25'b01110110_00110100_10101010_0;
      patterns[30263] = 25'b01110110_00110101_10101011_0;
      patterns[30264] = 25'b01110110_00110110_10101100_0;
      patterns[30265] = 25'b01110110_00110111_10101101_0;
      patterns[30266] = 25'b01110110_00111000_10101110_0;
      patterns[30267] = 25'b01110110_00111001_10101111_0;
      patterns[30268] = 25'b01110110_00111010_10110000_0;
      patterns[30269] = 25'b01110110_00111011_10110001_0;
      patterns[30270] = 25'b01110110_00111100_10110010_0;
      patterns[30271] = 25'b01110110_00111101_10110011_0;
      patterns[30272] = 25'b01110110_00111110_10110100_0;
      patterns[30273] = 25'b01110110_00111111_10110101_0;
      patterns[30274] = 25'b01110110_01000000_10110110_0;
      patterns[30275] = 25'b01110110_01000001_10110111_0;
      patterns[30276] = 25'b01110110_01000010_10111000_0;
      patterns[30277] = 25'b01110110_01000011_10111001_0;
      patterns[30278] = 25'b01110110_01000100_10111010_0;
      patterns[30279] = 25'b01110110_01000101_10111011_0;
      patterns[30280] = 25'b01110110_01000110_10111100_0;
      patterns[30281] = 25'b01110110_01000111_10111101_0;
      patterns[30282] = 25'b01110110_01001000_10111110_0;
      patterns[30283] = 25'b01110110_01001001_10111111_0;
      patterns[30284] = 25'b01110110_01001010_11000000_0;
      patterns[30285] = 25'b01110110_01001011_11000001_0;
      patterns[30286] = 25'b01110110_01001100_11000010_0;
      patterns[30287] = 25'b01110110_01001101_11000011_0;
      patterns[30288] = 25'b01110110_01001110_11000100_0;
      patterns[30289] = 25'b01110110_01001111_11000101_0;
      patterns[30290] = 25'b01110110_01010000_11000110_0;
      patterns[30291] = 25'b01110110_01010001_11000111_0;
      patterns[30292] = 25'b01110110_01010010_11001000_0;
      patterns[30293] = 25'b01110110_01010011_11001001_0;
      patterns[30294] = 25'b01110110_01010100_11001010_0;
      patterns[30295] = 25'b01110110_01010101_11001011_0;
      patterns[30296] = 25'b01110110_01010110_11001100_0;
      patterns[30297] = 25'b01110110_01010111_11001101_0;
      patterns[30298] = 25'b01110110_01011000_11001110_0;
      patterns[30299] = 25'b01110110_01011001_11001111_0;
      patterns[30300] = 25'b01110110_01011010_11010000_0;
      patterns[30301] = 25'b01110110_01011011_11010001_0;
      patterns[30302] = 25'b01110110_01011100_11010010_0;
      patterns[30303] = 25'b01110110_01011101_11010011_0;
      patterns[30304] = 25'b01110110_01011110_11010100_0;
      patterns[30305] = 25'b01110110_01011111_11010101_0;
      patterns[30306] = 25'b01110110_01100000_11010110_0;
      patterns[30307] = 25'b01110110_01100001_11010111_0;
      patterns[30308] = 25'b01110110_01100010_11011000_0;
      patterns[30309] = 25'b01110110_01100011_11011001_0;
      patterns[30310] = 25'b01110110_01100100_11011010_0;
      patterns[30311] = 25'b01110110_01100101_11011011_0;
      patterns[30312] = 25'b01110110_01100110_11011100_0;
      patterns[30313] = 25'b01110110_01100111_11011101_0;
      patterns[30314] = 25'b01110110_01101000_11011110_0;
      patterns[30315] = 25'b01110110_01101001_11011111_0;
      patterns[30316] = 25'b01110110_01101010_11100000_0;
      patterns[30317] = 25'b01110110_01101011_11100001_0;
      patterns[30318] = 25'b01110110_01101100_11100010_0;
      patterns[30319] = 25'b01110110_01101101_11100011_0;
      patterns[30320] = 25'b01110110_01101110_11100100_0;
      patterns[30321] = 25'b01110110_01101111_11100101_0;
      patterns[30322] = 25'b01110110_01110000_11100110_0;
      patterns[30323] = 25'b01110110_01110001_11100111_0;
      patterns[30324] = 25'b01110110_01110010_11101000_0;
      patterns[30325] = 25'b01110110_01110011_11101001_0;
      patterns[30326] = 25'b01110110_01110100_11101010_0;
      patterns[30327] = 25'b01110110_01110101_11101011_0;
      patterns[30328] = 25'b01110110_01110110_11101100_0;
      patterns[30329] = 25'b01110110_01110111_11101101_0;
      patterns[30330] = 25'b01110110_01111000_11101110_0;
      patterns[30331] = 25'b01110110_01111001_11101111_0;
      patterns[30332] = 25'b01110110_01111010_11110000_0;
      patterns[30333] = 25'b01110110_01111011_11110001_0;
      patterns[30334] = 25'b01110110_01111100_11110010_0;
      patterns[30335] = 25'b01110110_01111101_11110011_0;
      patterns[30336] = 25'b01110110_01111110_11110100_0;
      patterns[30337] = 25'b01110110_01111111_11110101_0;
      patterns[30338] = 25'b01110110_10000000_11110110_0;
      patterns[30339] = 25'b01110110_10000001_11110111_0;
      patterns[30340] = 25'b01110110_10000010_11111000_0;
      patterns[30341] = 25'b01110110_10000011_11111001_0;
      patterns[30342] = 25'b01110110_10000100_11111010_0;
      patterns[30343] = 25'b01110110_10000101_11111011_0;
      patterns[30344] = 25'b01110110_10000110_11111100_0;
      patterns[30345] = 25'b01110110_10000111_11111101_0;
      patterns[30346] = 25'b01110110_10001000_11111110_0;
      patterns[30347] = 25'b01110110_10001001_11111111_0;
      patterns[30348] = 25'b01110110_10001010_00000000_1;
      patterns[30349] = 25'b01110110_10001011_00000001_1;
      patterns[30350] = 25'b01110110_10001100_00000010_1;
      patterns[30351] = 25'b01110110_10001101_00000011_1;
      patterns[30352] = 25'b01110110_10001110_00000100_1;
      patterns[30353] = 25'b01110110_10001111_00000101_1;
      patterns[30354] = 25'b01110110_10010000_00000110_1;
      patterns[30355] = 25'b01110110_10010001_00000111_1;
      patterns[30356] = 25'b01110110_10010010_00001000_1;
      patterns[30357] = 25'b01110110_10010011_00001001_1;
      patterns[30358] = 25'b01110110_10010100_00001010_1;
      patterns[30359] = 25'b01110110_10010101_00001011_1;
      patterns[30360] = 25'b01110110_10010110_00001100_1;
      patterns[30361] = 25'b01110110_10010111_00001101_1;
      patterns[30362] = 25'b01110110_10011000_00001110_1;
      patterns[30363] = 25'b01110110_10011001_00001111_1;
      patterns[30364] = 25'b01110110_10011010_00010000_1;
      patterns[30365] = 25'b01110110_10011011_00010001_1;
      patterns[30366] = 25'b01110110_10011100_00010010_1;
      patterns[30367] = 25'b01110110_10011101_00010011_1;
      patterns[30368] = 25'b01110110_10011110_00010100_1;
      patterns[30369] = 25'b01110110_10011111_00010101_1;
      patterns[30370] = 25'b01110110_10100000_00010110_1;
      patterns[30371] = 25'b01110110_10100001_00010111_1;
      patterns[30372] = 25'b01110110_10100010_00011000_1;
      patterns[30373] = 25'b01110110_10100011_00011001_1;
      patterns[30374] = 25'b01110110_10100100_00011010_1;
      patterns[30375] = 25'b01110110_10100101_00011011_1;
      patterns[30376] = 25'b01110110_10100110_00011100_1;
      patterns[30377] = 25'b01110110_10100111_00011101_1;
      patterns[30378] = 25'b01110110_10101000_00011110_1;
      patterns[30379] = 25'b01110110_10101001_00011111_1;
      patterns[30380] = 25'b01110110_10101010_00100000_1;
      patterns[30381] = 25'b01110110_10101011_00100001_1;
      patterns[30382] = 25'b01110110_10101100_00100010_1;
      patterns[30383] = 25'b01110110_10101101_00100011_1;
      patterns[30384] = 25'b01110110_10101110_00100100_1;
      patterns[30385] = 25'b01110110_10101111_00100101_1;
      patterns[30386] = 25'b01110110_10110000_00100110_1;
      patterns[30387] = 25'b01110110_10110001_00100111_1;
      patterns[30388] = 25'b01110110_10110010_00101000_1;
      patterns[30389] = 25'b01110110_10110011_00101001_1;
      patterns[30390] = 25'b01110110_10110100_00101010_1;
      patterns[30391] = 25'b01110110_10110101_00101011_1;
      patterns[30392] = 25'b01110110_10110110_00101100_1;
      patterns[30393] = 25'b01110110_10110111_00101101_1;
      patterns[30394] = 25'b01110110_10111000_00101110_1;
      patterns[30395] = 25'b01110110_10111001_00101111_1;
      patterns[30396] = 25'b01110110_10111010_00110000_1;
      patterns[30397] = 25'b01110110_10111011_00110001_1;
      patterns[30398] = 25'b01110110_10111100_00110010_1;
      patterns[30399] = 25'b01110110_10111101_00110011_1;
      patterns[30400] = 25'b01110110_10111110_00110100_1;
      patterns[30401] = 25'b01110110_10111111_00110101_1;
      patterns[30402] = 25'b01110110_11000000_00110110_1;
      patterns[30403] = 25'b01110110_11000001_00110111_1;
      patterns[30404] = 25'b01110110_11000010_00111000_1;
      patterns[30405] = 25'b01110110_11000011_00111001_1;
      patterns[30406] = 25'b01110110_11000100_00111010_1;
      patterns[30407] = 25'b01110110_11000101_00111011_1;
      patterns[30408] = 25'b01110110_11000110_00111100_1;
      patterns[30409] = 25'b01110110_11000111_00111101_1;
      patterns[30410] = 25'b01110110_11001000_00111110_1;
      patterns[30411] = 25'b01110110_11001001_00111111_1;
      patterns[30412] = 25'b01110110_11001010_01000000_1;
      patterns[30413] = 25'b01110110_11001011_01000001_1;
      patterns[30414] = 25'b01110110_11001100_01000010_1;
      patterns[30415] = 25'b01110110_11001101_01000011_1;
      patterns[30416] = 25'b01110110_11001110_01000100_1;
      patterns[30417] = 25'b01110110_11001111_01000101_1;
      patterns[30418] = 25'b01110110_11010000_01000110_1;
      patterns[30419] = 25'b01110110_11010001_01000111_1;
      patterns[30420] = 25'b01110110_11010010_01001000_1;
      patterns[30421] = 25'b01110110_11010011_01001001_1;
      patterns[30422] = 25'b01110110_11010100_01001010_1;
      patterns[30423] = 25'b01110110_11010101_01001011_1;
      patterns[30424] = 25'b01110110_11010110_01001100_1;
      patterns[30425] = 25'b01110110_11010111_01001101_1;
      patterns[30426] = 25'b01110110_11011000_01001110_1;
      patterns[30427] = 25'b01110110_11011001_01001111_1;
      patterns[30428] = 25'b01110110_11011010_01010000_1;
      patterns[30429] = 25'b01110110_11011011_01010001_1;
      patterns[30430] = 25'b01110110_11011100_01010010_1;
      patterns[30431] = 25'b01110110_11011101_01010011_1;
      patterns[30432] = 25'b01110110_11011110_01010100_1;
      patterns[30433] = 25'b01110110_11011111_01010101_1;
      patterns[30434] = 25'b01110110_11100000_01010110_1;
      patterns[30435] = 25'b01110110_11100001_01010111_1;
      patterns[30436] = 25'b01110110_11100010_01011000_1;
      patterns[30437] = 25'b01110110_11100011_01011001_1;
      patterns[30438] = 25'b01110110_11100100_01011010_1;
      patterns[30439] = 25'b01110110_11100101_01011011_1;
      patterns[30440] = 25'b01110110_11100110_01011100_1;
      patterns[30441] = 25'b01110110_11100111_01011101_1;
      patterns[30442] = 25'b01110110_11101000_01011110_1;
      patterns[30443] = 25'b01110110_11101001_01011111_1;
      patterns[30444] = 25'b01110110_11101010_01100000_1;
      patterns[30445] = 25'b01110110_11101011_01100001_1;
      patterns[30446] = 25'b01110110_11101100_01100010_1;
      patterns[30447] = 25'b01110110_11101101_01100011_1;
      patterns[30448] = 25'b01110110_11101110_01100100_1;
      patterns[30449] = 25'b01110110_11101111_01100101_1;
      patterns[30450] = 25'b01110110_11110000_01100110_1;
      patterns[30451] = 25'b01110110_11110001_01100111_1;
      patterns[30452] = 25'b01110110_11110010_01101000_1;
      patterns[30453] = 25'b01110110_11110011_01101001_1;
      patterns[30454] = 25'b01110110_11110100_01101010_1;
      patterns[30455] = 25'b01110110_11110101_01101011_1;
      patterns[30456] = 25'b01110110_11110110_01101100_1;
      patterns[30457] = 25'b01110110_11110111_01101101_1;
      patterns[30458] = 25'b01110110_11111000_01101110_1;
      patterns[30459] = 25'b01110110_11111001_01101111_1;
      patterns[30460] = 25'b01110110_11111010_01110000_1;
      patterns[30461] = 25'b01110110_11111011_01110001_1;
      patterns[30462] = 25'b01110110_11111100_01110010_1;
      patterns[30463] = 25'b01110110_11111101_01110011_1;
      patterns[30464] = 25'b01110110_11111110_01110100_1;
      patterns[30465] = 25'b01110110_11111111_01110101_1;
      patterns[30466] = 25'b01110111_00000000_01110111_0;
      patterns[30467] = 25'b01110111_00000001_01111000_0;
      patterns[30468] = 25'b01110111_00000010_01111001_0;
      patterns[30469] = 25'b01110111_00000011_01111010_0;
      patterns[30470] = 25'b01110111_00000100_01111011_0;
      patterns[30471] = 25'b01110111_00000101_01111100_0;
      patterns[30472] = 25'b01110111_00000110_01111101_0;
      patterns[30473] = 25'b01110111_00000111_01111110_0;
      patterns[30474] = 25'b01110111_00001000_01111111_0;
      patterns[30475] = 25'b01110111_00001001_10000000_0;
      patterns[30476] = 25'b01110111_00001010_10000001_0;
      patterns[30477] = 25'b01110111_00001011_10000010_0;
      patterns[30478] = 25'b01110111_00001100_10000011_0;
      patterns[30479] = 25'b01110111_00001101_10000100_0;
      patterns[30480] = 25'b01110111_00001110_10000101_0;
      patterns[30481] = 25'b01110111_00001111_10000110_0;
      patterns[30482] = 25'b01110111_00010000_10000111_0;
      patterns[30483] = 25'b01110111_00010001_10001000_0;
      patterns[30484] = 25'b01110111_00010010_10001001_0;
      patterns[30485] = 25'b01110111_00010011_10001010_0;
      patterns[30486] = 25'b01110111_00010100_10001011_0;
      patterns[30487] = 25'b01110111_00010101_10001100_0;
      patterns[30488] = 25'b01110111_00010110_10001101_0;
      patterns[30489] = 25'b01110111_00010111_10001110_0;
      patterns[30490] = 25'b01110111_00011000_10001111_0;
      patterns[30491] = 25'b01110111_00011001_10010000_0;
      patterns[30492] = 25'b01110111_00011010_10010001_0;
      patterns[30493] = 25'b01110111_00011011_10010010_0;
      patterns[30494] = 25'b01110111_00011100_10010011_0;
      patterns[30495] = 25'b01110111_00011101_10010100_0;
      patterns[30496] = 25'b01110111_00011110_10010101_0;
      patterns[30497] = 25'b01110111_00011111_10010110_0;
      patterns[30498] = 25'b01110111_00100000_10010111_0;
      patterns[30499] = 25'b01110111_00100001_10011000_0;
      patterns[30500] = 25'b01110111_00100010_10011001_0;
      patterns[30501] = 25'b01110111_00100011_10011010_0;
      patterns[30502] = 25'b01110111_00100100_10011011_0;
      patterns[30503] = 25'b01110111_00100101_10011100_0;
      patterns[30504] = 25'b01110111_00100110_10011101_0;
      patterns[30505] = 25'b01110111_00100111_10011110_0;
      patterns[30506] = 25'b01110111_00101000_10011111_0;
      patterns[30507] = 25'b01110111_00101001_10100000_0;
      patterns[30508] = 25'b01110111_00101010_10100001_0;
      patterns[30509] = 25'b01110111_00101011_10100010_0;
      patterns[30510] = 25'b01110111_00101100_10100011_0;
      patterns[30511] = 25'b01110111_00101101_10100100_0;
      patterns[30512] = 25'b01110111_00101110_10100101_0;
      patterns[30513] = 25'b01110111_00101111_10100110_0;
      patterns[30514] = 25'b01110111_00110000_10100111_0;
      patterns[30515] = 25'b01110111_00110001_10101000_0;
      patterns[30516] = 25'b01110111_00110010_10101001_0;
      patterns[30517] = 25'b01110111_00110011_10101010_0;
      patterns[30518] = 25'b01110111_00110100_10101011_0;
      patterns[30519] = 25'b01110111_00110101_10101100_0;
      patterns[30520] = 25'b01110111_00110110_10101101_0;
      patterns[30521] = 25'b01110111_00110111_10101110_0;
      patterns[30522] = 25'b01110111_00111000_10101111_0;
      patterns[30523] = 25'b01110111_00111001_10110000_0;
      patterns[30524] = 25'b01110111_00111010_10110001_0;
      patterns[30525] = 25'b01110111_00111011_10110010_0;
      patterns[30526] = 25'b01110111_00111100_10110011_0;
      patterns[30527] = 25'b01110111_00111101_10110100_0;
      patterns[30528] = 25'b01110111_00111110_10110101_0;
      patterns[30529] = 25'b01110111_00111111_10110110_0;
      patterns[30530] = 25'b01110111_01000000_10110111_0;
      patterns[30531] = 25'b01110111_01000001_10111000_0;
      patterns[30532] = 25'b01110111_01000010_10111001_0;
      patterns[30533] = 25'b01110111_01000011_10111010_0;
      patterns[30534] = 25'b01110111_01000100_10111011_0;
      patterns[30535] = 25'b01110111_01000101_10111100_0;
      patterns[30536] = 25'b01110111_01000110_10111101_0;
      patterns[30537] = 25'b01110111_01000111_10111110_0;
      patterns[30538] = 25'b01110111_01001000_10111111_0;
      patterns[30539] = 25'b01110111_01001001_11000000_0;
      patterns[30540] = 25'b01110111_01001010_11000001_0;
      patterns[30541] = 25'b01110111_01001011_11000010_0;
      patterns[30542] = 25'b01110111_01001100_11000011_0;
      patterns[30543] = 25'b01110111_01001101_11000100_0;
      patterns[30544] = 25'b01110111_01001110_11000101_0;
      patterns[30545] = 25'b01110111_01001111_11000110_0;
      patterns[30546] = 25'b01110111_01010000_11000111_0;
      patterns[30547] = 25'b01110111_01010001_11001000_0;
      patterns[30548] = 25'b01110111_01010010_11001001_0;
      patterns[30549] = 25'b01110111_01010011_11001010_0;
      patterns[30550] = 25'b01110111_01010100_11001011_0;
      patterns[30551] = 25'b01110111_01010101_11001100_0;
      patterns[30552] = 25'b01110111_01010110_11001101_0;
      patterns[30553] = 25'b01110111_01010111_11001110_0;
      patterns[30554] = 25'b01110111_01011000_11001111_0;
      patterns[30555] = 25'b01110111_01011001_11010000_0;
      patterns[30556] = 25'b01110111_01011010_11010001_0;
      patterns[30557] = 25'b01110111_01011011_11010010_0;
      patterns[30558] = 25'b01110111_01011100_11010011_0;
      patterns[30559] = 25'b01110111_01011101_11010100_0;
      patterns[30560] = 25'b01110111_01011110_11010101_0;
      patterns[30561] = 25'b01110111_01011111_11010110_0;
      patterns[30562] = 25'b01110111_01100000_11010111_0;
      patterns[30563] = 25'b01110111_01100001_11011000_0;
      patterns[30564] = 25'b01110111_01100010_11011001_0;
      patterns[30565] = 25'b01110111_01100011_11011010_0;
      patterns[30566] = 25'b01110111_01100100_11011011_0;
      patterns[30567] = 25'b01110111_01100101_11011100_0;
      patterns[30568] = 25'b01110111_01100110_11011101_0;
      patterns[30569] = 25'b01110111_01100111_11011110_0;
      patterns[30570] = 25'b01110111_01101000_11011111_0;
      patterns[30571] = 25'b01110111_01101001_11100000_0;
      patterns[30572] = 25'b01110111_01101010_11100001_0;
      patterns[30573] = 25'b01110111_01101011_11100010_0;
      patterns[30574] = 25'b01110111_01101100_11100011_0;
      patterns[30575] = 25'b01110111_01101101_11100100_0;
      patterns[30576] = 25'b01110111_01101110_11100101_0;
      patterns[30577] = 25'b01110111_01101111_11100110_0;
      patterns[30578] = 25'b01110111_01110000_11100111_0;
      patterns[30579] = 25'b01110111_01110001_11101000_0;
      patterns[30580] = 25'b01110111_01110010_11101001_0;
      patterns[30581] = 25'b01110111_01110011_11101010_0;
      patterns[30582] = 25'b01110111_01110100_11101011_0;
      patterns[30583] = 25'b01110111_01110101_11101100_0;
      patterns[30584] = 25'b01110111_01110110_11101101_0;
      patterns[30585] = 25'b01110111_01110111_11101110_0;
      patterns[30586] = 25'b01110111_01111000_11101111_0;
      patterns[30587] = 25'b01110111_01111001_11110000_0;
      patterns[30588] = 25'b01110111_01111010_11110001_0;
      patterns[30589] = 25'b01110111_01111011_11110010_0;
      patterns[30590] = 25'b01110111_01111100_11110011_0;
      patterns[30591] = 25'b01110111_01111101_11110100_0;
      patterns[30592] = 25'b01110111_01111110_11110101_0;
      patterns[30593] = 25'b01110111_01111111_11110110_0;
      patterns[30594] = 25'b01110111_10000000_11110111_0;
      patterns[30595] = 25'b01110111_10000001_11111000_0;
      patterns[30596] = 25'b01110111_10000010_11111001_0;
      patterns[30597] = 25'b01110111_10000011_11111010_0;
      patterns[30598] = 25'b01110111_10000100_11111011_0;
      patterns[30599] = 25'b01110111_10000101_11111100_0;
      patterns[30600] = 25'b01110111_10000110_11111101_0;
      patterns[30601] = 25'b01110111_10000111_11111110_0;
      patterns[30602] = 25'b01110111_10001000_11111111_0;
      patterns[30603] = 25'b01110111_10001001_00000000_1;
      patterns[30604] = 25'b01110111_10001010_00000001_1;
      patterns[30605] = 25'b01110111_10001011_00000010_1;
      patterns[30606] = 25'b01110111_10001100_00000011_1;
      patterns[30607] = 25'b01110111_10001101_00000100_1;
      patterns[30608] = 25'b01110111_10001110_00000101_1;
      patterns[30609] = 25'b01110111_10001111_00000110_1;
      patterns[30610] = 25'b01110111_10010000_00000111_1;
      patterns[30611] = 25'b01110111_10010001_00001000_1;
      patterns[30612] = 25'b01110111_10010010_00001001_1;
      patterns[30613] = 25'b01110111_10010011_00001010_1;
      patterns[30614] = 25'b01110111_10010100_00001011_1;
      patterns[30615] = 25'b01110111_10010101_00001100_1;
      patterns[30616] = 25'b01110111_10010110_00001101_1;
      patterns[30617] = 25'b01110111_10010111_00001110_1;
      patterns[30618] = 25'b01110111_10011000_00001111_1;
      patterns[30619] = 25'b01110111_10011001_00010000_1;
      patterns[30620] = 25'b01110111_10011010_00010001_1;
      patterns[30621] = 25'b01110111_10011011_00010010_1;
      patterns[30622] = 25'b01110111_10011100_00010011_1;
      patterns[30623] = 25'b01110111_10011101_00010100_1;
      patterns[30624] = 25'b01110111_10011110_00010101_1;
      patterns[30625] = 25'b01110111_10011111_00010110_1;
      patterns[30626] = 25'b01110111_10100000_00010111_1;
      patterns[30627] = 25'b01110111_10100001_00011000_1;
      patterns[30628] = 25'b01110111_10100010_00011001_1;
      patterns[30629] = 25'b01110111_10100011_00011010_1;
      patterns[30630] = 25'b01110111_10100100_00011011_1;
      patterns[30631] = 25'b01110111_10100101_00011100_1;
      patterns[30632] = 25'b01110111_10100110_00011101_1;
      patterns[30633] = 25'b01110111_10100111_00011110_1;
      patterns[30634] = 25'b01110111_10101000_00011111_1;
      patterns[30635] = 25'b01110111_10101001_00100000_1;
      patterns[30636] = 25'b01110111_10101010_00100001_1;
      patterns[30637] = 25'b01110111_10101011_00100010_1;
      patterns[30638] = 25'b01110111_10101100_00100011_1;
      patterns[30639] = 25'b01110111_10101101_00100100_1;
      patterns[30640] = 25'b01110111_10101110_00100101_1;
      patterns[30641] = 25'b01110111_10101111_00100110_1;
      patterns[30642] = 25'b01110111_10110000_00100111_1;
      patterns[30643] = 25'b01110111_10110001_00101000_1;
      patterns[30644] = 25'b01110111_10110010_00101001_1;
      patterns[30645] = 25'b01110111_10110011_00101010_1;
      patterns[30646] = 25'b01110111_10110100_00101011_1;
      patterns[30647] = 25'b01110111_10110101_00101100_1;
      patterns[30648] = 25'b01110111_10110110_00101101_1;
      patterns[30649] = 25'b01110111_10110111_00101110_1;
      patterns[30650] = 25'b01110111_10111000_00101111_1;
      patterns[30651] = 25'b01110111_10111001_00110000_1;
      patterns[30652] = 25'b01110111_10111010_00110001_1;
      patterns[30653] = 25'b01110111_10111011_00110010_1;
      patterns[30654] = 25'b01110111_10111100_00110011_1;
      patterns[30655] = 25'b01110111_10111101_00110100_1;
      patterns[30656] = 25'b01110111_10111110_00110101_1;
      patterns[30657] = 25'b01110111_10111111_00110110_1;
      patterns[30658] = 25'b01110111_11000000_00110111_1;
      patterns[30659] = 25'b01110111_11000001_00111000_1;
      patterns[30660] = 25'b01110111_11000010_00111001_1;
      patterns[30661] = 25'b01110111_11000011_00111010_1;
      patterns[30662] = 25'b01110111_11000100_00111011_1;
      patterns[30663] = 25'b01110111_11000101_00111100_1;
      patterns[30664] = 25'b01110111_11000110_00111101_1;
      patterns[30665] = 25'b01110111_11000111_00111110_1;
      patterns[30666] = 25'b01110111_11001000_00111111_1;
      patterns[30667] = 25'b01110111_11001001_01000000_1;
      patterns[30668] = 25'b01110111_11001010_01000001_1;
      patterns[30669] = 25'b01110111_11001011_01000010_1;
      patterns[30670] = 25'b01110111_11001100_01000011_1;
      patterns[30671] = 25'b01110111_11001101_01000100_1;
      patterns[30672] = 25'b01110111_11001110_01000101_1;
      patterns[30673] = 25'b01110111_11001111_01000110_1;
      patterns[30674] = 25'b01110111_11010000_01000111_1;
      patterns[30675] = 25'b01110111_11010001_01001000_1;
      patterns[30676] = 25'b01110111_11010010_01001001_1;
      patterns[30677] = 25'b01110111_11010011_01001010_1;
      patterns[30678] = 25'b01110111_11010100_01001011_1;
      patterns[30679] = 25'b01110111_11010101_01001100_1;
      patterns[30680] = 25'b01110111_11010110_01001101_1;
      patterns[30681] = 25'b01110111_11010111_01001110_1;
      patterns[30682] = 25'b01110111_11011000_01001111_1;
      patterns[30683] = 25'b01110111_11011001_01010000_1;
      patterns[30684] = 25'b01110111_11011010_01010001_1;
      patterns[30685] = 25'b01110111_11011011_01010010_1;
      patterns[30686] = 25'b01110111_11011100_01010011_1;
      patterns[30687] = 25'b01110111_11011101_01010100_1;
      patterns[30688] = 25'b01110111_11011110_01010101_1;
      patterns[30689] = 25'b01110111_11011111_01010110_1;
      patterns[30690] = 25'b01110111_11100000_01010111_1;
      patterns[30691] = 25'b01110111_11100001_01011000_1;
      patterns[30692] = 25'b01110111_11100010_01011001_1;
      patterns[30693] = 25'b01110111_11100011_01011010_1;
      patterns[30694] = 25'b01110111_11100100_01011011_1;
      patterns[30695] = 25'b01110111_11100101_01011100_1;
      patterns[30696] = 25'b01110111_11100110_01011101_1;
      patterns[30697] = 25'b01110111_11100111_01011110_1;
      patterns[30698] = 25'b01110111_11101000_01011111_1;
      patterns[30699] = 25'b01110111_11101001_01100000_1;
      patterns[30700] = 25'b01110111_11101010_01100001_1;
      patterns[30701] = 25'b01110111_11101011_01100010_1;
      patterns[30702] = 25'b01110111_11101100_01100011_1;
      patterns[30703] = 25'b01110111_11101101_01100100_1;
      patterns[30704] = 25'b01110111_11101110_01100101_1;
      patterns[30705] = 25'b01110111_11101111_01100110_1;
      patterns[30706] = 25'b01110111_11110000_01100111_1;
      patterns[30707] = 25'b01110111_11110001_01101000_1;
      patterns[30708] = 25'b01110111_11110010_01101001_1;
      patterns[30709] = 25'b01110111_11110011_01101010_1;
      patterns[30710] = 25'b01110111_11110100_01101011_1;
      patterns[30711] = 25'b01110111_11110101_01101100_1;
      patterns[30712] = 25'b01110111_11110110_01101101_1;
      patterns[30713] = 25'b01110111_11110111_01101110_1;
      patterns[30714] = 25'b01110111_11111000_01101111_1;
      patterns[30715] = 25'b01110111_11111001_01110000_1;
      patterns[30716] = 25'b01110111_11111010_01110001_1;
      patterns[30717] = 25'b01110111_11111011_01110010_1;
      patterns[30718] = 25'b01110111_11111100_01110011_1;
      patterns[30719] = 25'b01110111_11111101_01110100_1;
      patterns[30720] = 25'b01110111_11111110_01110101_1;
      patterns[30721] = 25'b01110111_11111111_01110110_1;
      patterns[30722] = 25'b01111000_00000000_01111000_0;
      patterns[30723] = 25'b01111000_00000001_01111001_0;
      patterns[30724] = 25'b01111000_00000010_01111010_0;
      patterns[30725] = 25'b01111000_00000011_01111011_0;
      patterns[30726] = 25'b01111000_00000100_01111100_0;
      patterns[30727] = 25'b01111000_00000101_01111101_0;
      patterns[30728] = 25'b01111000_00000110_01111110_0;
      patterns[30729] = 25'b01111000_00000111_01111111_0;
      patterns[30730] = 25'b01111000_00001000_10000000_0;
      patterns[30731] = 25'b01111000_00001001_10000001_0;
      patterns[30732] = 25'b01111000_00001010_10000010_0;
      patterns[30733] = 25'b01111000_00001011_10000011_0;
      patterns[30734] = 25'b01111000_00001100_10000100_0;
      patterns[30735] = 25'b01111000_00001101_10000101_0;
      patterns[30736] = 25'b01111000_00001110_10000110_0;
      patterns[30737] = 25'b01111000_00001111_10000111_0;
      patterns[30738] = 25'b01111000_00010000_10001000_0;
      patterns[30739] = 25'b01111000_00010001_10001001_0;
      patterns[30740] = 25'b01111000_00010010_10001010_0;
      patterns[30741] = 25'b01111000_00010011_10001011_0;
      patterns[30742] = 25'b01111000_00010100_10001100_0;
      patterns[30743] = 25'b01111000_00010101_10001101_0;
      patterns[30744] = 25'b01111000_00010110_10001110_0;
      patterns[30745] = 25'b01111000_00010111_10001111_0;
      patterns[30746] = 25'b01111000_00011000_10010000_0;
      patterns[30747] = 25'b01111000_00011001_10010001_0;
      patterns[30748] = 25'b01111000_00011010_10010010_0;
      patterns[30749] = 25'b01111000_00011011_10010011_0;
      patterns[30750] = 25'b01111000_00011100_10010100_0;
      patterns[30751] = 25'b01111000_00011101_10010101_0;
      patterns[30752] = 25'b01111000_00011110_10010110_0;
      patterns[30753] = 25'b01111000_00011111_10010111_0;
      patterns[30754] = 25'b01111000_00100000_10011000_0;
      patterns[30755] = 25'b01111000_00100001_10011001_0;
      patterns[30756] = 25'b01111000_00100010_10011010_0;
      patterns[30757] = 25'b01111000_00100011_10011011_0;
      patterns[30758] = 25'b01111000_00100100_10011100_0;
      patterns[30759] = 25'b01111000_00100101_10011101_0;
      patterns[30760] = 25'b01111000_00100110_10011110_0;
      patterns[30761] = 25'b01111000_00100111_10011111_0;
      patterns[30762] = 25'b01111000_00101000_10100000_0;
      patterns[30763] = 25'b01111000_00101001_10100001_0;
      patterns[30764] = 25'b01111000_00101010_10100010_0;
      patterns[30765] = 25'b01111000_00101011_10100011_0;
      patterns[30766] = 25'b01111000_00101100_10100100_0;
      patterns[30767] = 25'b01111000_00101101_10100101_0;
      patterns[30768] = 25'b01111000_00101110_10100110_0;
      patterns[30769] = 25'b01111000_00101111_10100111_0;
      patterns[30770] = 25'b01111000_00110000_10101000_0;
      patterns[30771] = 25'b01111000_00110001_10101001_0;
      patterns[30772] = 25'b01111000_00110010_10101010_0;
      patterns[30773] = 25'b01111000_00110011_10101011_0;
      patterns[30774] = 25'b01111000_00110100_10101100_0;
      patterns[30775] = 25'b01111000_00110101_10101101_0;
      patterns[30776] = 25'b01111000_00110110_10101110_0;
      patterns[30777] = 25'b01111000_00110111_10101111_0;
      patterns[30778] = 25'b01111000_00111000_10110000_0;
      patterns[30779] = 25'b01111000_00111001_10110001_0;
      patterns[30780] = 25'b01111000_00111010_10110010_0;
      patterns[30781] = 25'b01111000_00111011_10110011_0;
      patterns[30782] = 25'b01111000_00111100_10110100_0;
      patterns[30783] = 25'b01111000_00111101_10110101_0;
      patterns[30784] = 25'b01111000_00111110_10110110_0;
      patterns[30785] = 25'b01111000_00111111_10110111_0;
      patterns[30786] = 25'b01111000_01000000_10111000_0;
      patterns[30787] = 25'b01111000_01000001_10111001_0;
      patterns[30788] = 25'b01111000_01000010_10111010_0;
      patterns[30789] = 25'b01111000_01000011_10111011_0;
      patterns[30790] = 25'b01111000_01000100_10111100_0;
      patterns[30791] = 25'b01111000_01000101_10111101_0;
      patterns[30792] = 25'b01111000_01000110_10111110_0;
      patterns[30793] = 25'b01111000_01000111_10111111_0;
      patterns[30794] = 25'b01111000_01001000_11000000_0;
      patterns[30795] = 25'b01111000_01001001_11000001_0;
      patterns[30796] = 25'b01111000_01001010_11000010_0;
      patterns[30797] = 25'b01111000_01001011_11000011_0;
      patterns[30798] = 25'b01111000_01001100_11000100_0;
      patterns[30799] = 25'b01111000_01001101_11000101_0;
      patterns[30800] = 25'b01111000_01001110_11000110_0;
      patterns[30801] = 25'b01111000_01001111_11000111_0;
      patterns[30802] = 25'b01111000_01010000_11001000_0;
      patterns[30803] = 25'b01111000_01010001_11001001_0;
      patterns[30804] = 25'b01111000_01010010_11001010_0;
      patterns[30805] = 25'b01111000_01010011_11001011_0;
      patterns[30806] = 25'b01111000_01010100_11001100_0;
      patterns[30807] = 25'b01111000_01010101_11001101_0;
      patterns[30808] = 25'b01111000_01010110_11001110_0;
      patterns[30809] = 25'b01111000_01010111_11001111_0;
      patterns[30810] = 25'b01111000_01011000_11010000_0;
      patterns[30811] = 25'b01111000_01011001_11010001_0;
      patterns[30812] = 25'b01111000_01011010_11010010_0;
      patterns[30813] = 25'b01111000_01011011_11010011_0;
      patterns[30814] = 25'b01111000_01011100_11010100_0;
      patterns[30815] = 25'b01111000_01011101_11010101_0;
      patterns[30816] = 25'b01111000_01011110_11010110_0;
      patterns[30817] = 25'b01111000_01011111_11010111_0;
      patterns[30818] = 25'b01111000_01100000_11011000_0;
      patterns[30819] = 25'b01111000_01100001_11011001_0;
      patterns[30820] = 25'b01111000_01100010_11011010_0;
      patterns[30821] = 25'b01111000_01100011_11011011_0;
      patterns[30822] = 25'b01111000_01100100_11011100_0;
      patterns[30823] = 25'b01111000_01100101_11011101_0;
      patterns[30824] = 25'b01111000_01100110_11011110_0;
      patterns[30825] = 25'b01111000_01100111_11011111_0;
      patterns[30826] = 25'b01111000_01101000_11100000_0;
      patterns[30827] = 25'b01111000_01101001_11100001_0;
      patterns[30828] = 25'b01111000_01101010_11100010_0;
      patterns[30829] = 25'b01111000_01101011_11100011_0;
      patterns[30830] = 25'b01111000_01101100_11100100_0;
      patterns[30831] = 25'b01111000_01101101_11100101_0;
      patterns[30832] = 25'b01111000_01101110_11100110_0;
      patterns[30833] = 25'b01111000_01101111_11100111_0;
      patterns[30834] = 25'b01111000_01110000_11101000_0;
      patterns[30835] = 25'b01111000_01110001_11101001_0;
      patterns[30836] = 25'b01111000_01110010_11101010_0;
      patterns[30837] = 25'b01111000_01110011_11101011_0;
      patterns[30838] = 25'b01111000_01110100_11101100_0;
      patterns[30839] = 25'b01111000_01110101_11101101_0;
      patterns[30840] = 25'b01111000_01110110_11101110_0;
      patterns[30841] = 25'b01111000_01110111_11101111_0;
      patterns[30842] = 25'b01111000_01111000_11110000_0;
      patterns[30843] = 25'b01111000_01111001_11110001_0;
      patterns[30844] = 25'b01111000_01111010_11110010_0;
      patterns[30845] = 25'b01111000_01111011_11110011_0;
      patterns[30846] = 25'b01111000_01111100_11110100_0;
      patterns[30847] = 25'b01111000_01111101_11110101_0;
      patterns[30848] = 25'b01111000_01111110_11110110_0;
      patterns[30849] = 25'b01111000_01111111_11110111_0;
      patterns[30850] = 25'b01111000_10000000_11111000_0;
      patterns[30851] = 25'b01111000_10000001_11111001_0;
      patterns[30852] = 25'b01111000_10000010_11111010_0;
      patterns[30853] = 25'b01111000_10000011_11111011_0;
      patterns[30854] = 25'b01111000_10000100_11111100_0;
      patterns[30855] = 25'b01111000_10000101_11111101_0;
      patterns[30856] = 25'b01111000_10000110_11111110_0;
      patterns[30857] = 25'b01111000_10000111_11111111_0;
      patterns[30858] = 25'b01111000_10001000_00000000_1;
      patterns[30859] = 25'b01111000_10001001_00000001_1;
      patterns[30860] = 25'b01111000_10001010_00000010_1;
      patterns[30861] = 25'b01111000_10001011_00000011_1;
      patterns[30862] = 25'b01111000_10001100_00000100_1;
      patterns[30863] = 25'b01111000_10001101_00000101_1;
      patterns[30864] = 25'b01111000_10001110_00000110_1;
      patterns[30865] = 25'b01111000_10001111_00000111_1;
      patterns[30866] = 25'b01111000_10010000_00001000_1;
      patterns[30867] = 25'b01111000_10010001_00001001_1;
      patterns[30868] = 25'b01111000_10010010_00001010_1;
      patterns[30869] = 25'b01111000_10010011_00001011_1;
      patterns[30870] = 25'b01111000_10010100_00001100_1;
      patterns[30871] = 25'b01111000_10010101_00001101_1;
      patterns[30872] = 25'b01111000_10010110_00001110_1;
      patterns[30873] = 25'b01111000_10010111_00001111_1;
      patterns[30874] = 25'b01111000_10011000_00010000_1;
      patterns[30875] = 25'b01111000_10011001_00010001_1;
      patterns[30876] = 25'b01111000_10011010_00010010_1;
      patterns[30877] = 25'b01111000_10011011_00010011_1;
      patterns[30878] = 25'b01111000_10011100_00010100_1;
      patterns[30879] = 25'b01111000_10011101_00010101_1;
      patterns[30880] = 25'b01111000_10011110_00010110_1;
      patterns[30881] = 25'b01111000_10011111_00010111_1;
      patterns[30882] = 25'b01111000_10100000_00011000_1;
      patterns[30883] = 25'b01111000_10100001_00011001_1;
      patterns[30884] = 25'b01111000_10100010_00011010_1;
      patterns[30885] = 25'b01111000_10100011_00011011_1;
      patterns[30886] = 25'b01111000_10100100_00011100_1;
      patterns[30887] = 25'b01111000_10100101_00011101_1;
      patterns[30888] = 25'b01111000_10100110_00011110_1;
      patterns[30889] = 25'b01111000_10100111_00011111_1;
      patterns[30890] = 25'b01111000_10101000_00100000_1;
      patterns[30891] = 25'b01111000_10101001_00100001_1;
      patterns[30892] = 25'b01111000_10101010_00100010_1;
      patterns[30893] = 25'b01111000_10101011_00100011_1;
      patterns[30894] = 25'b01111000_10101100_00100100_1;
      patterns[30895] = 25'b01111000_10101101_00100101_1;
      patterns[30896] = 25'b01111000_10101110_00100110_1;
      patterns[30897] = 25'b01111000_10101111_00100111_1;
      patterns[30898] = 25'b01111000_10110000_00101000_1;
      patterns[30899] = 25'b01111000_10110001_00101001_1;
      patterns[30900] = 25'b01111000_10110010_00101010_1;
      patterns[30901] = 25'b01111000_10110011_00101011_1;
      patterns[30902] = 25'b01111000_10110100_00101100_1;
      patterns[30903] = 25'b01111000_10110101_00101101_1;
      patterns[30904] = 25'b01111000_10110110_00101110_1;
      patterns[30905] = 25'b01111000_10110111_00101111_1;
      patterns[30906] = 25'b01111000_10111000_00110000_1;
      patterns[30907] = 25'b01111000_10111001_00110001_1;
      patterns[30908] = 25'b01111000_10111010_00110010_1;
      patterns[30909] = 25'b01111000_10111011_00110011_1;
      patterns[30910] = 25'b01111000_10111100_00110100_1;
      patterns[30911] = 25'b01111000_10111101_00110101_1;
      patterns[30912] = 25'b01111000_10111110_00110110_1;
      patterns[30913] = 25'b01111000_10111111_00110111_1;
      patterns[30914] = 25'b01111000_11000000_00111000_1;
      patterns[30915] = 25'b01111000_11000001_00111001_1;
      patterns[30916] = 25'b01111000_11000010_00111010_1;
      patterns[30917] = 25'b01111000_11000011_00111011_1;
      patterns[30918] = 25'b01111000_11000100_00111100_1;
      patterns[30919] = 25'b01111000_11000101_00111101_1;
      patterns[30920] = 25'b01111000_11000110_00111110_1;
      patterns[30921] = 25'b01111000_11000111_00111111_1;
      patterns[30922] = 25'b01111000_11001000_01000000_1;
      patterns[30923] = 25'b01111000_11001001_01000001_1;
      patterns[30924] = 25'b01111000_11001010_01000010_1;
      patterns[30925] = 25'b01111000_11001011_01000011_1;
      patterns[30926] = 25'b01111000_11001100_01000100_1;
      patterns[30927] = 25'b01111000_11001101_01000101_1;
      patterns[30928] = 25'b01111000_11001110_01000110_1;
      patterns[30929] = 25'b01111000_11001111_01000111_1;
      patterns[30930] = 25'b01111000_11010000_01001000_1;
      patterns[30931] = 25'b01111000_11010001_01001001_1;
      patterns[30932] = 25'b01111000_11010010_01001010_1;
      patterns[30933] = 25'b01111000_11010011_01001011_1;
      patterns[30934] = 25'b01111000_11010100_01001100_1;
      patterns[30935] = 25'b01111000_11010101_01001101_1;
      patterns[30936] = 25'b01111000_11010110_01001110_1;
      patterns[30937] = 25'b01111000_11010111_01001111_1;
      patterns[30938] = 25'b01111000_11011000_01010000_1;
      patterns[30939] = 25'b01111000_11011001_01010001_1;
      patterns[30940] = 25'b01111000_11011010_01010010_1;
      patterns[30941] = 25'b01111000_11011011_01010011_1;
      patterns[30942] = 25'b01111000_11011100_01010100_1;
      patterns[30943] = 25'b01111000_11011101_01010101_1;
      patterns[30944] = 25'b01111000_11011110_01010110_1;
      patterns[30945] = 25'b01111000_11011111_01010111_1;
      patterns[30946] = 25'b01111000_11100000_01011000_1;
      patterns[30947] = 25'b01111000_11100001_01011001_1;
      patterns[30948] = 25'b01111000_11100010_01011010_1;
      patterns[30949] = 25'b01111000_11100011_01011011_1;
      patterns[30950] = 25'b01111000_11100100_01011100_1;
      patterns[30951] = 25'b01111000_11100101_01011101_1;
      patterns[30952] = 25'b01111000_11100110_01011110_1;
      patterns[30953] = 25'b01111000_11100111_01011111_1;
      patterns[30954] = 25'b01111000_11101000_01100000_1;
      patterns[30955] = 25'b01111000_11101001_01100001_1;
      patterns[30956] = 25'b01111000_11101010_01100010_1;
      patterns[30957] = 25'b01111000_11101011_01100011_1;
      patterns[30958] = 25'b01111000_11101100_01100100_1;
      patterns[30959] = 25'b01111000_11101101_01100101_1;
      patterns[30960] = 25'b01111000_11101110_01100110_1;
      patterns[30961] = 25'b01111000_11101111_01100111_1;
      patterns[30962] = 25'b01111000_11110000_01101000_1;
      patterns[30963] = 25'b01111000_11110001_01101001_1;
      patterns[30964] = 25'b01111000_11110010_01101010_1;
      patterns[30965] = 25'b01111000_11110011_01101011_1;
      patterns[30966] = 25'b01111000_11110100_01101100_1;
      patterns[30967] = 25'b01111000_11110101_01101101_1;
      patterns[30968] = 25'b01111000_11110110_01101110_1;
      patterns[30969] = 25'b01111000_11110111_01101111_1;
      patterns[30970] = 25'b01111000_11111000_01110000_1;
      patterns[30971] = 25'b01111000_11111001_01110001_1;
      patterns[30972] = 25'b01111000_11111010_01110010_1;
      patterns[30973] = 25'b01111000_11111011_01110011_1;
      patterns[30974] = 25'b01111000_11111100_01110100_1;
      patterns[30975] = 25'b01111000_11111101_01110101_1;
      patterns[30976] = 25'b01111000_11111110_01110110_1;
      patterns[30977] = 25'b01111000_11111111_01110111_1;
      patterns[30978] = 25'b01111001_00000000_01111001_0;
      patterns[30979] = 25'b01111001_00000001_01111010_0;
      patterns[30980] = 25'b01111001_00000010_01111011_0;
      patterns[30981] = 25'b01111001_00000011_01111100_0;
      patterns[30982] = 25'b01111001_00000100_01111101_0;
      patterns[30983] = 25'b01111001_00000101_01111110_0;
      patterns[30984] = 25'b01111001_00000110_01111111_0;
      patterns[30985] = 25'b01111001_00000111_10000000_0;
      patterns[30986] = 25'b01111001_00001000_10000001_0;
      patterns[30987] = 25'b01111001_00001001_10000010_0;
      patterns[30988] = 25'b01111001_00001010_10000011_0;
      patterns[30989] = 25'b01111001_00001011_10000100_0;
      patterns[30990] = 25'b01111001_00001100_10000101_0;
      patterns[30991] = 25'b01111001_00001101_10000110_0;
      patterns[30992] = 25'b01111001_00001110_10000111_0;
      patterns[30993] = 25'b01111001_00001111_10001000_0;
      patterns[30994] = 25'b01111001_00010000_10001001_0;
      patterns[30995] = 25'b01111001_00010001_10001010_0;
      patterns[30996] = 25'b01111001_00010010_10001011_0;
      patterns[30997] = 25'b01111001_00010011_10001100_0;
      patterns[30998] = 25'b01111001_00010100_10001101_0;
      patterns[30999] = 25'b01111001_00010101_10001110_0;
      patterns[31000] = 25'b01111001_00010110_10001111_0;
      patterns[31001] = 25'b01111001_00010111_10010000_0;
      patterns[31002] = 25'b01111001_00011000_10010001_0;
      patterns[31003] = 25'b01111001_00011001_10010010_0;
      patterns[31004] = 25'b01111001_00011010_10010011_0;
      patterns[31005] = 25'b01111001_00011011_10010100_0;
      patterns[31006] = 25'b01111001_00011100_10010101_0;
      patterns[31007] = 25'b01111001_00011101_10010110_0;
      patterns[31008] = 25'b01111001_00011110_10010111_0;
      patterns[31009] = 25'b01111001_00011111_10011000_0;
      patterns[31010] = 25'b01111001_00100000_10011001_0;
      patterns[31011] = 25'b01111001_00100001_10011010_0;
      patterns[31012] = 25'b01111001_00100010_10011011_0;
      patterns[31013] = 25'b01111001_00100011_10011100_0;
      patterns[31014] = 25'b01111001_00100100_10011101_0;
      patterns[31015] = 25'b01111001_00100101_10011110_0;
      patterns[31016] = 25'b01111001_00100110_10011111_0;
      patterns[31017] = 25'b01111001_00100111_10100000_0;
      patterns[31018] = 25'b01111001_00101000_10100001_0;
      patterns[31019] = 25'b01111001_00101001_10100010_0;
      patterns[31020] = 25'b01111001_00101010_10100011_0;
      patterns[31021] = 25'b01111001_00101011_10100100_0;
      patterns[31022] = 25'b01111001_00101100_10100101_0;
      patterns[31023] = 25'b01111001_00101101_10100110_0;
      patterns[31024] = 25'b01111001_00101110_10100111_0;
      patterns[31025] = 25'b01111001_00101111_10101000_0;
      patterns[31026] = 25'b01111001_00110000_10101001_0;
      patterns[31027] = 25'b01111001_00110001_10101010_0;
      patterns[31028] = 25'b01111001_00110010_10101011_0;
      patterns[31029] = 25'b01111001_00110011_10101100_0;
      patterns[31030] = 25'b01111001_00110100_10101101_0;
      patterns[31031] = 25'b01111001_00110101_10101110_0;
      patterns[31032] = 25'b01111001_00110110_10101111_0;
      patterns[31033] = 25'b01111001_00110111_10110000_0;
      patterns[31034] = 25'b01111001_00111000_10110001_0;
      patterns[31035] = 25'b01111001_00111001_10110010_0;
      patterns[31036] = 25'b01111001_00111010_10110011_0;
      patterns[31037] = 25'b01111001_00111011_10110100_0;
      patterns[31038] = 25'b01111001_00111100_10110101_0;
      patterns[31039] = 25'b01111001_00111101_10110110_0;
      patterns[31040] = 25'b01111001_00111110_10110111_0;
      patterns[31041] = 25'b01111001_00111111_10111000_0;
      patterns[31042] = 25'b01111001_01000000_10111001_0;
      patterns[31043] = 25'b01111001_01000001_10111010_0;
      patterns[31044] = 25'b01111001_01000010_10111011_0;
      patterns[31045] = 25'b01111001_01000011_10111100_0;
      patterns[31046] = 25'b01111001_01000100_10111101_0;
      patterns[31047] = 25'b01111001_01000101_10111110_0;
      patterns[31048] = 25'b01111001_01000110_10111111_0;
      patterns[31049] = 25'b01111001_01000111_11000000_0;
      patterns[31050] = 25'b01111001_01001000_11000001_0;
      patterns[31051] = 25'b01111001_01001001_11000010_0;
      patterns[31052] = 25'b01111001_01001010_11000011_0;
      patterns[31053] = 25'b01111001_01001011_11000100_0;
      patterns[31054] = 25'b01111001_01001100_11000101_0;
      patterns[31055] = 25'b01111001_01001101_11000110_0;
      patterns[31056] = 25'b01111001_01001110_11000111_0;
      patterns[31057] = 25'b01111001_01001111_11001000_0;
      patterns[31058] = 25'b01111001_01010000_11001001_0;
      patterns[31059] = 25'b01111001_01010001_11001010_0;
      patterns[31060] = 25'b01111001_01010010_11001011_0;
      patterns[31061] = 25'b01111001_01010011_11001100_0;
      patterns[31062] = 25'b01111001_01010100_11001101_0;
      patterns[31063] = 25'b01111001_01010101_11001110_0;
      patterns[31064] = 25'b01111001_01010110_11001111_0;
      patterns[31065] = 25'b01111001_01010111_11010000_0;
      patterns[31066] = 25'b01111001_01011000_11010001_0;
      patterns[31067] = 25'b01111001_01011001_11010010_0;
      patterns[31068] = 25'b01111001_01011010_11010011_0;
      patterns[31069] = 25'b01111001_01011011_11010100_0;
      patterns[31070] = 25'b01111001_01011100_11010101_0;
      patterns[31071] = 25'b01111001_01011101_11010110_0;
      patterns[31072] = 25'b01111001_01011110_11010111_0;
      patterns[31073] = 25'b01111001_01011111_11011000_0;
      patterns[31074] = 25'b01111001_01100000_11011001_0;
      patterns[31075] = 25'b01111001_01100001_11011010_0;
      patterns[31076] = 25'b01111001_01100010_11011011_0;
      patterns[31077] = 25'b01111001_01100011_11011100_0;
      patterns[31078] = 25'b01111001_01100100_11011101_0;
      patterns[31079] = 25'b01111001_01100101_11011110_0;
      patterns[31080] = 25'b01111001_01100110_11011111_0;
      patterns[31081] = 25'b01111001_01100111_11100000_0;
      patterns[31082] = 25'b01111001_01101000_11100001_0;
      patterns[31083] = 25'b01111001_01101001_11100010_0;
      patterns[31084] = 25'b01111001_01101010_11100011_0;
      patterns[31085] = 25'b01111001_01101011_11100100_0;
      patterns[31086] = 25'b01111001_01101100_11100101_0;
      patterns[31087] = 25'b01111001_01101101_11100110_0;
      patterns[31088] = 25'b01111001_01101110_11100111_0;
      patterns[31089] = 25'b01111001_01101111_11101000_0;
      patterns[31090] = 25'b01111001_01110000_11101001_0;
      patterns[31091] = 25'b01111001_01110001_11101010_0;
      patterns[31092] = 25'b01111001_01110010_11101011_0;
      patterns[31093] = 25'b01111001_01110011_11101100_0;
      patterns[31094] = 25'b01111001_01110100_11101101_0;
      patterns[31095] = 25'b01111001_01110101_11101110_0;
      patterns[31096] = 25'b01111001_01110110_11101111_0;
      patterns[31097] = 25'b01111001_01110111_11110000_0;
      patterns[31098] = 25'b01111001_01111000_11110001_0;
      patterns[31099] = 25'b01111001_01111001_11110010_0;
      patterns[31100] = 25'b01111001_01111010_11110011_0;
      patterns[31101] = 25'b01111001_01111011_11110100_0;
      patterns[31102] = 25'b01111001_01111100_11110101_0;
      patterns[31103] = 25'b01111001_01111101_11110110_0;
      patterns[31104] = 25'b01111001_01111110_11110111_0;
      patterns[31105] = 25'b01111001_01111111_11111000_0;
      patterns[31106] = 25'b01111001_10000000_11111001_0;
      patterns[31107] = 25'b01111001_10000001_11111010_0;
      patterns[31108] = 25'b01111001_10000010_11111011_0;
      patterns[31109] = 25'b01111001_10000011_11111100_0;
      patterns[31110] = 25'b01111001_10000100_11111101_0;
      patterns[31111] = 25'b01111001_10000101_11111110_0;
      patterns[31112] = 25'b01111001_10000110_11111111_0;
      patterns[31113] = 25'b01111001_10000111_00000000_1;
      patterns[31114] = 25'b01111001_10001000_00000001_1;
      patterns[31115] = 25'b01111001_10001001_00000010_1;
      patterns[31116] = 25'b01111001_10001010_00000011_1;
      patterns[31117] = 25'b01111001_10001011_00000100_1;
      patterns[31118] = 25'b01111001_10001100_00000101_1;
      patterns[31119] = 25'b01111001_10001101_00000110_1;
      patterns[31120] = 25'b01111001_10001110_00000111_1;
      patterns[31121] = 25'b01111001_10001111_00001000_1;
      patterns[31122] = 25'b01111001_10010000_00001001_1;
      patterns[31123] = 25'b01111001_10010001_00001010_1;
      patterns[31124] = 25'b01111001_10010010_00001011_1;
      patterns[31125] = 25'b01111001_10010011_00001100_1;
      patterns[31126] = 25'b01111001_10010100_00001101_1;
      patterns[31127] = 25'b01111001_10010101_00001110_1;
      patterns[31128] = 25'b01111001_10010110_00001111_1;
      patterns[31129] = 25'b01111001_10010111_00010000_1;
      patterns[31130] = 25'b01111001_10011000_00010001_1;
      patterns[31131] = 25'b01111001_10011001_00010010_1;
      patterns[31132] = 25'b01111001_10011010_00010011_1;
      patterns[31133] = 25'b01111001_10011011_00010100_1;
      patterns[31134] = 25'b01111001_10011100_00010101_1;
      patterns[31135] = 25'b01111001_10011101_00010110_1;
      patterns[31136] = 25'b01111001_10011110_00010111_1;
      patterns[31137] = 25'b01111001_10011111_00011000_1;
      patterns[31138] = 25'b01111001_10100000_00011001_1;
      patterns[31139] = 25'b01111001_10100001_00011010_1;
      patterns[31140] = 25'b01111001_10100010_00011011_1;
      patterns[31141] = 25'b01111001_10100011_00011100_1;
      patterns[31142] = 25'b01111001_10100100_00011101_1;
      patterns[31143] = 25'b01111001_10100101_00011110_1;
      patterns[31144] = 25'b01111001_10100110_00011111_1;
      patterns[31145] = 25'b01111001_10100111_00100000_1;
      patterns[31146] = 25'b01111001_10101000_00100001_1;
      patterns[31147] = 25'b01111001_10101001_00100010_1;
      patterns[31148] = 25'b01111001_10101010_00100011_1;
      patterns[31149] = 25'b01111001_10101011_00100100_1;
      patterns[31150] = 25'b01111001_10101100_00100101_1;
      patterns[31151] = 25'b01111001_10101101_00100110_1;
      patterns[31152] = 25'b01111001_10101110_00100111_1;
      patterns[31153] = 25'b01111001_10101111_00101000_1;
      patterns[31154] = 25'b01111001_10110000_00101001_1;
      patterns[31155] = 25'b01111001_10110001_00101010_1;
      patterns[31156] = 25'b01111001_10110010_00101011_1;
      patterns[31157] = 25'b01111001_10110011_00101100_1;
      patterns[31158] = 25'b01111001_10110100_00101101_1;
      patterns[31159] = 25'b01111001_10110101_00101110_1;
      patterns[31160] = 25'b01111001_10110110_00101111_1;
      patterns[31161] = 25'b01111001_10110111_00110000_1;
      patterns[31162] = 25'b01111001_10111000_00110001_1;
      patterns[31163] = 25'b01111001_10111001_00110010_1;
      patterns[31164] = 25'b01111001_10111010_00110011_1;
      patterns[31165] = 25'b01111001_10111011_00110100_1;
      patterns[31166] = 25'b01111001_10111100_00110101_1;
      patterns[31167] = 25'b01111001_10111101_00110110_1;
      patterns[31168] = 25'b01111001_10111110_00110111_1;
      patterns[31169] = 25'b01111001_10111111_00111000_1;
      patterns[31170] = 25'b01111001_11000000_00111001_1;
      patterns[31171] = 25'b01111001_11000001_00111010_1;
      patterns[31172] = 25'b01111001_11000010_00111011_1;
      patterns[31173] = 25'b01111001_11000011_00111100_1;
      patterns[31174] = 25'b01111001_11000100_00111101_1;
      patterns[31175] = 25'b01111001_11000101_00111110_1;
      patterns[31176] = 25'b01111001_11000110_00111111_1;
      patterns[31177] = 25'b01111001_11000111_01000000_1;
      patterns[31178] = 25'b01111001_11001000_01000001_1;
      patterns[31179] = 25'b01111001_11001001_01000010_1;
      patterns[31180] = 25'b01111001_11001010_01000011_1;
      patterns[31181] = 25'b01111001_11001011_01000100_1;
      patterns[31182] = 25'b01111001_11001100_01000101_1;
      patterns[31183] = 25'b01111001_11001101_01000110_1;
      patterns[31184] = 25'b01111001_11001110_01000111_1;
      patterns[31185] = 25'b01111001_11001111_01001000_1;
      patterns[31186] = 25'b01111001_11010000_01001001_1;
      patterns[31187] = 25'b01111001_11010001_01001010_1;
      patterns[31188] = 25'b01111001_11010010_01001011_1;
      patterns[31189] = 25'b01111001_11010011_01001100_1;
      patterns[31190] = 25'b01111001_11010100_01001101_1;
      patterns[31191] = 25'b01111001_11010101_01001110_1;
      patterns[31192] = 25'b01111001_11010110_01001111_1;
      patterns[31193] = 25'b01111001_11010111_01010000_1;
      patterns[31194] = 25'b01111001_11011000_01010001_1;
      patterns[31195] = 25'b01111001_11011001_01010010_1;
      patterns[31196] = 25'b01111001_11011010_01010011_1;
      patterns[31197] = 25'b01111001_11011011_01010100_1;
      patterns[31198] = 25'b01111001_11011100_01010101_1;
      patterns[31199] = 25'b01111001_11011101_01010110_1;
      patterns[31200] = 25'b01111001_11011110_01010111_1;
      patterns[31201] = 25'b01111001_11011111_01011000_1;
      patterns[31202] = 25'b01111001_11100000_01011001_1;
      patterns[31203] = 25'b01111001_11100001_01011010_1;
      patterns[31204] = 25'b01111001_11100010_01011011_1;
      patterns[31205] = 25'b01111001_11100011_01011100_1;
      patterns[31206] = 25'b01111001_11100100_01011101_1;
      patterns[31207] = 25'b01111001_11100101_01011110_1;
      patterns[31208] = 25'b01111001_11100110_01011111_1;
      patterns[31209] = 25'b01111001_11100111_01100000_1;
      patterns[31210] = 25'b01111001_11101000_01100001_1;
      patterns[31211] = 25'b01111001_11101001_01100010_1;
      patterns[31212] = 25'b01111001_11101010_01100011_1;
      patterns[31213] = 25'b01111001_11101011_01100100_1;
      patterns[31214] = 25'b01111001_11101100_01100101_1;
      patterns[31215] = 25'b01111001_11101101_01100110_1;
      patterns[31216] = 25'b01111001_11101110_01100111_1;
      patterns[31217] = 25'b01111001_11101111_01101000_1;
      patterns[31218] = 25'b01111001_11110000_01101001_1;
      patterns[31219] = 25'b01111001_11110001_01101010_1;
      patterns[31220] = 25'b01111001_11110010_01101011_1;
      patterns[31221] = 25'b01111001_11110011_01101100_1;
      patterns[31222] = 25'b01111001_11110100_01101101_1;
      patterns[31223] = 25'b01111001_11110101_01101110_1;
      patterns[31224] = 25'b01111001_11110110_01101111_1;
      patterns[31225] = 25'b01111001_11110111_01110000_1;
      patterns[31226] = 25'b01111001_11111000_01110001_1;
      patterns[31227] = 25'b01111001_11111001_01110010_1;
      patterns[31228] = 25'b01111001_11111010_01110011_1;
      patterns[31229] = 25'b01111001_11111011_01110100_1;
      patterns[31230] = 25'b01111001_11111100_01110101_1;
      patterns[31231] = 25'b01111001_11111101_01110110_1;
      patterns[31232] = 25'b01111001_11111110_01110111_1;
      patterns[31233] = 25'b01111001_11111111_01111000_1;
      patterns[31234] = 25'b01111010_00000000_01111010_0;
      patterns[31235] = 25'b01111010_00000001_01111011_0;
      patterns[31236] = 25'b01111010_00000010_01111100_0;
      patterns[31237] = 25'b01111010_00000011_01111101_0;
      patterns[31238] = 25'b01111010_00000100_01111110_0;
      patterns[31239] = 25'b01111010_00000101_01111111_0;
      patterns[31240] = 25'b01111010_00000110_10000000_0;
      patterns[31241] = 25'b01111010_00000111_10000001_0;
      patterns[31242] = 25'b01111010_00001000_10000010_0;
      patterns[31243] = 25'b01111010_00001001_10000011_0;
      patterns[31244] = 25'b01111010_00001010_10000100_0;
      patterns[31245] = 25'b01111010_00001011_10000101_0;
      patterns[31246] = 25'b01111010_00001100_10000110_0;
      patterns[31247] = 25'b01111010_00001101_10000111_0;
      patterns[31248] = 25'b01111010_00001110_10001000_0;
      patterns[31249] = 25'b01111010_00001111_10001001_0;
      patterns[31250] = 25'b01111010_00010000_10001010_0;
      patterns[31251] = 25'b01111010_00010001_10001011_0;
      patterns[31252] = 25'b01111010_00010010_10001100_0;
      patterns[31253] = 25'b01111010_00010011_10001101_0;
      patterns[31254] = 25'b01111010_00010100_10001110_0;
      patterns[31255] = 25'b01111010_00010101_10001111_0;
      patterns[31256] = 25'b01111010_00010110_10010000_0;
      patterns[31257] = 25'b01111010_00010111_10010001_0;
      patterns[31258] = 25'b01111010_00011000_10010010_0;
      patterns[31259] = 25'b01111010_00011001_10010011_0;
      patterns[31260] = 25'b01111010_00011010_10010100_0;
      patterns[31261] = 25'b01111010_00011011_10010101_0;
      patterns[31262] = 25'b01111010_00011100_10010110_0;
      patterns[31263] = 25'b01111010_00011101_10010111_0;
      patterns[31264] = 25'b01111010_00011110_10011000_0;
      patterns[31265] = 25'b01111010_00011111_10011001_0;
      patterns[31266] = 25'b01111010_00100000_10011010_0;
      patterns[31267] = 25'b01111010_00100001_10011011_0;
      patterns[31268] = 25'b01111010_00100010_10011100_0;
      patterns[31269] = 25'b01111010_00100011_10011101_0;
      patterns[31270] = 25'b01111010_00100100_10011110_0;
      patterns[31271] = 25'b01111010_00100101_10011111_0;
      patterns[31272] = 25'b01111010_00100110_10100000_0;
      patterns[31273] = 25'b01111010_00100111_10100001_0;
      patterns[31274] = 25'b01111010_00101000_10100010_0;
      patterns[31275] = 25'b01111010_00101001_10100011_0;
      patterns[31276] = 25'b01111010_00101010_10100100_0;
      patterns[31277] = 25'b01111010_00101011_10100101_0;
      patterns[31278] = 25'b01111010_00101100_10100110_0;
      patterns[31279] = 25'b01111010_00101101_10100111_0;
      patterns[31280] = 25'b01111010_00101110_10101000_0;
      patterns[31281] = 25'b01111010_00101111_10101001_0;
      patterns[31282] = 25'b01111010_00110000_10101010_0;
      patterns[31283] = 25'b01111010_00110001_10101011_0;
      patterns[31284] = 25'b01111010_00110010_10101100_0;
      patterns[31285] = 25'b01111010_00110011_10101101_0;
      patterns[31286] = 25'b01111010_00110100_10101110_0;
      patterns[31287] = 25'b01111010_00110101_10101111_0;
      patterns[31288] = 25'b01111010_00110110_10110000_0;
      patterns[31289] = 25'b01111010_00110111_10110001_0;
      patterns[31290] = 25'b01111010_00111000_10110010_0;
      patterns[31291] = 25'b01111010_00111001_10110011_0;
      patterns[31292] = 25'b01111010_00111010_10110100_0;
      patterns[31293] = 25'b01111010_00111011_10110101_0;
      patterns[31294] = 25'b01111010_00111100_10110110_0;
      patterns[31295] = 25'b01111010_00111101_10110111_0;
      patterns[31296] = 25'b01111010_00111110_10111000_0;
      patterns[31297] = 25'b01111010_00111111_10111001_0;
      patterns[31298] = 25'b01111010_01000000_10111010_0;
      patterns[31299] = 25'b01111010_01000001_10111011_0;
      patterns[31300] = 25'b01111010_01000010_10111100_0;
      patterns[31301] = 25'b01111010_01000011_10111101_0;
      patterns[31302] = 25'b01111010_01000100_10111110_0;
      patterns[31303] = 25'b01111010_01000101_10111111_0;
      patterns[31304] = 25'b01111010_01000110_11000000_0;
      patterns[31305] = 25'b01111010_01000111_11000001_0;
      patterns[31306] = 25'b01111010_01001000_11000010_0;
      patterns[31307] = 25'b01111010_01001001_11000011_0;
      patterns[31308] = 25'b01111010_01001010_11000100_0;
      patterns[31309] = 25'b01111010_01001011_11000101_0;
      patterns[31310] = 25'b01111010_01001100_11000110_0;
      patterns[31311] = 25'b01111010_01001101_11000111_0;
      patterns[31312] = 25'b01111010_01001110_11001000_0;
      patterns[31313] = 25'b01111010_01001111_11001001_0;
      patterns[31314] = 25'b01111010_01010000_11001010_0;
      patterns[31315] = 25'b01111010_01010001_11001011_0;
      patterns[31316] = 25'b01111010_01010010_11001100_0;
      patterns[31317] = 25'b01111010_01010011_11001101_0;
      patterns[31318] = 25'b01111010_01010100_11001110_0;
      patterns[31319] = 25'b01111010_01010101_11001111_0;
      patterns[31320] = 25'b01111010_01010110_11010000_0;
      patterns[31321] = 25'b01111010_01010111_11010001_0;
      patterns[31322] = 25'b01111010_01011000_11010010_0;
      patterns[31323] = 25'b01111010_01011001_11010011_0;
      patterns[31324] = 25'b01111010_01011010_11010100_0;
      patterns[31325] = 25'b01111010_01011011_11010101_0;
      patterns[31326] = 25'b01111010_01011100_11010110_0;
      patterns[31327] = 25'b01111010_01011101_11010111_0;
      patterns[31328] = 25'b01111010_01011110_11011000_0;
      patterns[31329] = 25'b01111010_01011111_11011001_0;
      patterns[31330] = 25'b01111010_01100000_11011010_0;
      patterns[31331] = 25'b01111010_01100001_11011011_0;
      patterns[31332] = 25'b01111010_01100010_11011100_0;
      patterns[31333] = 25'b01111010_01100011_11011101_0;
      patterns[31334] = 25'b01111010_01100100_11011110_0;
      patterns[31335] = 25'b01111010_01100101_11011111_0;
      patterns[31336] = 25'b01111010_01100110_11100000_0;
      patterns[31337] = 25'b01111010_01100111_11100001_0;
      patterns[31338] = 25'b01111010_01101000_11100010_0;
      patterns[31339] = 25'b01111010_01101001_11100011_0;
      patterns[31340] = 25'b01111010_01101010_11100100_0;
      patterns[31341] = 25'b01111010_01101011_11100101_0;
      patterns[31342] = 25'b01111010_01101100_11100110_0;
      patterns[31343] = 25'b01111010_01101101_11100111_0;
      patterns[31344] = 25'b01111010_01101110_11101000_0;
      patterns[31345] = 25'b01111010_01101111_11101001_0;
      patterns[31346] = 25'b01111010_01110000_11101010_0;
      patterns[31347] = 25'b01111010_01110001_11101011_0;
      patterns[31348] = 25'b01111010_01110010_11101100_0;
      patterns[31349] = 25'b01111010_01110011_11101101_0;
      patterns[31350] = 25'b01111010_01110100_11101110_0;
      patterns[31351] = 25'b01111010_01110101_11101111_0;
      patterns[31352] = 25'b01111010_01110110_11110000_0;
      patterns[31353] = 25'b01111010_01110111_11110001_0;
      patterns[31354] = 25'b01111010_01111000_11110010_0;
      patterns[31355] = 25'b01111010_01111001_11110011_0;
      patterns[31356] = 25'b01111010_01111010_11110100_0;
      patterns[31357] = 25'b01111010_01111011_11110101_0;
      patterns[31358] = 25'b01111010_01111100_11110110_0;
      patterns[31359] = 25'b01111010_01111101_11110111_0;
      patterns[31360] = 25'b01111010_01111110_11111000_0;
      patterns[31361] = 25'b01111010_01111111_11111001_0;
      patterns[31362] = 25'b01111010_10000000_11111010_0;
      patterns[31363] = 25'b01111010_10000001_11111011_0;
      patterns[31364] = 25'b01111010_10000010_11111100_0;
      patterns[31365] = 25'b01111010_10000011_11111101_0;
      patterns[31366] = 25'b01111010_10000100_11111110_0;
      patterns[31367] = 25'b01111010_10000101_11111111_0;
      patterns[31368] = 25'b01111010_10000110_00000000_1;
      patterns[31369] = 25'b01111010_10000111_00000001_1;
      patterns[31370] = 25'b01111010_10001000_00000010_1;
      patterns[31371] = 25'b01111010_10001001_00000011_1;
      patterns[31372] = 25'b01111010_10001010_00000100_1;
      patterns[31373] = 25'b01111010_10001011_00000101_1;
      patterns[31374] = 25'b01111010_10001100_00000110_1;
      patterns[31375] = 25'b01111010_10001101_00000111_1;
      patterns[31376] = 25'b01111010_10001110_00001000_1;
      patterns[31377] = 25'b01111010_10001111_00001001_1;
      patterns[31378] = 25'b01111010_10010000_00001010_1;
      patterns[31379] = 25'b01111010_10010001_00001011_1;
      patterns[31380] = 25'b01111010_10010010_00001100_1;
      patterns[31381] = 25'b01111010_10010011_00001101_1;
      patterns[31382] = 25'b01111010_10010100_00001110_1;
      patterns[31383] = 25'b01111010_10010101_00001111_1;
      patterns[31384] = 25'b01111010_10010110_00010000_1;
      patterns[31385] = 25'b01111010_10010111_00010001_1;
      patterns[31386] = 25'b01111010_10011000_00010010_1;
      patterns[31387] = 25'b01111010_10011001_00010011_1;
      patterns[31388] = 25'b01111010_10011010_00010100_1;
      patterns[31389] = 25'b01111010_10011011_00010101_1;
      patterns[31390] = 25'b01111010_10011100_00010110_1;
      patterns[31391] = 25'b01111010_10011101_00010111_1;
      patterns[31392] = 25'b01111010_10011110_00011000_1;
      patterns[31393] = 25'b01111010_10011111_00011001_1;
      patterns[31394] = 25'b01111010_10100000_00011010_1;
      patterns[31395] = 25'b01111010_10100001_00011011_1;
      patterns[31396] = 25'b01111010_10100010_00011100_1;
      patterns[31397] = 25'b01111010_10100011_00011101_1;
      patterns[31398] = 25'b01111010_10100100_00011110_1;
      patterns[31399] = 25'b01111010_10100101_00011111_1;
      patterns[31400] = 25'b01111010_10100110_00100000_1;
      patterns[31401] = 25'b01111010_10100111_00100001_1;
      patterns[31402] = 25'b01111010_10101000_00100010_1;
      patterns[31403] = 25'b01111010_10101001_00100011_1;
      patterns[31404] = 25'b01111010_10101010_00100100_1;
      patterns[31405] = 25'b01111010_10101011_00100101_1;
      patterns[31406] = 25'b01111010_10101100_00100110_1;
      patterns[31407] = 25'b01111010_10101101_00100111_1;
      patterns[31408] = 25'b01111010_10101110_00101000_1;
      patterns[31409] = 25'b01111010_10101111_00101001_1;
      patterns[31410] = 25'b01111010_10110000_00101010_1;
      patterns[31411] = 25'b01111010_10110001_00101011_1;
      patterns[31412] = 25'b01111010_10110010_00101100_1;
      patterns[31413] = 25'b01111010_10110011_00101101_1;
      patterns[31414] = 25'b01111010_10110100_00101110_1;
      patterns[31415] = 25'b01111010_10110101_00101111_1;
      patterns[31416] = 25'b01111010_10110110_00110000_1;
      patterns[31417] = 25'b01111010_10110111_00110001_1;
      patterns[31418] = 25'b01111010_10111000_00110010_1;
      patterns[31419] = 25'b01111010_10111001_00110011_1;
      patterns[31420] = 25'b01111010_10111010_00110100_1;
      patterns[31421] = 25'b01111010_10111011_00110101_1;
      patterns[31422] = 25'b01111010_10111100_00110110_1;
      patterns[31423] = 25'b01111010_10111101_00110111_1;
      patterns[31424] = 25'b01111010_10111110_00111000_1;
      patterns[31425] = 25'b01111010_10111111_00111001_1;
      patterns[31426] = 25'b01111010_11000000_00111010_1;
      patterns[31427] = 25'b01111010_11000001_00111011_1;
      patterns[31428] = 25'b01111010_11000010_00111100_1;
      patterns[31429] = 25'b01111010_11000011_00111101_1;
      patterns[31430] = 25'b01111010_11000100_00111110_1;
      patterns[31431] = 25'b01111010_11000101_00111111_1;
      patterns[31432] = 25'b01111010_11000110_01000000_1;
      patterns[31433] = 25'b01111010_11000111_01000001_1;
      patterns[31434] = 25'b01111010_11001000_01000010_1;
      patterns[31435] = 25'b01111010_11001001_01000011_1;
      patterns[31436] = 25'b01111010_11001010_01000100_1;
      patterns[31437] = 25'b01111010_11001011_01000101_1;
      patterns[31438] = 25'b01111010_11001100_01000110_1;
      patterns[31439] = 25'b01111010_11001101_01000111_1;
      patterns[31440] = 25'b01111010_11001110_01001000_1;
      patterns[31441] = 25'b01111010_11001111_01001001_1;
      patterns[31442] = 25'b01111010_11010000_01001010_1;
      patterns[31443] = 25'b01111010_11010001_01001011_1;
      patterns[31444] = 25'b01111010_11010010_01001100_1;
      patterns[31445] = 25'b01111010_11010011_01001101_1;
      patterns[31446] = 25'b01111010_11010100_01001110_1;
      patterns[31447] = 25'b01111010_11010101_01001111_1;
      patterns[31448] = 25'b01111010_11010110_01010000_1;
      patterns[31449] = 25'b01111010_11010111_01010001_1;
      patterns[31450] = 25'b01111010_11011000_01010010_1;
      patterns[31451] = 25'b01111010_11011001_01010011_1;
      patterns[31452] = 25'b01111010_11011010_01010100_1;
      patterns[31453] = 25'b01111010_11011011_01010101_1;
      patterns[31454] = 25'b01111010_11011100_01010110_1;
      patterns[31455] = 25'b01111010_11011101_01010111_1;
      patterns[31456] = 25'b01111010_11011110_01011000_1;
      patterns[31457] = 25'b01111010_11011111_01011001_1;
      patterns[31458] = 25'b01111010_11100000_01011010_1;
      patterns[31459] = 25'b01111010_11100001_01011011_1;
      patterns[31460] = 25'b01111010_11100010_01011100_1;
      patterns[31461] = 25'b01111010_11100011_01011101_1;
      patterns[31462] = 25'b01111010_11100100_01011110_1;
      patterns[31463] = 25'b01111010_11100101_01011111_1;
      patterns[31464] = 25'b01111010_11100110_01100000_1;
      patterns[31465] = 25'b01111010_11100111_01100001_1;
      patterns[31466] = 25'b01111010_11101000_01100010_1;
      patterns[31467] = 25'b01111010_11101001_01100011_1;
      patterns[31468] = 25'b01111010_11101010_01100100_1;
      patterns[31469] = 25'b01111010_11101011_01100101_1;
      patterns[31470] = 25'b01111010_11101100_01100110_1;
      patterns[31471] = 25'b01111010_11101101_01100111_1;
      patterns[31472] = 25'b01111010_11101110_01101000_1;
      patterns[31473] = 25'b01111010_11101111_01101001_1;
      patterns[31474] = 25'b01111010_11110000_01101010_1;
      patterns[31475] = 25'b01111010_11110001_01101011_1;
      patterns[31476] = 25'b01111010_11110010_01101100_1;
      patterns[31477] = 25'b01111010_11110011_01101101_1;
      patterns[31478] = 25'b01111010_11110100_01101110_1;
      patterns[31479] = 25'b01111010_11110101_01101111_1;
      patterns[31480] = 25'b01111010_11110110_01110000_1;
      patterns[31481] = 25'b01111010_11110111_01110001_1;
      patterns[31482] = 25'b01111010_11111000_01110010_1;
      patterns[31483] = 25'b01111010_11111001_01110011_1;
      patterns[31484] = 25'b01111010_11111010_01110100_1;
      patterns[31485] = 25'b01111010_11111011_01110101_1;
      patterns[31486] = 25'b01111010_11111100_01110110_1;
      patterns[31487] = 25'b01111010_11111101_01110111_1;
      patterns[31488] = 25'b01111010_11111110_01111000_1;
      patterns[31489] = 25'b01111010_11111111_01111001_1;
      patterns[31490] = 25'b01111011_00000000_01111011_0;
      patterns[31491] = 25'b01111011_00000001_01111100_0;
      patterns[31492] = 25'b01111011_00000010_01111101_0;
      patterns[31493] = 25'b01111011_00000011_01111110_0;
      patterns[31494] = 25'b01111011_00000100_01111111_0;
      patterns[31495] = 25'b01111011_00000101_10000000_0;
      patterns[31496] = 25'b01111011_00000110_10000001_0;
      patterns[31497] = 25'b01111011_00000111_10000010_0;
      patterns[31498] = 25'b01111011_00001000_10000011_0;
      patterns[31499] = 25'b01111011_00001001_10000100_0;
      patterns[31500] = 25'b01111011_00001010_10000101_0;
      patterns[31501] = 25'b01111011_00001011_10000110_0;
      patterns[31502] = 25'b01111011_00001100_10000111_0;
      patterns[31503] = 25'b01111011_00001101_10001000_0;
      patterns[31504] = 25'b01111011_00001110_10001001_0;
      patterns[31505] = 25'b01111011_00001111_10001010_0;
      patterns[31506] = 25'b01111011_00010000_10001011_0;
      patterns[31507] = 25'b01111011_00010001_10001100_0;
      patterns[31508] = 25'b01111011_00010010_10001101_0;
      patterns[31509] = 25'b01111011_00010011_10001110_0;
      patterns[31510] = 25'b01111011_00010100_10001111_0;
      patterns[31511] = 25'b01111011_00010101_10010000_0;
      patterns[31512] = 25'b01111011_00010110_10010001_0;
      patterns[31513] = 25'b01111011_00010111_10010010_0;
      patterns[31514] = 25'b01111011_00011000_10010011_0;
      patterns[31515] = 25'b01111011_00011001_10010100_0;
      patterns[31516] = 25'b01111011_00011010_10010101_0;
      patterns[31517] = 25'b01111011_00011011_10010110_0;
      patterns[31518] = 25'b01111011_00011100_10010111_0;
      patterns[31519] = 25'b01111011_00011101_10011000_0;
      patterns[31520] = 25'b01111011_00011110_10011001_0;
      patterns[31521] = 25'b01111011_00011111_10011010_0;
      patterns[31522] = 25'b01111011_00100000_10011011_0;
      patterns[31523] = 25'b01111011_00100001_10011100_0;
      patterns[31524] = 25'b01111011_00100010_10011101_0;
      patterns[31525] = 25'b01111011_00100011_10011110_0;
      patterns[31526] = 25'b01111011_00100100_10011111_0;
      patterns[31527] = 25'b01111011_00100101_10100000_0;
      patterns[31528] = 25'b01111011_00100110_10100001_0;
      patterns[31529] = 25'b01111011_00100111_10100010_0;
      patterns[31530] = 25'b01111011_00101000_10100011_0;
      patterns[31531] = 25'b01111011_00101001_10100100_0;
      patterns[31532] = 25'b01111011_00101010_10100101_0;
      patterns[31533] = 25'b01111011_00101011_10100110_0;
      patterns[31534] = 25'b01111011_00101100_10100111_0;
      patterns[31535] = 25'b01111011_00101101_10101000_0;
      patterns[31536] = 25'b01111011_00101110_10101001_0;
      patterns[31537] = 25'b01111011_00101111_10101010_0;
      patterns[31538] = 25'b01111011_00110000_10101011_0;
      patterns[31539] = 25'b01111011_00110001_10101100_0;
      patterns[31540] = 25'b01111011_00110010_10101101_0;
      patterns[31541] = 25'b01111011_00110011_10101110_0;
      patterns[31542] = 25'b01111011_00110100_10101111_0;
      patterns[31543] = 25'b01111011_00110101_10110000_0;
      patterns[31544] = 25'b01111011_00110110_10110001_0;
      patterns[31545] = 25'b01111011_00110111_10110010_0;
      patterns[31546] = 25'b01111011_00111000_10110011_0;
      patterns[31547] = 25'b01111011_00111001_10110100_0;
      patterns[31548] = 25'b01111011_00111010_10110101_0;
      patterns[31549] = 25'b01111011_00111011_10110110_0;
      patterns[31550] = 25'b01111011_00111100_10110111_0;
      patterns[31551] = 25'b01111011_00111101_10111000_0;
      patterns[31552] = 25'b01111011_00111110_10111001_0;
      patterns[31553] = 25'b01111011_00111111_10111010_0;
      patterns[31554] = 25'b01111011_01000000_10111011_0;
      patterns[31555] = 25'b01111011_01000001_10111100_0;
      patterns[31556] = 25'b01111011_01000010_10111101_0;
      patterns[31557] = 25'b01111011_01000011_10111110_0;
      patterns[31558] = 25'b01111011_01000100_10111111_0;
      patterns[31559] = 25'b01111011_01000101_11000000_0;
      patterns[31560] = 25'b01111011_01000110_11000001_0;
      patterns[31561] = 25'b01111011_01000111_11000010_0;
      patterns[31562] = 25'b01111011_01001000_11000011_0;
      patterns[31563] = 25'b01111011_01001001_11000100_0;
      patterns[31564] = 25'b01111011_01001010_11000101_0;
      patterns[31565] = 25'b01111011_01001011_11000110_0;
      patterns[31566] = 25'b01111011_01001100_11000111_0;
      patterns[31567] = 25'b01111011_01001101_11001000_0;
      patterns[31568] = 25'b01111011_01001110_11001001_0;
      patterns[31569] = 25'b01111011_01001111_11001010_0;
      patterns[31570] = 25'b01111011_01010000_11001011_0;
      patterns[31571] = 25'b01111011_01010001_11001100_0;
      patterns[31572] = 25'b01111011_01010010_11001101_0;
      patterns[31573] = 25'b01111011_01010011_11001110_0;
      patterns[31574] = 25'b01111011_01010100_11001111_0;
      patterns[31575] = 25'b01111011_01010101_11010000_0;
      patterns[31576] = 25'b01111011_01010110_11010001_0;
      patterns[31577] = 25'b01111011_01010111_11010010_0;
      patterns[31578] = 25'b01111011_01011000_11010011_0;
      patterns[31579] = 25'b01111011_01011001_11010100_0;
      patterns[31580] = 25'b01111011_01011010_11010101_0;
      patterns[31581] = 25'b01111011_01011011_11010110_0;
      patterns[31582] = 25'b01111011_01011100_11010111_0;
      patterns[31583] = 25'b01111011_01011101_11011000_0;
      patterns[31584] = 25'b01111011_01011110_11011001_0;
      patterns[31585] = 25'b01111011_01011111_11011010_0;
      patterns[31586] = 25'b01111011_01100000_11011011_0;
      patterns[31587] = 25'b01111011_01100001_11011100_0;
      patterns[31588] = 25'b01111011_01100010_11011101_0;
      patterns[31589] = 25'b01111011_01100011_11011110_0;
      patterns[31590] = 25'b01111011_01100100_11011111_0;
      patterns[31591] = 25'b01111011_01100101_11100000_0;
      patterns[31592] = 25'b01111011_01100110_11100001_0;
      patterns[31593] = 25'b01111011_01100111_11100010_0;
      patterns[31594] = 25'b01111011_01101000_11100011_0;
      patterns[31595] = 25'b01111011_01101001_11100100_0;
      patterns[31596] = 25'b01111011_01101010_11100101_0;
      patterns[31597] = 25'b01111011_01101011_11100110_0;
      patterns[31598] = 25'b01111011_01101100_11100111_0;
      patterns[31599] = 25'b01111011_01101101_11101000_0;
      patterns[31600] = 25'b01111011_01101110_11101001_0;
      patterns[31601] = 25'b01111011_01101111_11101010_0;
      patterns[31602] = 25'b01111011_01110000_11101011_0;
      patterns[31603] = 25'b01111011_01110001_11101100_0;
      patterns[31604] = 25'b01111011_01110010_11101101_0;
      patterns[31605] = 25'b01111011_01110011_11101110_0;
      patterns[31606] = 25'b01111011_01110100_11101111_0;
      patterns[31607] = 25'b01111011_01110101_11110000_0;
      patterns[31608] = 25'b01111011_01110110_11110001_0;
      patterns[31609] = 25'b01111011_01110111_11110010_0;
      patterns[31610] = 25'b01111011_01111000_11110011_0;
      patterns[31611] = 25'b01111011_01111001_11110100_0;
      patterns[31612] = 25'b01111011_01111010_11110101_0;
      patterns[31613] = 25'b01111011_01111011_11110110_0;
      patterns[31614] = 25'b01111011_01111100_11110111_0;
      patterns[31615] = 25'b01111011_01111101_11111000_0;
      patterns[31616] = 25'b01111011_01111110_11111001_0;
      patterns[31617] = 25'b01111011_01111111_11111010_0;
      patterns[31618] = 25'b01111011_10000000_11111011_0;
      patterns[31619] = 25'b01111011_10000001_11111100_0;
      patterns[31620] = 25'b01111011_10000010_11111101_0;
      patterns[31621] = 25'b01111011_10000011_11111110_0;
      patterns[31622] = 25'b01111011_10000100_11111111_0;
      patterns[31623] = 25'b01111011_10000101_00000000_1;
      patterns[31624] = 25'b01111011_10000110_00000001_1;
      patterns[31625] = 25'b01111011_10000111_00000010_1;
      patterns[31626] = 25'b01111011_10001000_00000011_1;
      patterns[31627] = 25'b01111011_10001001_00000100_1;
      patterns[31628] = 25'b01111011_10001010_00000101_1;
      patterns[31629] = 25'b01111011_10001011_00000110_1;
      patterns[31630] = 25'b01111011_10001100_00000111_1;
      patterns[31631] = 25'b01111011_10001101_00001000_1;
      patterns[31632] = 25'b01111011_10001110_00001001_1;
      patterns[31633] = 25'b01111011_10001111_00001010_1;
      patterns[31634] = 25'b01111011_10010000_00001011_1;
      patterns[31635] = 25'b01111011_10010001_00001100_1;
      patterns[31636] = 25'b01111011_10010010_00001101_1;
      patterns[31637] = 25'b01111011_10010011_00001110_1;
      patterns[31638] = 25'b01111011_10010100_00001111_1;
      patterns[31639] = 25'b01111011_10010101_00010000_1;
      patterns[31640] = 25'b01111011_10010110_00010001_1;
      patterns[31641] = 25'b01111011_10010111_00010010_1;
      patterns[31642] = 25'b01111011_10011000_00010011_1;
      patterns[31643] = 25'b01111011_10011001_00010100_1;
      patterns[31644] = 25'b01111011_10011010_00010101_1;
      patterns[31645] = 25'b01111011_10011011_00010110_1;
      patterns[31646] = 25'b01111011_10011100_00010111_1;
      patterns[31647] = 25'b01111011_10011101_00011000_1;
      patterns[31648] = 25'b01111011_10011110_00011001_1;
      patterns[31649] = 25'b01111011_10011111_00011010_1;
      patterns[31650] = 25'b01111011_10100000_00011011_1;
      patterns[31651] = 25'b01111011_10100001_00011100_1;
      patterns[31652] = 25'b01111011_10100010_00011101_1;
      patterns[31653] = 25'b01111011_10100011_00011110_1;
      patterns[31654] = 25'b01111011_10100100_00011111_1;
      patterns[31655] = 25'b01111011_10100101_00100000_1;
      patterns[31656] = 25'b01111011_10100110_00100001_1;
      patterns[31657] = 25'b01111011_10100111_00100010_1;
      patterns[31658] = 25'b01111011_10101000_00100011_1;
      patterns[31659] = 25'b01111011_10101001_00100100_1;
      patterns[31660] = 25'b01111011_10101010_00100101_1;
      patterns[31661] = 25'b01111011_10101011_00100110_1;
      patterns[31662] = 25'b01111011_10101100_00100111_1;
      patterns[31663] = 25'b01111011_10101101_00101000_1;
      patterns[31664] = 25'b01111011_10101110_00101001_1;
      patterns[31665] = 25'b01111011_10101111_00101010_1;
      patterns[31666] = 25'b01111011_10110000_00101011_1;
      patterns[31667] = 25'b01111011_10110001_00101100_1;
      patterns[31668] = 25'b01111011_10110010_00101101_1;
      patterns[31669] = 25'b01111011_10110011_00101110_1;
      patterns[31670] = 25'b01111011_10110100_00101111_1;
      patterns[31671] = 25'b01111011_10110101_00110000_1;
      patterns[31672] = 25'b01111011_10110110_00110001_1;
      patterns[31673] = 25'b01111011_10110111_00110010_1;
      patterns[31674] = 25'b01111011_10111000_00110011_1;
      patterns[31675] = 25'b01111011_10111001_00110100_1;
      patterns[31676] = 25'b01111011_10111010_00110101_1;
      patterns[31677] = 25'b01111011_10111011_00110110_1;
      patterns[31678] = 25'b01111011_10111100_00110111_1;
      patterns[31679] = 25'b01111011_10111101_00111000_1;
      patterns[31680] = 25'b01111011_10111110_00111001_1;
      patterns[31681] = 25'b01111011_10111111_00111010_1;
      patterns[31682] = 25'b01111011_11000000_00111011_1;
      patterns[31683] = 25'b01111011_11000001_00111100_1;
      patterns[31684] = 25'b01111011_11000010_00111101_1;
      patterns[31685] = 25'b01111011_11000011_00111110_1;
      patterns[31686] = 25'b01111011_11000100_00111111_1;
      patterns[31687] = 25'b01111011_11000101_01000000_1;
      patterns[31688] = 25'b01111011_11000110_01000001_1;
      patterns[31689] = 25'b01111011_11000111_01000010_1;
      patterns[31690] = 25'b01111011_11001000_01000011_1;
      patterns[31691] = 25'b01111011_11001001_01000100_1;
      patterns[31692] = 25'b01111011_11001010_01000101_1;
      patterns[31693] = 25'b01111011_11001011_01000110_1;
      patterns[31694] = 25'b01111011_11001100_01000111_1;
      patterns[31695] = 25'b01111011_11001101_01001000_1;
      patterns[31696] = 25'b01111011_11001110_01001001_1;
      patterns[31697] = 25'b01111011_11001111_01001010_1;
      patterns[31698] = 25'b01111011_11010000_01001011_1;
      patterns[31699] = 25'b01111011_11010001_01001100_1;
      patterns[31700] = 25'b01111011_11010010_01001101_1;
      patterns[31701] = 25'b01111011_11010011_01001110_1;
      patterns[31702] = 25'b01111011_11010100_01001111_1;
      patterns[31703] = 25'b01111011_11010101_01010000_1;
      patterns[31704] = 25'b01111011_11010110_01010001_1;
      patterns[31705] = 25'b01111011_11010111_01010010_1;
      patterns[31706] = 25'b01111011_11011000_01010011_1;
      patterns[31707] = 25'b01111011_11011001_01010100_1;
      patterns[31708] = 25'b01111011_11011010_01010101_1;
      patterns[31709] = 25'b01111011_11011011_01010110_1;
      patterns[31710] = 25'b01111011_11011100_01010111_1;
      patterns[31711] = 25'b01111011_11011101_01011000_1;
      patterns[31712] = 25'b01111011_11011110_01011001_1;
      patterns[31713] = 25'b01111011_11011111_01011010_1;
      patterns[31714] = 25'b01111011_11100000_01011011_1;
      patterns[31715] = 25'b01111011_11100001_01011100_1;
      patterns[31716] = 25'b01111011_11100010_01011101_1;
      patterns[31717] = 25'b01111011_11100011_01011110_1;
      patterns[31718] = 25'b01111011_11100100_01011111_1;
      patterns[31719] = 25'b01111011_11100101_01100000_1;
      patterns[31720] = 25'b01111011_11100110_01100001_1;
      patterns[31721] = 25'b01111011_11100111_01100010_1;
      patterns[31722] = 25'b01111011_11101000_01100011_1;
      patterns[31723] = 25'b01111011_11101001_01100100_1;
      patterns[31724] = 25'b01111011_11101010_01100101_1;
      patterns[31725] = 25'b01111011_11101011_01100110_1;
      patterns[31726] = 25'b01111011_11101100_01100111_1;
      patterns[31727] = 25'b01111011_11101101_01101000_1;
      patterns[31728] = 25'b01111011_11101110_01101001_1;
      patterns[31729] = 25'b01111011_11101111_01101010_1;
      patterns[31730] = 25'b01111011_11110000_01101011_1;
      patterns[31731] = 25'b01111011_11110001_01101100_1;
      patterns[31732] = 25'b01111011_11110010_01101101_1;
      patterns[31733] = 25'b01111011_11110011_01101110_1;
      patterns[31734] = 25'b01111011_11110100_01101111_1;
      patterns[31735] = 25'b01111011_11110101_01110000_1;
      patterns[31736] = 25'b01111011_11110110_01110001_1;
      patterns[31737] = 25'b01111011_11110111_01110010_1;
      patterns[31738] = 25'b01111011_11111000_01110011_1;
      patterns[31739] = 25'b01111011_11111001_01110100_1;
      patterns[31740] = 25'b01111011_11111010_01110101_1;
      patterns[31741] = 25'b01111011_11111011_01110110_1;
      patterns[31742] = 25'b01111011_11111100_01110111_1;
      patterns[31743] = 25'b01111011_11111101_01111000_1;
      patterns[31744] = 25'b01111011_11111110_01111001_1;
      patterns[31745] = 25'b01111011_11111111_01111010_1;
      patterns[31746] = 25'b01111100_00000000_01111100_0;
      patterns[31747] = 25'b01111100_00000001_01111101_0;
      patterns[31748] = 25'b01111100_00000010_01111110_0;
      patterns[31749] = 25'b01111100_00000011_01111111_0;
      patterns[31750] = 25'b01111100_00000100_10000000_0;
      patterns[31751] = 25'b01111100_00000101_10000001_0;
      patterns[31752] = 25'b01111100_00000110_10000010_0;
      patterns[31753] = 25'b01111100_00000111_10000011_0;
      patterns[31754] = 25'b01111100_00001000_10000100_0;
      patterns[31755] = 25'b01111100_00001001_10000101_0;
      patterns[31756] = 25'b01111100_00001010_10000110_0;
      patterns[31757] = 25'b01111100_00001011_10000111_0;
      patterns[31758] = 25'b01111100_00001100_10001000_0;
      patterns[31759] = 25'b01111100_00001101_10001001_0;
      patterns[31760] = 25'b01111100_00001110_10001010_0;
      patterns[31761] = 25'b01111100_00001111_10001011_0;
      patterns[31762] = 25'b01111100_00010000_10001100_0;
      patterns[31763] = 25'b01111100_00010001_10001101_0;
      patterns[31764] = 25'b01111100_00010010_10001110_0;
      patterns[31765] = 25'b01111100_00010011_10001111_0;
      patterns[31766] = 25'b01111100_00010100_10010000_0;
      patterns[31767] = 25'b01111100_00010101_10010001_0;
      patterns[31768] = 25'b01111100_00010110_10010010_0;
      patterns[31769] = 25'b01111100_00010111_10010011_0;
      patterns[31770] = 25'b01111100_00011000_10010100_0;
      patterns[31771] = 25'b01111100_00011001_10010101_0;
      patterns[31772] = 25'b01111100_00011010_10010110_0;
      patterns[31773] = 25'b01111100_00011011_10010111_0;
      patterns[31774] = 25'b01111100_00011100_10011000_0;
      patterns[31775] = 25'b01111100_00011101_10011001_0;
      patterns[31776] = 25'b01111100_00011110_10011010_0;
      patterns[31777] = 25'b01111100_00011111_10011011_0;
      patterns[31778] = 25'b01111100_00100000_10011100_0;
      patterns[31779] = 25'b01111100_00100001_10011101_0;
      patterns[31780] = 25'b01111100_00100010_10011110_0;
      patterns[31781] = 25'b01111100_00100011_10011111_0;
      patterns[31782] = 25'b01111100_00100100_10100000_0;
      patterns[31783] = 25'b01111100_00100101_10100001_0;
      patterns[31784] = 25'b01111100_00100110_10100010_0;
      patterns[31785] = 25'b01111100_00100111_10100011_0;
      patterns[31786] = 25'b01111100_00101000_10100100_0;
      patterns[31787] = 25'b01111100_00101001_10100101_0;
      patterns[31788] = 25'b01111100_00101010_10100110_0;
      patterns[31789] = 25'b01111100_00101011_10100111_0;
      patterns[31790] = 25'b01111100_00101100_10101000_0;
      patterns[31791] = 25'b01111100_00101101_10101001_0;
      patterns[31792] = 25'b01111100_00101110_10101010_0;
      patterns[31793] = 25'b01111100_00101111_10101011_0;
      patterns[31794] = 25'b01111100_00110000_10101100_0;
      patterns[31795] = 25'b01111100_00110001_10101101_0;
      patterns[31796] = 25'b01111100_00110010_10101110_0;
      patterns[31797] = 25'b01111100_00110011_10101111_0;
      patterns[31798] = 25'b01111100_00110100_10110000_0;
      patterns[31799] = 25'b01111100_00110101_10110001_0;
      patterns[31800] = 25'b01111100_00110110_10110010_0;
      patterns[31801] = 25'b01111100_00110111_10110011_0;
      patterns[31802] = 25'b01111100_00111000_10110100_0;
      patterns[31803] = 25'b01111100_00111001_10110101_0;
      patterns[31804] = 25'b01111100_00111010_10110110_0;
      patterns[31805] = 25'b01111100_00111011_10110111_0;
      patterns[31806] = 25'b01111100_00111100_10111000_0;
      patterns[31807] = 25'b01111100_00111101_10111001_0;
      patterns[31808] = 25'b01111100_00111110_10111010_0;
      patterns[31809] = 25'b01111100_00111111_10111011_0;
      patterns[31810] = 25'b01111100_01000000_10111100_0;
      patterns[31811] = 25'b01111100_01000001_10111101_0;
      patterns[31812] = 25'b01111100_01000010_10111110_0;
      patterns[31813] = 25'b01111100_01000011_10111111_0;
      patterns[31814] = 25'b01111100_01000100_11000000_0;
      patterns[31815] = 25'b01111100_01000101_11000001_0;
      patterns[31816] = 25'b01111100_01000110_11000010_0;
      patterns[31817] = 25'b01111100_01000111_11000011_0;
      patterns[31818] = 25'b01111100_01001000_11000100_0;
      patterns[31819] = 25'b01111100_01001001_11000101_0;
      patterns[31820] = 25'b01111100_01001010_11000110_0;
      patterns[31821] = 25'b01111100_01001011_11000111_0;
      patterns[31822] = 25'b01111100_01001100_11001000_0;
      patterns[31823] = 25'b01111100_01001101_11001001_0;
      patterns[31824] = 25'b01111100_01001110_11001010_0;
      patterns[31825] = 25'b01111100_01001111_11001011_0;
      patterns[31826] = 25'b01111100_01010000_11001100_0;
      patterns[31827] = 25'b01111100_01010001_11001101_0;
      patterns[31828] = 25'b01111100_01010010_11001110_0;
      patterns[31829] = 25'b01111100_01010011_11001111_0;
      patterns[31830] = 25'b01111100_01010100_11010000_0;
      patterns[31831] = 25'b01111100_01010101_11010001_0;
      patterns[31832] = 25'b01111100_01010110_11010010_0;
      patterns[31833] = 25'b01111100_01010111_11010011_0;
      patterns[31834] = 25'b01111100_01011000_11010100_0;
      patterns[31835] = 25'b01111100_01011001_11010101_0;
      patterns[31836] = 25'b01111100_01011010_11010110_0;
      patterns[31837] = 25'b01111100_01011011_11010111_0;
      patterns[31838] = 25'b01111100_01011100_11011000_0;
      patterns[31839] = 25'b01111100_01011101_11011001_0;
      patterns[31840] = 25'b01111100_01011110_11011010_0;
      patterns[31841] = 25'b01111100_01011111_11011011_0;
      patterns[31842] = 25'b01111100_01100000_11011100_0;
      patterns[31843] = 25'b01111100_01100001_11011101_0;
      patterns[31844] = 25'b01111100_01100010_11011110_0;
      patterns[31845] = 25'b01111100_01100011_11011111_0;
      patterns[31846] = 25'b01111100_01100100_11100000_0;
      patterns[31847] = 25'b01111100_01100101_11100001_0;
      patterns[31848] = 25'b01111100_01100110_11100010_0;
      patterns[31849] = 25'b01111100_01100111_11100011_0;
      patterns[31850] = 25'b01111100_01101000_11100100_0;
      patterns[31851] = 25'b01111100_01101001_11100101_0;
      patterns[31852] = 25'b01111100_01101010_11100110_0;
      patterns[31853] = 25'b01111100_01101011_11100111_0;
      patterns[31854] = 25'b01111100_01101100_11101000_0;
      patterns[31855] = 25'b01111100_01101101_11101001_0;
      patterns[31856] = 25'b01111100_01101110_11101010_0;
      patterns[31857] = 25'b01111100_01101111_11101011_0;
      patterns[31858] = 25'b01111100_01110000_11101100_0;
      patterns[31859] = 25'b01111100_01110001_11101101_0;
      patterns[31860] = 25'b01111100_01110010_11101110_0;
      patterns[31861] = 25'b01111100_01110011_11101111_0;
      patterns[31862] = 25'b01111100_01110100_11110000_0;
      patterns[31863] = 25'b01111100_01110101_11110001_0;
      patterns[31864] = 25'b01111100_01110110_11110010_0;
      patterns[31865] = 25'b01111100_01110111_11110011_0;
      patterns[31866] = 25'b01111100_01111000_11110100_0;
      patterns[31867] = 25'b01111100_01111001_11110101_0;
      patterns[31868] = 25'b01111100_01111010_11110110_0;
      patterns[31869] = 25'b01111100_01111011_11110111_0;
      patterns[31870] = 25'b01111100_01111100_11111000_0;
      patterns[31871] = 25'b01111100_01111101_11111001_0;
      patterns[31872] = 25'b01111100_01111110_11111010_0;
      patterns[31873] = 25'b01111100_01111111_11111011_0;
      patterns[31874] = 25'b01111100_10000000_11111100_0;
      patterns[31875] = 25'b01111100_10000001_11111101_0;
      patterns[31876] = 25'b01111100_10000010_11111110_0;
      patterns[31877] = 25'b01111100_10000011_11111111_0;
      patterns[31878] = 25'b01111100_10000100_00000000_1;
      patterns[31879] = 25'b01111100_10000101_00000001_1;
      patterns[31880] = 25'b01111100_10000110_00000010_1;
      patterns[31881] = 25'b01111100_10000111_00000011_1;
      patterns[31882] = 25'b01111100_10001000_00000100_1;
      patterns[31883] = 25'b01111100_10001001_00000101_1;
      patterns[31884] = 25'b01111100_10001010_00000110_1;
      patterns[31885] = 25'b01111100_10001011_00000111_1;
      patterns[31886] = 25'b01111100_10001100_00001000_1;
      patterns[31887] = 25'b01111100_10001101_00001001_1;
      patterns[31888] = 25'b01111100_10001110_00001010_1;
      patterns[31889] = 25'b01111100_10001111_00001011_1;
      patterns[31890] = 25'b01111100_10010000_00001100_1;
      patterns[31891] = 25'b01111100_10010001_00001101_1;
      patterns[31892] = 25'b01111100_10010010_00001110_1;
      patterns[31893] = 25'b01111100_10010011_00001111_1;
      patterns[31894] = 25'b01111100_10010100_00010000_1;
      patterns[31895] = 25'b01111100_10010101_00010001_1;
      patterns[31896] = 25'b01111100_10010110_00010010_1;
      patterns[31897] = 25'b01111100_10010111_00010011_1;
      patterns[31898] = 25'b01111100_10011000_00010100_1;
      patterns[31899] = 25'b01111100_10011001_00010101_1;
      patterns[31900] = 25'b01111100_10011010_00010110_1;
      patterns[31901] = 25'b01111100_10011011_00010111_1;
      patterns[31902] = 25'b01111100_10011100_00011000_1;
      patterns[31903] = 25'b01111100_10011101_00011001_1;
      patterns[31904] = 25'b01111100_10011110_00011010_1;
      patterns[31905] = 25'b01111100_10011111_00011011_1;
      patterns[31906] = 25'b01111100_10100000_00011100_1;
      patterns[31907] = 25'b01111100_10100001_00011101_1;
      patterns[31908] = 25'b01111100_10100010_00011110_1;
      patterns[31909] = 25'b01111100_10100011_00011111_1;
      patterns[31910] = 25'b01111100_10100100_00100000_1;
      patterns[31911] = 25'b01111100_10100101_00100001_1;
      patterns[31912] = 25'b01111100_10100110_00100010_1;
      patterns[31913] = 25'b01111100_10100111_00100011_1;
      patterns[31914] = 25'b01111100_10101000_00100100_1;
      patterns[31915] = 25'b01111100_10101001_00100101_1;
      patterns[31916] = 25'b01111100_10101010_00100110_1;
      patterns[31917] = 25'b01111100_10101011_00100111_1;
      patterns[31918] = 25'b01111100_10101100_00101000_1;
      patterns[31919] = 25'b01111100_10101101_00101001_1;
      patterns[31920] = 25'b01111100_10101110_00101010_1;
      patterns[31921] = 25'b01111100_10101111_00101011_1;
      patterns[31922] = 25'b01111100_10110000_00101100_1;
      patterns[31923] = 25'b01111100_10110001_00101101_1;
      patterns[31924] = 25'b01111100_10110010_00101110_1;
      patterns[31925] = 25'b01111100_10110011_00101111_1;
      patterns[31926] = 25'b01111100_10110100_00110000_1;
      patterns[31927] = 25'b01111100_10110101_00110001_1;
      patterns[31928] = 25'b01111100_10110110_00110010_1;
      patterns[31929] = 25'b01111100_10110111_00110011_1;
      patterns[31930] = 25'b01111100_10111000_00110100_1;
      patterns[31931] = 25'b01111100_10111001_00110101_1;
      patterns[31932] = 25'b01111100_10111010_00110110_1;
      patterns[31933] = 25'b01111100_10111011_00110111_1;
      patterns[31934] = 25'b01111100_10111100_00111000_1;
      patterns[31935] = 25'b01111100_10111101_00111001_1;
      patterns[31936] = 25'b01111100_10111110_00111010_1;
      patterns[31937] = 25'b01111100_10111111_00111011_1;
      patterns[31938] = 25'b01111100_11000000_00111100_1;
      patterns[31939] = 25'b01111100_11000001_00111101_1;
      patterns[31940] = 25'b01111100_11000010_00111110_1;
      patterns[31941] = 25'b01111100_11000011_00111111_1;
      patterns[31942] = 25'b01111100_11000100_01000000_1;
      patterns[31943] = 25'b01111100_11000101_01000001_1;
      patterns[31944] = 25'b01111100_11000110_01000010_1;
      patterns[31945] = 25'b01111100_11000111_01000011_1;
      patterns[31946] = 25'b01111100_11001000_01000100_1;
      patterns[31947] = 25'b01111100_11001001_01000101_1;
      patterns[31948] = 25'b01111100_11001010_01000110_1;
      patterns[31949] = 25'b01111100_11001011_01000111_1;
      patterns[31950] = 25'b01111100_11001100_01001000_1;
      patterns[31951] = 25'b01111100_11001101_01001001_1;
      patterns[31952] = 25'b01111100_11001110_01001010_1;
      patterns[31953] = 25'b01111100_11001111_01001011_1;
      patterns[31954] = 25'b01111100_11010000_01001100_1;
      patterns[31955] = 25'b01111100_11010001_01001101_1;
      patterns[31956] = 25'b01111100_11010010_01001110_1;
      patterns[31957] = 25'b01111100_11010011_01001111_1;
      patterns[31958] = 25'b01111100_11010100_01010000_1;
      patterns[31959] = 25'b01111100_11010101_01010001_1;
      patterns[31960] = 25'b01111100_11010110_01010010_1;
      patterns[31961] = 25'b01111100_11010111_01010011_1;
      patterns[31962] = 25'b01111100_11011000_01010100_1;
      patterns[31963] = 25'b01111100_11011001_01010101_1;
      patterns[31964] = 25'b01111100_11011010_01010110_1;
      patterns[31965] = 25'b01111100_11011011_01010111_1;
      patterns[31966] = 25'b01111100_11011100_01011000_1;
      patterns[31967] = 25'b01111100_11011101_01011001_1;
      patterns[31968] = 25'b01111100_11011110_01011010_1;
      patterns[31969] = 25'b01111100_11011111_01011011_1;
      patterns[31970] = 25'b01111100_11100000_01011100_1;
      patterns[31971] = 25'b01111100_11100001_01011101_1;
      patterns[31972] = 25'b01111100_11100010_01011110_1;
      patterns[31973] = 25'b01111100_11100011_01011111_1;
      patterns[31974] = 25'b01111100_11100100_01100000_1;
      patterns[31975] = 25'b01111100_11100101_01100001_1;
      patterns[31976] = 25'b01111100_11100110_01100010_1;
      patterns[31977] = 25'b01111100_11100111_01100011_1;
      patterns[31978] = 25'b01111100_11101000_01100100_1;
      patterns[31979] = 25'b01111100_11101001_01100101_1;
      patterns[31980] = 25'b01111100_11101010_01100110_1;
      patterns[31981] = 25'b01111100_11101011_01100111_1;
      patterns[31982] = 25'b01111100_11101100_01101000_1;
      patterns[31983] = 25'b01111100_11101101_01101001_1;
      patterns[31984] = 25'b01111100_11101110_01101010_1;
      patterns[31985] = 25'b01111100_11101111_01101011_1;
      patterns[31986] = 25'b01111100_11110000_01101100_1;
      patterns[31987] = 25'b01111100_11110001_01101101_1;
      patterns[31988] = 25'b01111100_11110010_01101110_1;
      patterns[31989] = 25'b01111100_11110011_01101111_1;
      patterns[31990] = 25'b01111100_11110100_01110000_1;
      patterns[31991] = 25'b01111100_11110101_01110001_1;
      patterns[31992] = 25'b01111100_11110110_01110010_1;
      patterns[31993] = 25'b01111100_11110111_01110011_1;
      patterns[31994] = 25'b01111100_11111000_01110100_1;
      patterns[31995] = 25'b01111100_11111001_01110101_1;
      patterns[31996] = 25'b01111100_11111010_01110110_1;
      patterns[31997] = 25'b01111100_11111011_01110111_1;
      patterns[31998] = 25'b01111100_11111100_01111000_1;
      patterns[31999] = 25'b01111100_11111101_01111001_1;
      patterns[32000] = 25'b01111100_11111110_01111010_1;
      patterns[32001] = 25'b01111100_11111111_01111011_1;
      patterns[32002] = 25'b01111101_00000000_01111101_0;
      patterns[32003] = 25'b01111101_00000001_01111110_0;
      patterns[32004] = 25'b01111101_00000010_01111111_0;
      patterns[32005] = 25'b01111101_00000011_10000000_0;
      patterns[32006] = 25'b01111101_00000100_10000001_0;
      patterns[32007] = 25'b01111101_00000101_10000010_0;
      patterns[32008] = 25'b01111101_00000110_10000011_0;
      patterns[32009] = 25'b01111101_00000111_10000100_0;
      patterns[32010] = 25'b01111101_00001000_10000101_0;
      patterns[32011] = 25'b01111101_00001001_10000110_0;
      patterns[32012] = 25'b01111101_00001010_10000111_0;
      patterns[32013] = 25'b01111101_00001011_10001000_0;
      patterns[32014] = 25'b01111101_00001100_10001001_0;
      patterns[32015] = 25'b01111101_00001101_10001010_0;
      patterns[32016] = 25'b01111101_00001110_10001011_0;
      patterns[32017] = 25'b01111101_00001111_10001100_0;
      patterns[32018] = 25'b01111101_00010000_10001101_0;
      patterns[32019] = 25'b01111101_00010001_10001110_0;
      patterns[32020] = 25'b01111101_00010010_10001111_0;
      patterns[32021] = 25'b01111101_00010011_10010000_0;
      patterns[32022] = 25'b01111101_00010100_10010001_0;
      patterns[32023] = 25'b01111101_00010101_10010010_0;
      patterns[32024] = 25'b01111101_00010110_10010011_0;
      patterns[32025] = 25'b01111101_00010111_10010100_0;
      patterns[32026] = 25'b01111101_00011000_10010101_0;
      patterns[32027] = 25'b01111101_00011001_10010110_0;
      patterns[32028] = 25'b01111101_00011010_10010111_0;
      patterns[32029] = 25'b01111101_00011011_10011000_0;
      patterns[32030] = 25'b01111101_00011100_10011001_0;
      patterns[32031] = 25'b01111101_00011101_10011010_0;
      patterns[32032] = 25'b01111101_00011110_10011011_0;
      patterns[32033] = 25'b01111101_00011111_10011100_0;
      patterns[32034] = 25'b01111101_00100000_10011101_0;
      patterns[32035] = 25'b01111101_00100001_10011110_0;
      patterns[32036] = 25'b01111101_00100010_10011111_0;
      patterns[32037] = 25'b01111101_00100011_10100000_0;
      patterns[32038] = 25'b01111101_00100100_10100001_0;
      patterns[32039] = 25'b01111101_00100101_10100010_0;
      patterns[32040] = 25'b01111101_00100110_10100011_0;
      patterns[32041] = 25'b01111101_00100111_10100100_0;
      patterns[32042] = 25'b01111101_00101000_10100101_0;
      patterns[32043] = 25'b01111101_00101001_10100110_0;
      patterns[32044] = 25'b01111101_00101010_10100111_0;
      patterns[32045] = 25'b01111101_00101011_10101000_0;
      patterns[32046] = 25'b01111101_00101100_10101001_0;
      patterns[32047] = 25'b01111101_00101101_10101010_0;
      patterns[32048] = 25'b01111101_00101110_10101011_0;
      patterns[32049] = 25'b01111101_00101111_10101100_0;
      patterns[32050] = 25'b01111101_00110000_10101101_0;
      patterns[32051] = 25'b01111101_00110001_10101110_0;
      patterns[32052] = 25'b01111101_00110010_10101111_0;
      patterns[32053] = 25'b01111101_00110011_10110000_0;
      patterns[32054] = 25'b01111101_00110100_10110001_0;
      patterns[32055] = 25'b01111101_00110101_10110010_0;
      patterns[32056] = 25'b01111101_00110110_10110011_0;
      patterns[32057] = 25'b01111101_00110111_10110100_0;
      patterns[32058] = 25'b01111101_00111000_10110101_0;
      patterns[32059] = 25'b01111101_00111001_10110110_0;
      patterns[32060] = 25'b01111101_00111010_10110111_0;
      patterns[32061] = 25'b01111101_00111011_10111000_0;
      patterns[32062] = 25'b01111101_00111100_10111001_0;
      patterns[32063] = 25'b01111101_00111101_10111010_0;
      patterns[32064] = 25'b01111101_00111110_10111011_0;
      patterns[32065] = 25'b01111101_00111111_10111100_0;
      patterns[32066] = 25'b01111101_01000000_10111101_0;
      patterns[32067] = 25'b01111101_01000001_10111110_0;
      patterns[32068] = 25'b01111101_01000010_10111111_0;
      patterns[32069] = 25'b01111101_01000011_11000000_0;
      patterns[32070] = 25'b01111101_01000100_11000001_0;
      patterns[32071] = 25'b01111101_01000101_11000010_0;
      patterns[32072] = 25'b01111101_01000110_11000011_0;
      patterns[32073] = 25'b01111101_01000111_11000100_0;
      patterns[32074] = 25'b01111101_01001000_11000101_0;
      patterns[32075] = 25'b01111101_01001001_11000110_0;
      patterns[32076] = 25'b01111101_01001010_11000111_0;
      patterns[32077] = 25'b01111101_01001011_11001000_0;
      patterns[32078] = 25'b01111101_01001100_11001001_0;
      patterns[32079] = 25'b01111101_01001101_11001010_0;
      patterns[32080] = 25'b01111101_01001110_11001011_0;
      patterns[32081] = 25'b01111101_01001111_11001100_0;
      patterns[32082] = 25'b01111101_01010000_11001101_0;
      patterns[32083] = 25'b01111101_01010001_11001110_0;
      patterns[32084] = 25'b01111101_01010010_11001111_0;
      patterns[32085] = 25'b01111101_01010011_11010000_0;
      patterns[32086] = 25'b01111101_01010100_11010001_0;
      patterns[32087] = 25'b01111101_01010101_11010010_0;
      patterns[32088] = 25'b01111101_01010110_11010011_0;
      patterns[32089] = 25'b01111101_01010111_11010100_0;
      patterns[32090] = 25'b01111101_01011000_11010101_0;
      patterns[32091] = 25'b01111101_01011001_11010110_0;
      patterns[32092] = 25'b01111101_01011010_11010111_0;
      patterns[32093] = 25'b01111101_01011011_11011000_0;
      patterns[32094] = 25'b01111101_01011100_11011001_0;
      patterns[32095] = 25'b01111101_01011101_11011010_0;
      patterns[32096] = 25'b01111101_01011110_11011011_0;
      patterns[32097] = 25'b01111101_01011111_11011100_0;
      patterns[32098] = 25'b01111101_01100000_11011101_0;
      patterns[32099] = 25'b01111101_01100001_11011110_0;
      patterns[32100] = 25'b01111101_01100010_11011111_0;
      patterns[32101] = 25'b01111101_01100011_11100000_0;
      patterns[32102] = 25'b01111101_01100100_11100001_0;
      patterns[32103] = 25'b01111101_01100101_11100010_0;
      patterns[32104] = 25'b01111101_01100110_11100011_0;
      patterns[32105] = 25'b01111101_01100111_11100100_0;
      patterns[32106] = 25'b01111101_01101000_11100101_0;
      patterns[32107] = 25'b01111101_01101001_11100110_0;
      patterns[32108] = 25'b01111101_01101010_11100111_0;
      patterns[32109] = 25'b01111101_01101011_11101000_0;
      patterns[32110] = 25'b01111101_01101100_11101001_0;
      patterns[32111] = 25'b01111101_01101101_11101010_0;
      patterns[32112] = 25'b01111101_01101110_11101011_0;
      patterns[32113] = 25'b01111101_01101111_11101100_0;
      patterns[32114] = 25'b01111101_01110000_11101101_0;
      patterns[32115] = 25'b01111101_01110001_11101110_0;
      patterns[32116] = 25'b01111101_01110010_11101111_0;
      patterns[32117] = 25'b01111101_01110011_11110000_0;
      patterns[32118] = 25'b01111101_01110100_11110001_0;
      patterns[32119] = 25'b01111101_01110101_11110010_0;
      patterns[32120] = 25'b01111101_01110110_11110011_0;
      patterns[32121] = 25'b01111101_01110111_11110100_0;
      patterns[32122] = 25'b01111101_01111000_11110101_0;
      patterns[32123] = 25'b01111101_01111001_11110110_0;
      patterns[32124] = 25'b01111101_01111010_11110111_0;
      patterns[32125] = 25'b01111101_01111011_11111000_0;
      patterns[32126] = 25'b01111101_01111100_11111001_0;
      patterns[32127] = 25'b01111101_01111101_11111010_0;
      patterns[32128] = 25'b01111101_01111110_11111011_0;
      patterns[32129] = 25'b01111101_01111111_11111100_0;
      patterns[32130] = 25'b01111101_10000000_11111101_0;
      patterns[32131] = 25'b01111101_10000001_11111110_0;
      patterns[32132] = 25'b01111101_10000010_11111111_0;
      patterns[32133] = 25'b01111101_10000011_00000000_1;
      patterns[32134] = 25'b01111101_10000100_00000001_1;
      patterns[32135] = 25'b01111101_10000101_00000010_1;
      patterns[32136] = 25'b01111101_10000110_00000011_1;
      patterns[32137] = 25'b01111101_10000111_00000100_1;
      patterns[32138] = 25'b01111101_10001000_00000101_1;
      patterns[32139] = 25'b01111101_10001001_00000110_1;
      patterns[32140] = 25'b01111101_10001010_00000111_1;
      patterns[32141] = 25'b01111101_10001011_00001000_1;
      patterns[32142] = 25'b01111101_10001100_00001001_1;
      patterns[32143] = 25'b01111101_10001101_00001010_1;
      patterns[32144] = 25'b01111101_10001110_00001011_1;
      patterns[32145] = 25'b01111101_10001111_00001100_1;
      patterns[32146] = 25'b01111101_10010000_00001101_1;
      patterns[32147] = 25'b01111101_10010001_00001110_1;
      patterns[32148] = 25'b01111101_10010010_00001111_1;
      patterns[32149] = 25'b01111101_10010011_00010000_1;
      patterns[32150] = 25'b01111101_10010100_00010001_1;
      patterns[32151] = 25'b01111101_10010101_00010010_1;
      patterns[32152] = 25'b01111101_10010110_00010011_1;
      patterns[32153] = 25'b01111101_10010111_00010100_1;
      patterns[32154] = 25'b01111101_10011000_00010101_1;
      patterns[32155] = 25'b01111101_10011001_00010110_1;
      patterns[32156] = 25'b01111101_10011010_00010111_1;
      patterns[32157] = 25'b01111101_10011011_00011000_1;
      patterns[32158] = 25'b01111101_10011100_00011001_1;
      patterns[32159] = 25'b01111101_10011101_00011010_1;
      patterns[32160] = 25'b01111101_10011110_00011011_1;
      patterns[32161] = 25'b01111101_10011111_00011100_1;
      patterns[32162] = 25'b01111101_10100000_00011101_1;
      patterns[32163] = 25'b01111101_10100001_00011110_1;
      patterns[32164] = 25'b01111101_10100010_00011111_1;
      patterns[32165] = 25'b01111101_10100011_00100000_1;
      patterns[32166] = 25'b01111101_10100100_00100001_1;
      patterns[32167] = 25'b01111101_10100101_00100010_1;
      patterns[32168] = 25'b01111101_10100110_00100011_1;
      patterns[32169] = 25'b01111101_10100111_00100100_1;
      patterns[32170] = 25'b01111101_10101000_00100101_1;
      patterns[32171] = 25'b01111101_10101001_00100110_1;
      patterns[32172] = 25'b01111101_10101010_00100111_1;
      patterns[32173] = 25'b01111101_10101011_00101000_1;
      patterns[32174] = 25'b01111101_10101100_00101001_1;
      patterns[32175] = 25'b01111101_10101101_00101010_1;
      patterns[32176] = 25'b01111101_10101110_00101011_1;
      patterns[32177] = 25'b01111101_10101111_00101100_1;
      patterns[32178] = 25'b01111101_10110000_00101101_1;
      patterns[32179] = 25'b01111101_10110001_00101110_1;
      patterns[32180] = 25'b01111101_10110010_00101111_1;
      patterns[32181] = 25'b01111101_10110011_00110000_1;
      patterns[32182] = 25'b01111101_10110100_00110001_1;
      patterns[32183] = 25'b01111101_10110101_00110010_1;
      patterns[32184] = 25'b01111101_10110110_00110011_1;
      patterns[32185] = 25'b01111101_10110111_00110100_1;
      patterns[32186] = 25'b01111101_10111000_00110101_1;
      patterns[32187] = 25'b01111101_10111001_00110110_1;
      patterns[32188] = 25'b01111101_10111010_00110111_1;
      patterns[32189] = 25'b01111101_10111011_00111000_1;
      patterns[32190] = 25'b01111101_10111100_00111001_1;
      patterns[32191] = 25'b01111101_10111101_00111010_1;
      patterns[32192] = 25'b01111101_10111110_00111011_1;
      patterns[32193] = 25'b01111101_10111111_00111100_1;
      patterns[32194] = 25'b01111101_11000000_00111101_1;
      patterns[32195] = 25'b01111101_11000001_00111110_1;
      patterns[32196] = 25'b01111101_11000010_00111111_1;
      patterns[32197] = 25'b01111101_11000011_01000000_1;
      patterns[32198] = 25'b01111101_11000100_01000001_1;
      patterns[32199] = 25'b01111101_11000101_01000010_1;
      patterns[32200] = 25'b01111101_11000110_01000011_1;
      patterns[32201] = 25'b01111101_11000111_01000100_1;
      patterns[32202] = 25'b01111101_11001000_01000101_1;
      patterns[32203] = 25'b01111101_11001001_01000110_1;
      patterns[32204] = 25'b01111101_11001010_01000111_1;
      patterns[32205] = 25'b01111101_11001011_01001000_1;
      patterns[32206] = 25'b01111101_11001100_01001001_1;
      patterns[32207] = 25'b01111101_11001101_01001010_1;
      patterns[32208] = 25'b01111101_11001110_01001011_1;
      patterns[32209] = 25'b01111101_11001111_01001100_1;
      patterns[32210] = 25'b01111101_11010000_01001101_1;
      patterns[32211] = 25'b01111101_11010001_01001110_1;
      patterns[32212] = 25'b01111101_11010010_01001111_1;
      patterns[32213] = 25'b01111101_11010011_01010000_1;
      patterns[32214] = 25'b01111101_11010100_01010001_1;
      patterns[32215] = 25'b01111101_11010101_01010010_1;
      patterns[32216] = 25'b01111101_11010110_01010011_1;
      patterns[32217] = 25'b01111101_11010111_01010100_1;
      patterns[32218] = 25'b01111101_11011000_01010101_1;
      patterns[32219] = 25'b01111101_11011001_01010110_1;
      patterns[32220] = 25'b01111101_11011010_01010111_1;
      patterns[32221] = 25'b01111101_11011011_01011000_1;
      patterns[32222] = 25'b01111101_11011100_01011001_1;
      patterns[32223] = 25'b01111101_11011101_01011010_1;
      patterns[32224] = 25'b01111101_11011110_01011011_1;
      patterns[32225] = 25'b01111101_11011111_01011100_1;
      patterns[32226] = 25'b01111101_11100000_01011101_1;
      patterns[32227] = 25'b01111101_11100001_01011110_1;
      patterns[32228] = 25'b01111101_11100010_01011111_1;
      patterns[32229] = 25'b01111101_11100011_01100000_1;
      patterns[32230] = 25'b01111101_11100100_01100001_1;
      patterns[32231] = 25'b01111101_11100101_01100010_1;
      patterns[32232] = 25'b01111101_11100110_01100011_1;
      patterns[32233] = 25'b01111101_11100111_01100100_1;
      patterns[32234] = 25'b01111101_11101000_01100101_1;
      patterns[32235] = 25'b01111101_11101001_01100110_1;
      patterns[32236] = 25'b01111101_11101010_01100111_1;
      patterns[32237] = 25'b01111101_11101011_01101000_1;
      patterns[32238] = 25'b01111101_11101100_01101001_1;
      patterns[32239] = 25'b01111101_11101101_01101010_1;
      patterns[32240] = 25'b01111101_11101110_01101011_1;
      patterns[32241] = 25'b01111101_11101111_01101100_1;
      patterns[32242] = 25'b01111101_11110000_01101101_1;
      patterns[32243] = 25'b01111101_11110001_01101110_1;
      patterns[32244] = 25'b01111101_11110010_01101111_1;
      patterns[32245] = 25'b01111101_11110011_01110000_1;
      patterns[32246] = 25'b01111101_11110100_01110001_1;
      patterns[32247] = 25'b01111101_11110101_01110010_1;
      patterns[32248] = 25'b01111101_11110110_01110011_1;
      patterns[32249] = 25'b01111101_11110111_01110100_1;
      patterns[32250] = 25'b01111101_11111000_01110101_1;
      patterns[32251] = 25'b01111101_11111001_01110110_1;
      patterns[32252] = 25'b01111101_11111010_01110111_1;
      patterns[32253] = 25'b01111101_11111011_01111000_1;
      patterns[32254] = 25'b01111101_11111100_01111001_1;
      patterns[32255] = 25'b01111101_11111101_01111010_1;
      patterns[32256] = 25'b01111101_11111110_01111011_1;
      patterns[32257] = 25'b01111101_11111111_01111100_1;
      patterns[32258] = 25'b01111110_00000000_01111110_0;
      patterns[32259] = 25'b01111110_00000001_01111111_0;
      patterns[32260] = 25'b01111110_00000010_10000000_0;
      patterns[32261] = 25'b01111110_00000011_10000001_0;
      patterns[32262] = 25'b01111110_00000100_10000010_0;
      patterns[32263] = 25'b01111110_00000101_10000011_0;
      patterns[32264] = 25'b01111110_00000110_10000100_0;
      patterns[32265] = 25'b01111110_00000111_10000101_0;
      patterns[32266] = 25'b01111110_00001000_10000110_0;
      patterns[32267] = 25'b01111110_00001001_10000111_0;
      patterns[32268] = 25'b01111110_00001010_10001000_0;
      patterns[32269] = 25'b01111110_00001011_10001001_0;
      patterns[32270] = 25'b01111110_00001100_10001010_0;
      patterns[32271] = 25'b01111110_00001101_10001011_0;
      patterns[32272] = 25'b01111110_00001110_10001100_0;
      patterns[32273] = 25'b01111110_00001111_10001101_0;
      patterns[32274] = 25'b01111110_00010000_10001110_0;
      patterns[32275] = 25'b01111110_00010001_10001111_0;
      patterns[32276] = 25'b01111110_00010010_10010000_0;
      patterns[32277] = 25'b01111110_00010011_10010001_0;
      patterns[32278] = 25'b01111110_00010100_10010010_0;
      patterns[32279] = 25'b01111110_00010101_10010011_0;
      patterns[32280] = 25'b01111110_00010110_10010100_0;
      patterns[32281] = 25'b01111110_00010111_10010101_0;
      patterns[32282] = 25'b01111110_00011000_10010110_0;
      patterns[32283] = 25'b01111110_00011001_10010111_0;
      patterns[32284] = 25'b01111110_00011010_10011000_0;
      patterns[32285] = 25'b01111110_00011011_10011001_0;
      patterns[32286] = 25'b01111110_00011100_10011010_0;
      patterns[32287] = 25'b01111110_00011101_10011011_0;
      patterns[32288] = 25'b01111110_00011110_10011100_0;
      patterns[32289] = 25'b01111110_00011111_10011101_0;
      patterns[32290] = 25'b01111110_00100000_10011110_0;
      patterns[32291] = 25'b01111110_00100001_10011111_0;
      patterns[32292] = 25'b01111110_00100010_10100000_0;
      patterns[32293] = 25'b01111110_00100011_10100001_0;
      patterns[32294] = 25'b01111110_00100100_10100010_0;
      patterns[32295] = 25'b01111110_00100101_10100011_0;
      patterns[32296] = 25'b01111110_00100110_10100100_0;
      patterns[32297] = 25'b01111110_00100111_10100101_0;
      patterns[32298] = 25'b01111110_00101000_10100110_0;
      patterns[32299] = 25'b01111110_00101001_10100111_0;
      patterns[32300] = 25'b01111110_00101010_10101000_0;
      patterns[32301] = 25'b01111110_00101011_10101001_0;
      patterns[32302] = 25'b01111110_00101100_10101010_0;
      patterns[32303] = 25'b01111110_00101101_10101011_0;
      patterns[32304] = 25'b01111110_00101110_10101100_0;
      patterns[32305] = 25'b01111110_00101111_10101101_0;
      patterns[32306] = 25'b01111110_00110000_10101110_0;
      patterns[32307] = 25'b01111110_00110001_10101111_0;
      patterns[32308] = 25'b01111110_00110010_10110000_0;
      patterns[32309] = 25'b01111110_00110011_10110001_0;
      patterns[32310] = 25'b01111110_00110100_10110010_0;
      patterns[32311] = 25'b01111110_00110101_10110011_0;
      patterns[32312] = 25'b01111110_00110110_10110100_0;
      patterns[32313] = 25'b01111110_00110111_10110101_0;
      patterns[32314] = 25'b01111110_00111000_10110110_0;
      patterns[32315] = 25'b01111110_00111001_10110111_0;
      patterns[32316] = 25'b01111110_00111010_10111000_0;
      patterns[32317] = 25'b01111110_00111011_10111001_0;
      patterns[32318] = 25'b01111110_00111100_10111010_0;
      patterns[32319] = 25'b01111110_00111101_10111011_0;
      patterns[32320] = 25'b01111110_00111110_10111100_0;
      patterns[32321] = 25'b01111110_00111111_10111101_0;
      patterns[32322] = 25'b01111110_01000000_10111110_0;
      patterns[32323] = 25'b01111110_01000001_10111111_0;
      patterns[32324] = 25'b01111110_01000010_11000000_0;
      patterns[32325] = 25'b01111110_01000011_11000001_0;
      patterns[32326] = 25'b01111110_01000100_11000010_0;
      patterns[32327] = 25'b01111110_01000101_11000011_0;
      patterns[32328] = 25'b01111110_01000110_11000100_0;
      patterns[32329] = 25'b01111110_01000111_11000101_0;
      patterns[32330] = 25'b01111110_01001000_11000110_0;
      patterns[32331] = 25'b01111110_01001001_11000111_0;
      patterns[32332] = 25'b01111110_01001010_11001000_0;
      patterns[32333] = 25'b01111110_01001011_11001001_0;
      patterns[32334] = 25'b01111110_01001100_11001010_0;
      patterns[32335] = 25'b01111110_01001101_11001011_0;
      patterns[32336] = 25'b01111110_01001110_11001100_0;
      patterns[32337] = 25'b01111110_01001111_11001101_0;
      patterns[32338] = 25'b01111110_01010000_11001110_0;
      patterns[32339] = 25'b01111110_01010001_11001111_0;
      patterns[32340] = 25'b01111110_01010010_11010000_0;
      patterns[32341] = 25'b01111110_01010011_11010001_0;
      patterns[32342] = 25'b01111110_01010100_11010010_0;
      patterns[32343] = 25'b01111110_01010101_11010011_0;
      patterns[32344] = 25'b01111110_01010110_11010100_0;
      patterns[32345] = 25'b01111110_01010111_11010101_0;
      patterns[32346] = 25'b01111110_01011000_11010110_0;
      patterns[32347] = 25'b01111110_01011001_11010111_0;
      patterns[32348] = 25'b01111110_01011010_11011000_0;
      patterns[32349] = 25'b01111110_01011011_11011001_0;
      patterns[32350] = 25'b01111110_01011100_11011010_0;
      patterns[32351] = 25'b01111110_01011101_11011011_0;
      patterns[32352] = 25'b01111110_01011110_11011100_0;
      patterns[32353] = 25'b01111110_01011111_11011101_0;
      patterns[32354] = 25'b01111110_01100000_11011110_0;
      patterns[32355] = 25'b01111110_01100001_11011111_0;
      patterns[32356] = 25'b01111110_01100010_11100000_0;
      patterns[32357] = 25'b01111110_01100011_11100001_0;
      patterns[32358] = 25'b01111110_01100100_11100010_0;
      patterns[32359] = 25'b01111110_01100101_11100011_0;
      patterns[32360] = 25'b01111110_01100110_11100100_0;
      patterns[32361] = 25'b01111110_01100111_11100101_0;
      patterns[32362] = 25'b01111110_01101000_11100110_0;
      patterns[32363] = 25'b01111110_01101001_11100111_0;
      patterns[32364] = 25'b01111110_01101010_11101000_0;
      patterns[32365] = 25'b01111110_01101011_11101001_0;
      patterns[32366] = 25'b01111110_01101100_11101010_0;
      patterns[32367] = 25'b01111110_01101101_11101011_0;
      patterns[32368] = 25'b01111110_01101110_11101100_0;
      patterns[32369] = 25'b01111110_01101111_11101101_0;
      patterns[32370] = 25'b01111110_01110000_11101110_0;
      patterns[32371] = 25'b01111110_01110001_11101111_0;
      patterns[32372] = 25'b01111110_01110010_11110000_0;
      patterns[32373] = 25'b01111110_01110011_11110001_0;
      patterns[32374] = 25'b01111110_01110100_11110010_0;
      patterns[32375] = 25'b01111110_01110101_11110011_0;
      patterns[32376] = 25'b01111110_01110110_11110100_0;
      patterns[32377] = 25'b01111110_01110111_11110101_0;
      patterns[32378] = 25'b01111110_01111000_11110110_0;
      patterns[32379] = 25'b01111110_01111001_11110111_0;
      patterns[32380] = 25'b01111110_01111010_11111000_0;
      patterns[32381] = 25'b01111110_01111011_11111001_0;
      patterns[32382] = 25'b01111110_01111100_11111010_0;
      patterns[32383] = 25'b01111110_01111101_11111011_0;
      patterns[32384] = 25'b01111110_01111110_11111100_0;
      patterns[32385] = 25'b01111110_01111111_11111101_0;
      patterns[32386] = 25'b01111110_10000000_11111110_0;
      patterns[32387] = 25'b01111110_10000001_11111111_0;
      patterns[32388] = 25'b01111110_10000010_00000000_1;
      patterns[32389] = 25'b01111110_10000011_00000001_1;
      patterns[32390] = 25'b01111110_10000100_00000010_1;
      patterns[32391] = 25'b01111110_10000101_00000011_1;
      patterns[32392] = 25'b01111110_10000110_00000100_1;
      patterns[32393] = 25'b01111110_10000111_00000101_1;
      patterns[32394] = 25'b01111110_10001000_00000110_1;
      patterns[32395] = 25'b01111110_10001001_00000111_1;
      patterns[32396] = 25'b01111110_10001010_00001000_1;
      patterns[32397] = 25'b01111110_10001011_00001001_1;
      patterns[32398] = 25'b01111110_10001100_00001010_1;
      patterns[32399] = 25'b01111110_10001101_00001011_1;
      patterns[32400] = 25'b01111110_10001110_00001100_1;
      patterns[32401] = 25'b01111110_10001111_00001101_1;
      patterns[32402] = 25'b01111110_10010000_00001110_1;
      patterns[32403] = 25'b01111110_10010001_00001111_1;
      patterns[32404] = 25'b01111110_10010010_00010000_1;
      patterns[32405] = 25'b01111110_10010011_00010001_1;
      patterns[32406] = 25'b01111110_10010100_00010010_1;
      patterns[32407] = 25'b01111110_10010101_00010011_1;
      patterns[32408] = 25'b01111110_10010110_00010100_1;
      patterns[32409] = 25'b01111110_10010111_00010101_1;
      patterns[32410] = 25'b01111110_10011000_00010110_1;
      patterns[32411] = 25'b01111110_10011001_00010111_1;
      patterns[32412] = 25'b01111110_10011010_00011000_1;
      patterns[32413] = 25'b01111110_10011011_00011001_1;
      patterns[32414] = 25'b01111110_10011100_00011010_1;
      patterns[32415] = 25'b01111110_10011101_00011011_1;
      patterns[32416] = 25'b01111110_10011110_00011100_1;
      patterns[32417] = 25'b01111110_10011111_00011101_1;
      patterns[32418] = 25'b01111110_10100000_00011110_1;
      patterns[32419] = 25'b01111110_10100001_00011111_1;
      patterns[32420] = 25'b01111110_10100010_00100000_1;
      patterns[32421] = 25'b01111110_10100011_00100001_1;
      patterns[32422] = 25'b01111110_10100100_00100010_1;
      patterns[32423] = 25'b01111110_10100101_00100011_1;
      patterns[32424] = 25'b01111110_10100110_00100100_1;
      patterns[32425] = 25'b01111110_10100111_00100101_1;
      patterns[32426] = 25'b01111110_10101000_00100110_1;
      patterns[32427] = 25'b01111110_10101001_00100111_1;
      patterns[32428] = 25'b01111110_10101010_00101000_1;
      patterns[32429] = 25'b01111110_10101011_00101001_1;
      patterns[32430] = 25'b01111110_10101100_00101010_1;
      patterns[32431] = 25'b01111110_10101101_00101011_1;
      patterns[32432] = 25'b01111110_10101110_00101100_1;
      patterns[32433] = 25'b01111110_10101111_00101101_1;
      patterns[32434] = 25'b01111110_10110000_00101110_1;
      patterns[32435] = 25'b01111110_10110001_00101111_1;
      patterns[32436] = 25'b01111110_10110010_00110000_1;
      patterns[32437] = 25'b01111110_10110011_00110001_1;
      patterns[32438] = 25'b01111110_10110100_00110010_1;
      patterns[32439] = 25'b01111110_10110101_00110011_1;
      patterns[32440] = 25'b01111110_10110110_00110100_1;
      patterns[32441] = 25'b01111110_10110111_00110101_1;
      patterns[32442] = 25'b01111110_10111000_00110110_1;
      patterns[32443] = 25'b01111110_10111001_00110111_1;
      patterns[32444] = 25'b01111110_10111010_00111000_1;
      patterns[32445] = 25'b01111110_10111011_00111001_1;
      patterns[32446] = 25'b01111110_10111100_00111010_1;
      patterns[32447] = 25'b01111110_10111101_00111011_1;
      patterns[32448] = 25'b01111110_10111110_00111100_1;
      patterns[32449] = 25'b01111110_10111111_00111101_1;
      patterns[32450] = 25'b01111110_11000000_00111110_1;
      patterns[32451] = 25'b01111110_11000001_00111111_1;
      patterns[32452] = 25'b01111110_11000010_01000000_1;
      patterns[32453] = 25'b01111110_11000011_01000001_1;
      patterns[32454] = 25'b01111110_11000100_01000010_1;
      patterns[32455] = 25'b01111110_11000101_01000011_1;
      patterns[32456] = 25'b01111110_11000110_01000100_1;
      patterns[32457] = 25'b01111110_11000111_01000101_1;
      patterns[32458] = 25'b01111110_11001000_01000110_1;
      patterns[32459] = 25'b01111110_11001001_01000111_1;
      patterns[32460] = 25'b01111110_11001010_01001000_1;
      patterns[32461] = 25'b01111110_11001011_01001001_1;
      patterns[32462] = 25'b01111110_11001100_01001010_1;
      patterns[32463] = 25'b01111110_11001101_01001011_1;
      patterns[32464] = 25'b01111110_11001110_01001100_1;
      patterns[32465] = 25'b01111110_11001111_01001101_1;
      patterns[32466] = 25'b01111110_11010000_01001110_1;
      patterns[32467] = 25'b01111110_11010001_01001111_1;
      patterns[32468] = 25'b01111110_11010010_01010000_1;
      patterns[32469] = 25'b01111110_11010011_01010001_1;
      patterns[32470] = 25'b01111110_11010100_01010010_1;
      patterns[32471] = 25'b01111110_11010101_01010011_1;
      patterns[32472] = 25'b01111110_11010110_01010100_1;
      patterns[32473] = 25'b01111110_11010111_01010101_1;
      patterns[32474] = 25'b01111110_11011000_01010110_1;
      patterns[32475] = 25'b01111110_11011001_01010111_1;
      patterns[32476] = 25'b01111110_11011010_01011000_1;
      patterns[32477] = 25'b01111110_11011011_01011001_1;
      patterns[32478] = 25'b01111110_11011100_01011010_1;
      patterns[32479] = 25'b01111110_11011101_01011011_1;
      patterns[32480] = 25'b01111110_11011110_01011100_1;
      patterns[32481] = 25'b01111110_11011111_01011101_1;
      patterns[32482] = 25'b01111110_11100000_01011110_1;
      patterns[32483] = 25'b01111110_11100001_01011111_1;
      patterns[32484] = 25'b01111110_11100010_01100000_1;
      patterns[32485] = 25'b01111110_11100011_01100001_1;
      patterns[32486] = 25'b01111110_11100100_01100010_1;
      patterns[32487] = 25'b01111110_11100101_01100011_1;
      patterns[32488] = 25'b01111110_11100110_01100100_1;
      patterns[32489] = 25'b01111110_11100111_01100101_1;
      patterns[32490] = 25'b01111110_11101000_01100110_1;
      patterns[32491] = 25'b01111110_11101001_01100111_1;
      patterns[32492] = 25'b01111110_11101010_01101000_1;
      patterns[32493] = 25'b01111110_11101011_01101001_1;
      patterns[32494] = 25'b01111110_11101100_01101010_1;
      patterns[32495] = 25'b01111110_11101101_01101011_1;
      patterns[32496] = 25'b01111110_11101110_01101100_1;
      patterns[32497] = 25'b01111110_11101111_01101101_1;
      patterns[32498] = 25'b01111110_11110000_01101110_1;
      patterns[32499] = 25'b01111110_11110001_01101111_1;
      patterns[32500] = 25'b01111110_11110010_01110000_1;
      patterns[32501] = 25'b01111110_11110011_01110001_1;
      patterns[32502] = 25'b01111110_11110100_01110010_1;
      patterns[32503] = 25'b01111110_11110101_01110011_1;
      patterns[32504] = 25'b01111110_11110110_01110100_1;
      patterns[32505] = 25'b01111110_11110111_01110101_1;
      patterns[32506] = 25'b01111110_11111000_01110110_1;
      patterns[32507] = 25'b01111110_11111001_01110111_1;
      patterns[32508] = 25'b01111110_11111010_01111000_1;
      patterns[32509] = 25'b01111110_11111011_01111001_1;
      patterns[32510] = 25'b01111110_11111100_01111010_1;
      patterns[32511] = 25'b01111110_11111101_01111011_1;
      patterns[32512] = 25'b01111110_11111110_01111100_1;
      patterns[32513] = 25'b01111110_11111111_01111101_1;
      patterns[32514] = 25'b01111111_00000000_01111111_0;
      patterns[32515] = 25'b01111111_00000001_10000000_0;
      patterns[32516] = 25'b01111111_00000010_10000001_0;
      patterns[32517] = 25'b01111111_00000011_10000010_0;
      patterns[32518] = 25'b01111111_00000100_10000011_0;
      patterns[32519] = 25'b01111111_00000101_10000100_0;
      patterns[32520] = 25'b01111111_00000110_10000101_0;
      patterns[32521] = 25'b01111111_00000111_10000110_0;
      patterns[32522] = 25'b01111111_00001000_10000111_0;
      patterns[32523] = 25'b01111111_00001001_10001000_0;
      patterns[32524] = 25'b01111111_00001010_10001001_0;
      patterns[32525] = 25'b01111111_00001011_10001010_0;
      patterns[32526] = 25'b01111111_00001100_10001011_0;
      patterns[32527] = 25'b01111111_00001101_10001100_0;
      patterns[32528] = 25'b01111111_00001110_10001101_0;
      patterns[32529] = 25'b01111111_00001111_10001110_0;
      patterns[32530] = 25'b01111111_00010000_10001111_0;
      patterns[32531] = 25'b01111111_00010001_10010000_0;
      patterns[32532] = 25'b01111111_00010010_10010001_0;
      patterns[32533] = 25'b01111111_00010011_10010010_0;
      patterns[32534] = 25'b01111111_00010100_10010011_0;
      patterns[32535] = 25'b01111111_00010101_10010100_0;
      patterns[32536] = 25'b01111111_00010110_10010101_0;
      patterns[32537] = 25'b01111111_00010111_10010110_0;
      patterns[32538] = 25'b01111111_00011000_10010111_0;
      patterns[32539] = 25'b01111111_00011001_10011000_0;
      patterns[32540] = 25'b01111111_00011010_10011001_0;
      patterns[32541] = 25'b01111111_00011011_10011010_0;
      patterns[32542] = 25'b01111111_00011100_10011011_0;
      patterns[32543] = 25'b01111111_00011101_10011100_0;
      patterns[32544] = 25'b01111111_00011110_10011101_0;
      patterns[32545] = 25'b01111111_00011111_10011110_0;
      patterns[32546] = 25'b01111111_00100000_10011111_0;
      patterns[32547] = 25'b01111111_00100001_10100000_0;
      patterns[32548] = 25'b01111111_00100010_10100001_0;
      patterns[32549] = 25'b01111111_00100011_10100010_0;
      patterns[32550] = 25'b01111111_00100100_10100011_0;
      patterns[32551] = 25'b01111111_00100101_10100100_0;
      patterns[32552] = 25'b01111111_00100110_10100101_0;
      patterns[32553] = 25'b01111111_00100111_10100110_0;
      patterns[32554] = 25'b01111111_00101000_10100111_0;
      patterns[32555] = 25'b01111111_00101001_10101000_0;
      patterns[32556] = 25'b01111111_00101010_10101001_0;
      patterns[32557] = 25'b01111111_00101011_10101010_0;
      patterns[32558] = 25'b01111111_00101100_10101011_0;
      patterns[32559] = 25'b01111111_00101101_10101100_0;
      patterns[32560] = 25'b01111111_00101110_10101101_0;
      patterns[32561] = 25'b01111111_00101111_10101110_0;
      patterns[32562] = 25'b01111111_00110000_10101111_0;
      patterns[32563] = 25'b01111111_00110001_10110000_0;
      patterns[32564] = 25'b01111111_00110010_10110001_0;
      patterns[32565] = 25'b01111111_00110011_10110010_0;
      patterns[32566] = 25'b01111111_00110100_10110011_0;
      patterns[32567] = 25'b01111111_00110101_10110100_0;
      patterns[32568] = 25'b01111111_00110110_10110101_0;
      patterns[32569] = 25'b01111111_00110111_10110110_0;
      patterns[32570] = 25'b01111111_00111000_10110111_0;
      patterns[32571] = 25'b01111111_00111001_10111000_0;
      patterns[32572] = 25'b01111111_00111010_10111001_0;
      patterns[32573] = 25'b01111111_00111011_10111010_0;
      patterns[32574] = 25'b01111111_00111100_10111011_0;
      patterns[32575] = 25'b01111111_00111101_10111100_0;
      patterns[32576] = 25'b01111111_00111110_10111101_0;
      patterns[32577] = 25'b01111111_00111111_10111110_0;
      patterns[32578] = 25'b01111111_01000000_10111111_0;
      patterns[32579] = 25'b01111111_01000001_11000000_0;
      patterns[32580] = 25'b01111111_01000010_11000001_0;
      patterns[32581] = 25'b01111111_01000011_11000010_0;
      patterns[32582] = 25'b01111111_01000100_11000011_0;
      patterns[32583] = 25'b01111111_01000101_11000100_0;
      patterns[32584] = 25'b01111111_01000110_11000101_0;
      patterns[32585] = 25'b01111111_01000111_11000110_0;
      patterns[32586] = 25'b01111111_01001000_11000111_0;
      patterns[32587] = 25'b01111111_01001001_11001000_0;
      patterns[32588] = 25'b01111111_01001010_11001001_0;
      patterns[32589] = 25'b01111111_01001011_11001010_0;
      patterns[32590] = 25'b01111111_01001100_11001011_0;
      patterns[32591] = 25'b01111111_01001101_11001100_0;
      patterns[32592] = 25'b01111111_01001110_11001101_0;
      patterns[32593] = 25'b01111111_01001111_11001110_0;
      patterns[32594] = 25'b01111111_01010000_11001111_0;
      patterns[32595] = 25'b01111111_01010001_11010000_0;
      patterns[32596] = 25'b01111111_01010010_11010001_0;
      patterns[32597] = 25'b01111111_01010011_11010010_0;
      patterns[32598] = 25'b01111111_01010100_11010011_0;
      patterns[32599] = 25'b01111111_01010101_11010100_0;
      patterns[32600] = 25'b01111111_01010110_11010101_0;
      patterns[32601] = 25'b01111111_01010111_11010110_0;
      patterns[32602] = 25'b01111111_01011000_11010111_0;
      patterns[32603] = 25'b01111111_01011001_11011000_0;
      patterns[32604] = 25'b01111111_01011010_11011001_0;
      patterns[32605] = 25'b01111111_01011011_11011010_0;
      patterns[32606] = 25'b01111111_01011100_11011011_0;
      patterns[32607] = 25'b01111111_01011101_11011100_0;
      patterns[32608] = 25'b01111111_01011110_11011101_0;
      patterns[32609] = 25'b01111111_01011111_11011110_0;
      patterns[32610] = 25'b01111111_01100000_11011111_0;
      patterns[32611] = 25'b01111111_01100001_11100000_0;
      patterns[32612] = 25'b01111111_01100010_11100001_0;
      patterns[32613] = 25'b01111111_01100011_11100010_0;
      patterns[32614] = 25'b01111111_01100100_11100011_0;
      patterns[32615] = 25'b01111111_01100101_11100100_0;
      patterns[32616] = 25'b01111111_01100110_11100101_0;
      patterns[32617] = 25'b01111111_01100111_11100110_0;
      patterns[32618] = 25'b01111111_01101000_11100111_0;
      patterns[32619] = 25'b01111111_01101001_11101000_0;
      patterns[32620] = 25'b01111111_01101010_11101001_0;
      patterns[32621] = 25'b01111111_01101011_11101010_0;
      patterns[32622] = 25'b01111111_01101100_11101011_0;
      patterns[32623] = 25'b01111111_01101101_11101100_0;
      patterns[32624] = 25'b01111111_01101110_11101101_0;
      patterns[32625] = 25'b01111111_01101111_11101110_0;
      patterns[32626] = 25'b01111111_01110000_11101111_0;
      patterns[32627] = 25'b01111111_01110001_11110000_0;
      patterns[32628] = 25'b01111111_01110010_11110001_0;
      patterns[32629] = 25'b01111111_01110011_11110010_0;
      patterns[32630] = 25'b01111111_01110100_11110011_0;
      patterns[32631] = 25'b01111111_01110101_11110100_0;
      patterns[32632] = 25'b01111111_01110110_11110101_0;
      patterns[32633] = 25'b01111111_01110111_11110110_0;
      patterns[32634] = 25'b01111111_01111000_11110111_0;
      patterns[32635] = 25'b01111111_01111001_11111000_0;
      patterns[32636] = 25'b01111111_01111010_11111001_0;
      patterns[32637] = 25'b01111111_01111011_11111010_0;
      patterns[32638] = 25'b01111111_01111100_11111011_0;
      patterns[32639] = 25'b01111111_01111101_11111100_0;
      patterns[32640] = 25'b01111111_01111110_11111101_0;
      patterns[32641] = 25'b01111111_01111111_11111110_0;
      patterns[32642] = 25'b01111111_10000000_11111111_0;
      patterns[32643] = 25'b01111111_10000001_00000000_1;
      patterns[32644] = 25'b01111111_10000010_00000001_1;
      patterns[32645] = 25'b01111111_10000011_00000010_1;
      patterns[32646] = 25'b01111111_10000100_00000011_1;
      patterns[32647] = 25'b01111111_10000101_00000100_1;
      patterns[32648] = 25'b01111111_10000110_00000101_1;
      patterns[32649] = 25'b01111111_10000111_00000110_1;
      patterns[32650] = 25'b01111111_10001000_00000111_1;
      patterns[32651] = 25'b01111111_10001001_00001000_1;
      patterns[32652] = 25'b01111111_10001010_00001001_1;
      patterns[32653] = 25'b01111111_10001011_00001010_1;
      patterns[32654] = 25'b01111111_10001100_00001011_1;
      patterns[32655] = 25'b01111111_10001101_00001100_1;
      patterns[32656] = 25'b01111111_10001110_00001101_1;
      patterns[32657] = 25'b01111111_10001111_00001110_1;
      patterns[32658] = 25'b01111111_10010000_00001111_1;
      patterns[32659] = 25'b01111111_10010001_00010000_1;
      patterns[32660] = 25'b01111111_10010010_00010001_1;
      patterns[32661] = 25'b01111111_10010011_00010010_1;
      patterns[32662] = 25'b01111111_10010100_00010011_1;
      patterns[32663] = 25'b01111111_10010101_00010100_1;
      patterns[32664] = 25'b01111111_10010110_00010101_1;
      patterns[32665] = 25'b01111111_10010111_00010110_1;
      patterns[32666] = 25'b01111111_10011000_00010111_1;
      patterns[32667] = 25'b01111111_10011001_00011000_1;
      patterns[32668] = 25'b01111111_10011010_00011001_1;
      patterns[32669] = 25'b01111111_10011011_00011010_1;
      patterns[32670] = 25'b01111111_10011100_00011011_1;
      patterns[32671] = 25'b01111111_10011101_00011100_1;
      patterns[32672] = 25'b01111111_10011110_00011101_1;
      patterns[32673] = 25'b01111111_10011111_00011110_1;
      patterns[32674] = 25'b01111111_10100000_00011111_1;
      patterns[32675] = 25'b01111111_10100001_00100000_1;
      patterns[32676] = 25'b01111111_10100010_00100001_1;
      patterns[32677] = 25'b01111111_10100011_00100010_1;
      patterns[32678] = 25'b01111111_10100100_00100011_1;
      patterns[32679] = 25'b01111111_10100101_00100100_1;
      patterns[32680] = 25'b01111111_10100110_00100101_1;
      patterns[32681] = 25'b01111111_10100111_00100110_1;
      patterns[32682] = 25'b01111111_10101000_00100111_1;
      patterns[32683] = 25'b01111111_10101001_00101000_1;
      patterns[32684] = 25'b01111111_10101010_00101001_1;
      patterns[32685] = 25'b01111111_10101011_00101010_1;
      patterns[32686] = 25'b01111111_10101100_00101011_1;
      patterns[32687] = 25'b01111111_10101101_00101100_1;
      patterns[32688] = 25'b01111111_10101110_00101101_1;
      patterns[32689] = 25'b01111111_10101111_00101110_1;
      patterns[32690] = 25'b01111111_10110000_00101111_1;
      patterns[32691] = 25'b01111111_10110001_00110000_1;
      patterns[32692] = 25'b01111111_10110010_00110001_1;
      patterns[32693] = 25'b01111111_10110011_00110010_1;
      patterns[32694] = 25'b01111111_10110100_00110011_1;
      patterns[32695] = 25'b01111111_10110101_00110100_1;
      patterns[32696] = 25'b01111111_10110110_00110101_1;
      patterns[32697] = 25'b01111111_10110111_00110110_1;
      patterns[32698] = 25'b01111111_10111000_00110111_1;
      patterns[32699] = 25'b01111111_10111001_00111000_1;
      patterns[32700] = 25'b01111111_10111010_00111001_1;
      patterns[32701] = 25'b01111111_10111011_00111010_1;
      patterns[32702] = 25'b01111111_10111100_00111011_1;
      patterns[32703] = 25'b01111111_10111101_00111100_1;
      patterns[32704] = 25'b01111111_10111110_00111101_1;
      patterns[32705] = 25'b01111111_10111111_00111110_1;
      patterns[32706] = 25'b01111111_11000000_00111111_1;
      patterns[32707] = 25'b01111111_11000001_01000000_1;
      patterns[32708] = 25'b01111111_11000010_01000001_1;
      patterns[32709] = 25'b01111111_11000011_01000010_1;
      patterns[32710] = 25'b01111111_11000100_01000011_1;
      patterns[32711] = 25'b01111111_11000101_01000100_1;
      patterns[32712] = 25'b01111111_11000110_01000101_1;
      patterns[32713] = 25'b01111111_11000111_01000110_1;
      patterns[32714] = 25'b01111111_11001000_01000111_1;
      patterns[32715] = 25'b01111111_11001001_01001000_1;
      patterns[32716] = 25'b01111111_11001010_01001001_1;
      patterns[32717] = 25'b01111111_11001011_01001010_1;
      patterns[32718] = 25'b01111111_11001100_01001011_1;
      patterns[32719] = 25'b01111111_11001101_01001100_1;
      patterns[32720] = 25'b01111111_11001110_01001101_1;
      patterns[32721] = 25'b01111111_11001111_01001110_1;
      patterns[32722] = 25'b01111111_11010000_01001111_1;
      patterns[32723] = 25'b01111111_11010001_01010000_1;
      patterns[32724] = 25'b01111111_11010010_01010001_1;
      patterns[32725] = 25'b01111111_11010011_01010010_1;
      patterns[32726] = 25'b01111111_11010100_01010011_1;
      patterns[32727] = 25'b01111111_11010101_01010100_1;
      patterns[32728] = 25'b01111111_11010110_01010101_1;
      patterns[32729] = 25'b01111111_11010111_01010110_1;
      patterns[32730] = 25'b01111111_11011000_01010111_1;
      patterns[32731] = 25'b01111111_11011001_01011000_1;
      patterns[32732] = 25'b01111111_11011010_01011001_1;
      patterns[32733] = 25'b01111111_11011011_01011010_1;
      patterns[32734] = 25'b01111111_11011100_01011011_1;
      patterns[32735] = 25'b01111111_11011101_01011100_1;
      patterns[32736] = 25'b01111111_11011110_01011101_1;
      patterns[32737] = 25'b01111111_11011111_01011110_1;
      patterns[32738] = 25'b01111111_11100000_01011111_1;
      patterns[32739] = 25'b01111111_11100001_01100000_1;
      patterns[32740] = 25'b01111111_11100010_01100001_1;
      patterns[32741] = 25'b01111111_11100011_01100010_1;
      patterns[32742] = 25'b01111111_11100100_01100011_1;
      patterns[32743] = 25'b01111111_11100101_01100100_1;
      patterns[32744] = 25'b01111111_11100110_01100101_1;
      patterns[32745] = 25'b01111111_11100111_01100110_1;
      patterns[32746] = 25'b01111111_11101000_01100111_1;
      patterns[32747] = 25'b01111111_11101001_01101000_1;
      patterns[32748] = 25'b01111111_11101010_01101001_1;
      patterns[32749] = 25'b01111111_11101011_01101010_1;
      patterns[32750] = 25'b01111111_11101100_01101011_1;
      patterns[32751] = 25'b01111111_11101101_01101100_1;
      patterns[32752] = 25'b01111111_11101110_01101101_1;
      patterns[32753] = 25'b01111111_11101111_01101110_1;
      patterns[32754] = 25'b01111111_11110000_01101111_1;
      patterns[32755] = 25'b01111111_11110001_01110000_1;
      patterns[32756] = 25'b01111111_11110010_01110001_1;
      patterns[32757] = 25'b01111111_11110011_01110010_1;
      patterns[32758] = 25'b01111111_11110100_01110011_1;
      patterns[32759] = 25'b01111111_11110101_01110100_1;
      patterns[32760] = 25'b01111111_11110110_01110101_1;
      patterns[32761] = 25'b01111111_11110111_01110110_1;
      patterns[32762] = 25'b01111111_11111000_01110111_1;
      patterns[32763] = 25'b01111111_11111001_01111000_1;
      patterns[32764] = 25'b01111111_11111010_01111001_1;
      patterns[32765] = 25'b01111111_11111011_01111010_1;
      patterns[32766] = 25'b01111111_11111100_01111011_1;
      patterns[32767] = 25'b01111111_11111101_01111100_1;
      patterns[32768] = 25'b01111111_11111110_01111101_1;
      patterns[32769] = 25'b01111111_11111111_01111110_1;
      patterns[32770] = 25'b10000000_00000000_10000000_0;
      patterns[32771] = 25'b10000000_00000001_10000001_0;
      patterns[32772] = 25'b10000000_00000010_10000010_0;
      patterns[32773] = 25'b10000000_00000011_10000011_0;
      patterns[32774] = 25'b10000000_00000100_10000100_0;
      patterns[32775] = 25'b10000000_00000101_10000101_0;
      patterns[32776] = 25'b10000000_00000110_10000110_0;
      patterns[32777] = 25'b10000000_00000111_10000111_0;
      patterns[32778] = 25'b10000000_00001000_10001000_0;
      patterns[32779] = 25'b10000000_00001001_10001001_0;
      patterns[32780] = 25'b10000000_00001010_10001010_0;
      patterns[32781] = 25'b10000000_00001011_10001011_0;
      patterns[32782] = 25'b10000000_00001100_10001100_0;
      patterns[32783] = 25'b10000000_00001101_10001101_0;
      patterns[32784] = 25'b10000000_00001110_10001110_0;
      patterns[32785] = 25'b10000000_00001111_10001111_0;
      patterns[32786] = 25'b10000000_00010000_10010000_0;
      patterns[32787] = 25'b10000000_00010001_10010001_0;
      patterns[32788] = 25'b10000000_00010010_10010010_0;
      patterns[32789] = 25'b10000000_00010011_10010011_0;
      patterns[32790] = 25'b10000000_00010100_10010100_0;
      patterns[32791] = 25'b10000000_00010101_10010101_0;
      patterns[32792] = 25'b10000000_00010110_10010110_0;
      patterns[32793] = 25'b10000000_00010111_10010111_0;
      patterns[32794] = 25'b10000000_00011000_10011000_0;
      patterns[32795] = 25'b10000000_00011001_10011001_0;
      patterns[32796] = 25'b10000000_00011010_10011010_0;
      patterns[32797] = 25'b10000000_00011011_10011011_0;
      patterns[32798] = 25'b10000000_00011100_10011100_0;
      patterns[32799] = 25'b10000000_00011101_10011101_0;
      patterns[32800] = 25'b10000000_00011110_10011110_0;
      patterns[32801] = 25'b10000000_00011111_10011111_0;
      patterns[32802] = 25'b10000000_00100000_10100000_0;
      patterns[32803] = 25'b10000000_00100001_10100001_0;
      patterns[32804] = 25'b10000000_00100010_10100010_0;
      patterns[32805] = 25'b10000000_00100011_10100011_0;
      patterns[32806] = 25'b10000000_00100100_10100100_0;
      patterns[32807] = 25'b10000000_00100101_10100101_0;
      patterns[32808] = 25'b10000000_00100110_10100110_0;
      patterns[32809] = 25'b10000000_00100111_10100111_0;
      patterns[32810] = 25'b10000000_00101000_10101000_0;
      patterns[32811] = 25'b10000000_00101001_10101001_0;
      patterns[32812] = 25'b10000000_00101010_10101010_0;
      patterns[32813] = 25'b10000000_00101011_10101011_0;
      patterns[32814] = 25'b10000000_00101100_10101100_0;
      patterns[32815] = 25'b10000000_00101101_10101101_0;
      patterns[32816] = 25'b10000000_00101110_10101110_0;
      patterns[32817] = 25'b10000000_00101111_10101111_0;
      patterns[32818] = 25'b10000000_00110000_10110000_0;
      patterns[32819] = 25'b10000000_00110001_10110001_0;
      patterns[32820] = 25'b10000000_00110010_10110010_0;
      patterns[32821] = 25'b10000000_00110011_10110011_0;
      patterns[32822] = 25'b10000000_00110100_10110100_0;
      patterns[32823] = 25'b10000000_00110101_10110101_0;
      patterns[32824] = 25'b10000000_00110110_10110110_0;
      patterns[32825] = 25'b10000000_00110111_10110111_0;
      patterns[32826] = 25'b10000000_00111000_10111000_0;
      patterns[32827] = 25'b10000000_00111001_10111001_0;
      patterns[32828] = 25'b10000000_00111010_10111010_0;
      patterns[32829] = 25'b10000000_00111011_10111011_0;
      patterns[32830] = 25'b10000000_00111100_10111100_0;
      patterns[32831] = 25'b10000000_00111101_10111101_0;
      patterns[32832] = 25'b10000000_00111110_10111110_0;
      patterns[32833] = 25'b10000000_00111111_10111111_0;
      patterns[32834] = 25'b10000000_01000000_11000000_0;
      patterns[32835] = 25'b10000000_01000001_11000001_0;
      patterns[32836] = 25'b10000000_01000010_11000010_0;
      patterns[32837] = 25'b10000000_01000011_11000011_0;
      patterns[32838] = 25'b10000000_01000100_11000100_0;
      patterns[32839] = 25'b10000000_01000101_11000101_0;
      patterns[32840] = 25'b10000000_01000110_11000110_0;
      patterns[32841] = 25'b10000000_01000111_11000111_0;
      patterns[32842] = 25'b10000000_01001000_11001000_0;
      patterns[32843] = 25'b10000000_01001001_11001001_0;
      patterns[32844] = 25'b10000000_01001010_11001010_0;
      patterns[32845] = 25'b10000000_01001011_11001011_0;
      patterns[32846] = 25'b10000000_01001100_11001100_0;
      patterns[32847] = 25'b10000000_01001101_11001101_0;
      patterns[32848] = 25'b10000000_01001110_11001110_0;
      patterns[32849] = 25'b10000000_01001111_11001111_0;
      patterns[32850] = 25'b10000000_01010000_11010000_0;
      patterns[32851] = 25'b10000000_01010001_11010001_0;
      patterns[32852] = 25'b10000000_01010010_11010010_0;
      patterns[32853] = 25'b10000000_01010011_11010011_0;
      patterns[32854] = 25'b10000000_01010100_11010100_0;
      patterns[32855] = 25'b10000000_01010101_11010101_0;
      patterns[32856] = 25'b10000000_01010110_11010110_0;
      patterns[32857] = 25'b10000000_01010111_11010111_0;
      patterns[32858] = 25'b10000000_01011000_11011000_0;
      patterns[32859] = 25'b10000000_01011001_11011001_0;
      patterns[32860] = 25'b10000000_01011010_11011010_0;
      patterns[32861] = 25'b10000000_01011011_11011011_0;
      patterns[32862] = 25'b10000000_01011100_11011100_0;
      patterns[32863] = 25'b10000000_01011101_11011101_0;
      patterns[32864] = 25'b10000000_01011110_11011110_0;
      patterns[32865] = 25'b10000000_01011111_11011111_0;
      patterns[32866] = 25'b10000000_01100000_11100000_0;
      patterns[32867] = 25'b10000000_01100001_11100001_0;
      patterns[32868] = 25'b10000000_01100010_11100010_0;
      patterns[32869] = 25'b10000000_01100011_11100011_0;
      patterns[32870] = 25'b10000000_01100100_11100100_0;
      patterns[32871] = 25'b10000000_01100101_11100101_0;
      patterns[32872] = 25'b10000000_01100110_11100110_0;
      patterns[32873] = 25'b10000000_01100111_11100111_0;
      patterns[32874] = 25'b10000000_01101000_11101000_0;
      patterns[32875] = 25'b10000000_01101001_11101001_0;
      patterns[32876] = 25'b10000000_01101010_11101010_0;
      patterns[32877] = 25'b10000000_01101011_11101011_0;
      patterns[32878] = 25'b10000000_01101100_11101100_0;
      patterns[32879] = 25'b10000000_01101101_11101101_0;
      patterns[32880] = 25'b10000000_01101110_11101110_0;
      patterns[32881] = 25'b10000000_01101111_11101111_0;
      patterns[32882] = 25'b10000000_01110000_11110000_0;
      patterns[32883] = 25'b10000000_01110001_11110001_0;
      patterns[32884] = 25'b10000000_01110010_11110010_0;
      patterns[32885] = 25'b10000000_01110011_11110011_0;
      patterns[32886] = 25'b10000000_01110100_11110100_0;
      patterns[32887] = 25'b10000000_01110101_11110101_0;
      patterns[32888] = 25'b10000000_01110110_11110110_0;
      patterns[32889] = 25'b10000000_01110111_11110111_0;
      patterns[32890] = 25'b10000000_01111000_11111000_0;
      patterns[32891] = 25'b10000000_01111001_11111001_0;
      patterns[32892] = 25'b10000000_01111010_11111010_0;
      patterns[32893] = 25'b10000000_01111011_11111011_0;
      patterns[32894] = 25'b10000000_01111100_11111100_0;
      patterns[32895] = 25'b10000000_01111101_11111101_0;
      patterns[32896] = 25'b10000000_01111110_11111110_0;
      patterns[32897] = 25'b10000000_01111111_11111111_0;
      patterns[32898] = 25'b10000000_10000000_00000000_1;
      patterns[32899] = 25'b10000000_10000001_00000001_1;
      patterns[32900] = 25'b10000000_10000010_00000010_1;
      patterns[32901] = 25'b10000000_10000011_00000011_1;
      patterns[32902] = 25'b10000000_10000100_00000100_1;
      patterns[32903] = 25'b10000000_10000101_00000101_1;
      patterns[32904] = 25'b10000000_10000110_00000110_1;
      patterns[32905] = 25'b10000000_10000111_00000111_1;
      patterns[32906] = 25'b10000000_10001000_00001000_1;
      patterns[32907] = 25'b10000000_10001001_00001001_1;
      patterns[32908] = 25'b10000000_10001010_00001010_1;
      patterns[32909] = 25'b10000000_10001011_00001011_1;
      patterns[32910] = 25'b10000000_10001100_00001100_1;
      patterns[32911] = 25'b10000000_10001101_00001101_1;
      patterns[32912] = 25'b10000000_10001110_00001110_1;
      patterns[32913] = 25'b10000000_10001111_00001111_1;
      patterns[32914] = 25'b10000000_10010000_00010000_1;
      patterns[32915] = 25'b10000000_10010001_00010001_1;
      patterns[32916] = 25'b10000000_10010010_00010010_1;
      patterns[32917] = 25'b10000000_10010011_00010011_1;
      patterns[32918] = 25'b10000000_10010100_00010100_1;
      patterns[32919] = 25'b10000000_10010101_00010101_1;
      patterns[32920] = 25'b10000000_10010110_00010110_1;
      patterns[32921] = 25'b10000000_10010111_00010111_1;
      patterns[32922] = 25'b10000000_10011000_00011000_1;
      patterns[32923] = 25'b10000000_10011001_00011001_1;
      patterns[32924] = 25'b10000000_10011010_00011010_1;
      patterns[32925] = 25'b10000000_10011011_00011011_1;
      patterns[32926] = 25'b10000000_10011100_00011100_1;
      patterns[32927] = 25'b10000000_10011101_00011101_1;
      patterns[32928] = 25'b10000000_10011110_00011110_1;
      patterns[32929] = 25'b10000000_10011111_00011111_1;
      patterns[32930] = 25'b10000000_10100000_00100000_1;
      patterns[32931] = 25'b10000000_10100001_00100001_1;
      patterns[32932] = 25'b10000000_10100010_00100010_1;
      patterns[32933] = 25'b10000000_10100011_00100011_1;
      patterns[32934] = 25'b10000000_10100100_00100100_1;
      patterns[32935] = 25'b10000000_10100101_00100101_1;
      patterns[32936] = 25'b10000000_10100110_00100110_1;
      patterns[32937] = 25'b10000000_10100111_00100111_1;
      patterns[32938] = 25'b10000000_10101000_00101000_1;
      patterns[32939] = 25'b10000000_10101001_00101001_1;
      patterns[32940] = 25'b10000000_10101010_00101010_1;
      patterns[32941] = 25'b10000000_10101011_00101011_1;
      patterns[32942] = 25'b10000000_10101100_00101100_1;
      patterns[32943] = 25'b10000000_10101101_00101101_1;
      patterns[32944] = 25'b10000000_10101110_00101110_1;
      patterns[32945] = 25'b10000000_10101111_00101111_1;
      patterns[32946] = 25'b10000000_10110000_00110000_1;
      patterns[32947] = 25'b10000000_10110001_00110001_1;
      patterns[32948] = 25'b10000000_10110010_00110010_1;
      patterns[32949] = 25'b10000000_10110011_00110011_1;
      patterns[32950] = 25'b10000000_10110100_00110100_1;
      patterns[32951] = 25'b10000000_10110101_00110101_1;
      patterns[32952] = 25'b10000000_10110110_00110110_1;
      patterns[32953] = 25'b10000000_10110111_00110111_1;
      patterns[32954] = 25'b10000000_10111000_00111000_1;
      patterns[32955] = 25'b10000000_10111001_00111001_1;
      patterns[32956] = 25'b10000000_10111010_00111010_1;
      patterns[32957] = 25'b10000000_10111011_00111011_1;
      patterns[32958] = 25'b10000000_10111100_00111100_1;
      patterns[32959] = 25'b10000000_10111101_00111101_1;
      patterns[32960] = 25'b10000000_10111110_00111110_1;
      patterns[32961] = 25'b10000000_10111111_00111111_1;
      patterns[32962] = 25'b10000000_11000000_01000000_1;
      patterns[32963] = 25'b10000000_11000001_01000001_1;
      patterns[32964] = 25'b10000000_11000010_01000010_1;
      patterns[32965] = 25'b10000000_11000011_01000011_1;
      patterns[32966] = 25'b10000000_11000100_01000100_1;
      patterns[32967] = 25'b10000000_11000101_01000101_1;
      patterns[32968] = 25'b10000000_11000110_01000110_1;
      patterns[32969] = 25'b10000000_11000111_01000111_1;
      patterns[32970] = 25'b10000000_11001000_01001000_1;
      patterns[32971] = 25'b10000000_11001001_01001001_1;
      patterns[32972] = 25'b10000000_11001010_01001010_1;
      patterns[32973] = 25'b10000000_11001011_01001011_1;
      patterns[32974] = 25'b10000000_11001100_01001100_1;
      patterns[32975] = 25'b10000000_11001101_01001101_1;
      patterns[32976] = 25'b10000000_11001110_01001110_1;
      patterns[32977] = 25'b10000000_11001111_01001111_1;
      patterns[32978] = 25'b10000000_11010000_01010000_1;
      patterns[32979] = 25'b10000000_11010001_01010001_1;
      patterns[32980] = 25'b10000000_11010010_01010010_1;
      patterns[32981] = 25'b10000000_11010011_01010011_1;
      patterns[32982] = 25'b10000000_11010100_01010100_1;
      patterns[32983] = 25'b10000000_11010101_01010101_1;
      patterns[32984] = 25'b10000000_11010110_01010110_1;
      patterns[32985] = 25'b10000000_11010111_01010111_1;
      patterns[32986] = 25'b10000000_11011000_01011000_1;
      patterns[32987] = 25'b10000000_11011001_01011001_1;
      patterns[32988] = 25'b10000000_11011010_01011010_1;
      patterns[32989] = 25'b10000000_11011011_01011011_1;
      patterns[32990] = 25'b10000000_11011100_01011100_1;
      patterns[32991] = 25'b10000000_11011101_01011101_1;
      patterns[32992] = 25'b10000000_11011110_01011110_1;
      patterns[32993] = 25'b10000000_11011111_01011111_1;
      patterns[32994] = 25'b10000000_11100000_01100000_1;
      patterns[32995] = 25'b10000000_11100001_01100001_1;
      patterns[32996] = 25'b10000000_11100010_01100010_1;
      patterns[32997] = 25'b10000000_11100011_01100011_1;
      patterns[32998] = 25'b10000000_11100100_01100100_1;
      patterns[32999] = 25'b10000000_11100101_01100101_1;
      patterns[33000] = 25'b10000000_11100110_01100110_1;
      patterns[33001] = 25'b10000000_11100111_01100111_1;
      patterns[33002] = 25'b10000000_11101000_01101000_1;
      patterns[33003] = 25'b10000000_11101001_01101001_1;
      patterns[33004] = 25'b10000000_11101010_01101010_1;
      patterns[33005] = 25'b10000000_11101011_01101011_1;
      patterns[33006] = 25'b10000000_11101100_01101100_1;
      patterns[33007] = 25'b10000000_11101101_01101101_1;
      patterns[33008] = 25'b10000000_11101110_01101110_1;
      patterns[33009] = 25'b10000000_11101111_01101111_1;
      patterns[33010] = 25'b10000000_11110000_01110000_1;
      patterns[33011] = 25'b10000000_11110001_01110001_1;
      patterns[33012] = 25'b10000000_11110010_01110010_1;
      patterns[33013] = 25'b10000000_11110011_01110011_1;
      patterns[33014] = 25'b10000000_11110100_01110100_1;
      patterns[33015] = 25'b10000000_11110101_01110101_1;
      patterns[33016] = 25'b10000000_11110110_01110110_1;
      patterns[33017] = 25'b10000000_11110111_01110111_1;
      patterns[33018] = 25'b10000000_11111000_01111000_1;
      patterns[33019] = 25'b10000000_11111001_01111001_1;
      patterns[33020] = 25'b10000000_11111010_01111010_1;
      patterns[33021] = 25'b10000000_11111011_01111011_1;
      patterns[33022] = 25'b10000000_11111100_01111100_1;
      patterns[33023] = 25'b10000000_11111101_01111101_1;
      patterns[33024] = 25'b10000000_11111110_01111110_1;
      patterns[33025] = 25'b10000000_11111111_01111111_1;
      patterns[33026] = 25'b10000001_00000000_10000001_0;
      patterns[33027] = 25'b10000001_00000001_10000010_0;
      patterns[33028] = 25'b10000001_00000010_10000011_0;
      patterns[33029] = 25'b10000001_00000011_10000100_0;
      patterns[33030] = 25'b10000001_00000100_10000101_0;
      patterns[33031] = 25'b10000001_00000101_10000110_0;
      patterns[33032] = 25'b10000001_00000110_10000111_0;
      patterns[33033] = 25'b10000001_00000111_10001000_0;
      patterns[33034] = 25'b10000001_00001000_10001001_0;
      patterns[33035] = 25'b10000001_00001001_10001010_0;
      patterns[33036] = 25'b10000001_00001010_10001011_0;
      patterns[33037] = 25'b10000001_00001011_10001100_0;
      patterns[33038] = 25'b10000001_00001100_10001101_0;
      patterns[33039] = 25'b10000001_00001101_10001110_0;
      patterns[33040] = 25'b10000001_00001110_10001111_0;
      patterns[33041] = 25'b10000001_00001111_10010000_0;
      patterns[33042] = 25'b10000001_00010000_10010001_0;
      patterns[33043] = 25'b10000001_00010001_10010010_0;
      patterns[33044] = 25'b10000001_00010010_10010011_0;
      patterns[33045] = 25'b10000001_00010011_10010100_0;
      patterns[33046] = 25'b10000001_00010100_10010101_0;
      patterns[33047] = 25'b10000001_00010101_10010110_0;
      patterns[33048] = 25'b10000001_00010110_10010111_0;
      patterns[33049] = 25'b10000001_00010111_10011000_0;
      patterns[33050] = 25'b10000001_00011000_10011001_0;
      patterns[33051] = 25'b10000001_00011001_10011010_0;
      patterns[33052] = 25'b10000001_00011010_10011011_0;
      patterns[33053] = 25'b10000001_00011011_10011100_0;
      patterns[33054] = 25'b10000001_00011100_10011101_0;
      patterns[33055] = 25'b10000001_00011101_10011110_0;
      patterns[33056] = 25'b10000001_00011110_10011111_0;
      patterns[33057] = 25'b10000001_00011111_10100000_0;
      patterns[33058] = 25'b10000001_00100000_10100001_0;
      patterns[33059] = 25'b10000001_00100001_10100010_0;
      patterns[33060] = 25'b10000001_00100010_10100011_0;
      patterns[33061] = 25'b10000001_00100011_10100100_0;
      patterns[33062] = 25'b10000001_00100100_10100101_0;
      patterns[33063] = 25'b10000001_00100101_10100110_0;
      patterns[33064] = 25'b10000001_00100110_10100111_0;
      patterns[33065] = 25'b10000001_00100111_10101000_0;
      patterns[33066] = 25'b10000001_00101000_10101001_0;
      patterns[33067] = 25'b10000001_00101001_10101010_0;
      patterns[33068] = 25'b10000001_00101010_10101011_0;
      patterns[33069] = 25'b10000001_00101011_10101100_0;
      patterns[33070] = 25'b10000001_00101100_10101101_0;
      patterns[33071] = 25'b10000001_00101101_10101110_0;
      patterns[33072] = 25'b10000001_00101110_10101111_0;
      patterns[33073] = 25'b10000001_00101111_10110000_0;
      patterns[33074] = 25'b10000001_00110000_10110001_0;
      patterns[33075] = 25'b10000001_00110001_10110010_0;
      patterns[33076] = 25'b10000001_00110010_10110011_0;
      patterns[33077] = 25'b10000001_00110011_10110100_0;
      patterns[33078] = 25'b10000001_00110100_10110101_0;
      patterns[33079] = 25'b10000001_00110101_10110110_0;
      patterns[33080] = 25'b10000001_00110110_10110111_0;
      patterns[33081] = 25'b10000001_00110111_10111000_0;
      patterns[33082] = 25'b10000001_00111000_10111001_0;
      patterns[33083] = 25'b10000001_00111001_10111010_0;
      patterns[33084] = 25'b10000001_00111010_10111011_0;
      patterns[33085] = 25'b10000001_00111011_10111100_0;
      patterns[33086] = 25'b10000001_00111100_10111101_0;
      patterns[33087] = 25'b10000001_00111101_10111110_0;
      patterns[33088] = 25'b10000001_00111110_10111111_0;
      patterns[33089] = 25'b10000001_00111111_11000000_0;
      patterns[33090] = 25'b10000001_01000000_11000001_0;
      patterns[33091] = 25'b10000001_01000001_11000010_0;
      patterns[33092] = 25'b10000001_01000010_11000011_0;
      patterns[33093] = 25'b10000001_01000011_11000100_0;
      patterns[33094] = 25'b10000001_01000100_11000101_0;
      patterns[33095] = 25'b10000001_01000101_11000110_0;
      patterns[33096] = 25'b10000001_01000110_11000111_0;
      patterns[33097] = 25'b10000001_01000111_11001000_0;
      patterns[33098] = 25'b10000001_01001000_11001001_0;
      patterns[33099] = 25'b10000001_01001001_11001010_0;
      patterns[33100] = 25'b10000001_01001010_11001011_0;
      patterns[33101] = 25'b10000001_01001011_11001100_0;
      patterns[33102] = 25'b10000001_01001100_11001101_0;
      patterns[33103] = 25'b10000001_01001101_11001110_0;
      patterns[33104] = 25'b10000001_01001110_11001111_0;
      patterns[33105] = 25'b10000001_01001111_11010000_0;
      patterns[33106] = 25'b10000001_01010000_11010001_0;
      patterns[33107] = 25'b10000001_01010001_11010010_0;
      patterns[33108] = 25'b10000001_01010010_11010011_0;
      patterns[33109] = 25'b10000001_01010011_11010100_0;
      patterns[33110] = 25'b10000001_01010100_11010101_0;
      patterns[33111] = 25'b10000001_01010101_11010110_0;
      patterns[33112] = 25'b10000001_01010110_11010111_0;
      patterns[33113] = 25'b10000001_01010111_11011000_0;
      patterns[33114] = 25'b10000001_01011000_11011001_0;
      patterns[33115] = 25'b10000001_01011001_11011010_0;
      patterns[33116] = 25'b10000001_01011010_11011011_0;
      patterns[33117] = 25'b10000001_01011011_11011100_0;
      patterns[33118] = 25'b10000001_01011100_11011101_0;
      patterns[33119] = 25'b10000001_01011101_11011110_0;
      patterns[33120] = 25'b10000001_01011110_11011111_0;
      patterns[33121] = 25'b10000001_01011111_11100000_0;
      patterns[33122] = 25'b10000001_01100000_11100001_0;
      patterns[33123] = 25'b10000001_01100001_11100010_0;
      patterns[33124] = 25'b10000001_01100010_11100011_0;
      patterns[33125] = 25'b10000001_01100011_11100100_0;
      patterns[33126] = 25'b10000001_01100100_11100101_0;
      patterns[33127] = 25'b10000001_01100101_11100110_0;
      patterns[33128] = 25'b10000001_01100110_11100111_0;
      patterns[33129] = 25'b10000001_01100111_11101000_0;
      patterns[33130] = 25'b10000001_01101000_11101001_0;
      patterns[33131] = 25'b10000001_01101001_11101010_0;
      patterns[33132] = 25'b10000001_01101010_11101011_0;
      patterns[33133] = 25'b10000001_01101011_11101100_0;
      patterns[33134] = 25'b10000001_01101100_11101101_0;
      patterns[33135] = 25'b10000001_01101101_11101110_0;
      patterns[33136] = 25'b10000001_01101110_11101111_0;
      patterns[33137] = 25'b10000001_01101111_11110000_0;
      patterns[33138] = 25'b10000001_01110000_11110001_0;
      patterns[33139] = 25'b10000001_01110001_11110010_0;
      patterns[33140] = 25'b10000001_01110010_11110011_0;
      patterns[33141] = 25'b10000001_01110011_11110100_0;
      patterns[33142] = 25'b10000001_01110100_11110101_0;
      patterns[33143] = 25'b10000001_01110101_11110110_0;
      patterns[33144] = 25'b10000001_01110110_11110111_0;
      patterns[33145] = 25'b10000001_01110111_11111000_0;
      patterns[33146] = 25'b10000001_01111000_11111001_0;
      patterns[33147] = 25'b10000001_01111001_11111010_0;
      patterns[33148] = 25'b10000001_01111010_11111011_0;
      patterns[33149] = 25'b10000001_01111011_11111100_0;
      patterns[33150] = 25'b10000001_01111100_11111101_0;
      patterns[33151] = 25'b10000001_01111101_11111110_0;
      patterns[33152] = 25'b10000001_01111110_11111111_0;
      patterns[33153] = 25'b10000001_01111111_00000000_1;
      patterns[33154] = 25'b10000001_10000000_00000001_1;
      patterns[33155] = 25'b10000001_10000001_00000010_1;
      patterns[33156] = 25'b10000001_10000010_00000011_1;
      patterns[33157] = 25'b10000001_10000011_00000100_1;
      patterns[33158] = 25'b10000001_10000100_00000101_1;
      patterns[33159] = 25'b10000001_10000101_00000110_1;
      patterns[33160] = 25'b10000001_10000110_00000111_1;
      patterns[33161] = 25'b10000001_10000111_00001000_1;
      patterns[33162] = 25'b10000001_10001000_00001001_1;
      patterns[33163] = 25'b10000001_10001001_00001010_1;
      patterns[33164] = 25'b10000001_10001010_00001011_1;
      patterns[33165] = 25'b10000001_10001011_00001100_1;
      patterns[33166] = 25'b10000001_10001100_00001101_1;
      patterns[33167] = 25'b10000001_10001101_00001110_1;
      patterns[33168] = 25'b10000001_10001110_00001111_1;
      patterns[33169] = 25'b10000001_10001111_00010000_1;
      patterns[33170] = 25'b10000001_10010000_00010001_1;
      patterns[33171] = 25'b10000001_10010001_00010010_1;
      patterns[33172] = 25'b10000001_10010010_00010011_1;
      patterns[33173] = 25'b10000001_10010011_00010100_1;
      patterns[33174] = 25'b10000001_10010100_00010101_1;
      patterns[33175] = 25'b10000001_10010101_00010110_1;
      patterns[33176] = 25'b10000001_10010110_00010111_1;
      patterns[33177] = 25'b10000001_10010111_00011000_1;
      patterns[33178] = 25'b10000001_10011000_00011001_1;
      patterns[33179] = 25'b10000001_10011001_00011010_1;
      patterns[33180] = 25'b10000001_10011010_00011011_1;
      patterns[33181] = 25'b10000001_10011011_00011100_1;
      patterns[33182] = 25'b10000001_10011100_00011101_1;
      patterns[33183] = 25'b10000001_10011101_00011110_1;
      patterns[33184] = 25'b10000001_10011110_00011111_1;
      patterns[33185] = 25'b10000001_10011111_00100000_1;
      patterns[33186] = 25'b10000001_10100000_00100001_1;
      patterns[33187] = 25'b10000001_10100001_00100010_1;
      patterns[33188] = 25'b10000001_10100010_00100011_1;
      patterns[33189] = 25'b10000001_10100011_00100100_1;
      patterns[33190] = 25'b10000001_10100100_00100101_1;
      patterns[33191] = 25'b10000001_10100101_00100110_1;
      patterns[33192] = 25'b10000001_10100110_00100111_1;
      patterns[33193] = 25'b10000001_10100111_00101000_1;
      patterns[33194] = 25'b10000001_10101000_00101001_1;
      patterns[33195] = 25'b10000001_10101001_00101010_1;
      patterns[33196] = 25'b10000001_10101010_00101011_1;
      patterns[33197] = 25'b10000001_10101011_00101100_1;
      patterns[33198] = 25'b10000001_10101100_00101101_1;
      patterns[33199] = 25'b10000001_10101101_00101110_1;
      patterns[33200] = 25'b10000001_10101110_00101111_1;
      patterns[33201] = 25'b10000001_10101111_00110000_1;
      patterns[33202] = 25'b10000001_10110000_00110001_1;
      patterns[33203] = 25'b10000001_10110001_00110010_1;
      patterns[33204] = 25'b10000001_10110010_00110011_1;
      patterns[33205] = 25'b10000001_10110011_00110100_1;
      patterns[33206] = 25'b10000001_10110100_00110101_1;
      patterns[33207] = 25'b10000001_10110101_00110110_1;
      patterns[33208] = 25'b10000001_10110110_00110111_1;
      patterns[33209] = 25'b10000001_10110111_00111000_1;
      patterns[33210] = 25'b10000001_10111000_00111001_1;
      patterns[33211] = 25'b10000001_10111001_00111010_1;
      patterns[33212] = 25'b10000001_10111010_00111011_1;
      patterns[33213] = 25'b10000001_10111011_00111100_1;
      patterns[33214] = 25'b10000001_10111100_00111101_1;
      patterns[33215] = 25'b10000001_10111101_00111110_1;
      patterns[33216] = 25'b10000001_10111110_00111111_1;
      patterns[33217] = 25'b10000001_10111111_01000000_1;
      patterns[33218] = 25'b10000001_11000000_01000001_1;
      patterns[33219] = 25'b10000001_11000001_01000010_1;
      patterns[33220] = 25'b10000001_11000010_01000011_1;
      patterns[33221] = 25'b10000001_11000011_01000100_1;
      patterns[33222] = 25'b10000001_11000100_01000101_1;
      patterns[33223] = 25'b10000001_11000101_01000110_1;
      patterns[33224] = 25'b10000001_11000110_01000111_1;
      patterns[33225] = 25'b10000001_11000111_01001000_1;
      patterns[33226] = 25'b10000001_11001000_01001001_1;
      patterns[33227] = 25'b10000001_11001001_01001010_1;
      patterns[33228] = 25'b10000001_11001010_01001011_1;
      patterns[33229] = 25'b10000001_11001011_01001100_1;
      patterns[33230] = 25'b10000001_11001100_01001101_1;
      patterns[33231] = 25'b10000001_11001101_01001110_1;
      patterns[33232] = 25'b10000001_11001110_01001111_1;
      patterns[33233] = 25'b10000001_11001111_01010000_1;
      patterns[33234] = 25'b10000001_11010000_01010001_1;
      patterns[33235] = 25'b10000001_11010001_01010010_1;
      patterns[33236] = 25'b10000001_11010010_01010011_1;
      patterns[33237] = 25'b10000001_11010011_01010100_1;
      patterns[33238] = 25'b10000001_11010100_01010101_1;
      patterns[33239] = 25'b10000001_11010101_01010110_1;
      patterns[33240] = 25'b10000001_11010110_01010111_1;
      patterns[33241] = 25'b10000001_11010111_01011000_1;
      patterns[33242] = 25'b10000001_11011000_01011001_1;
      patterns[33243] = 25'b10000001_11011001_01011010_1;
      patterns[33244] = 25'b10000001_11011010_01011011_1;
      patterns[33245] = 25'b10000001_11011011_01011100_1;
      patterns[33246] = 25'b10000001_11011100_01011101_1;
      patterns[33247] = 25'b10000001_11011101_01011110_1;
      patterns[33248] = 25'b10000001_11011110_01011111_1;
      patterns[33249] = 25'b10000001_11011111_01100000_1;
      patterns[33250] = 25'b10000001_11100000_01100001_1;
      patterns[33251] = 25'b10000001_11100001_01100010_1;
      patterns[33252] = 25'b10000001_11100010_01100011_1;
      patterns[33253] = 25'b10000001_11100011_01100100_1;
      patterns[33254] = 25'b10000001_11100100_01100101_1;
      patterns[33255] = 25'b10000001_11100101_01100110_1;
      patterns[33256] = 25'b10000001_11100110_01100111_1;
      patterns[33257] = 25'b10000001_11100111_01101000_1;
      patterns[33258] = 25'b10000001_11101000_01101001_1;
      patterns[33259] = 25'b10000001_11101001_01101010_1;
      patterns[33260] = 25'b10000001_11101010_01101011_1;
      patterns[33261] = 25'b10000001_11101011_01101100_1;
      patterns[33262] = 25'b10000001_11101100_01101101_1;
      patterns[33263] = 25'b10000001_11101101_01101110_1;
      patterns[33264] = 25'b10000001_11101110_01101111_1;
      patterns[33265] = 25'b10000001_11101111_01110000_1;
      patterns[33266] = 25'b10000001_11110000_01110001_1;
      patterns[33267] = 25'b10000001_11110001_01110010_1;
      patterns[33268] = 25'b10000001_11110010_01110011_1;
      patterns[33269] = 25'b10000001_11110011_01110100_1;
      patterns[33270] = 25'b10000001_11110100_01110101_1;
      patterns[33271] = 25'b10000001_11110101_01110110_1;
      patterns[33272] = 25'b10000001_11110110_01110111_1;
      patterns[33273] = 25'b10000001_11110111_01111000_1;
      patterns[33274] = 25'b10000001_11111000_01111001_1;
      patterns[33275] = 25'b10000001_11111001_01111010_1;
      patterns[33276] = 25'b10000001_11111010_01111011_1;
      patterns[33277] = 25'b10000001_11111011_01111100_1;
      patterns[33278] = 25'b10000001_11111100_01111101_1;
      patterns[33279] = 25'b10000001_11111101_01111110_1;
      patterns[33280] = 25'b10000001_11111110_01111111_1;
      patterns[33281] = 25'b10000001_11111111_10000000_1;
      patterns[33282] = 25'b10000010_00000000_10000010_0;
      patterns[33283] = 25'b10000010_00000001_10000011_0;
      patterns[33284] = 25'b10000010_00000010_10000100_0;
      patterns[33285] = 25'b10000010_00000011_10000101_0;
      patterns[33286] = 25'b10000010_00000100_10000110_0;
      patterns[33287] = 25'b10000010_00000101_10000111_0;
      patterns[33288] = 25'b10000010_00000110_10001000_0;
      patterns[33289] = 25'b10000010_00000111_10001001_0;
      patterns[33290] = 25'b10000010_00001000_10001010_0;
      patterns[33291] = 25'b10000010_00001001_10001011_0;
      patterns[33292] = 25'b10000010_00001010_10001100_0;
      patterns[33293] = 25'b10000010_00001011_10001101_0;
      patterns[33294] = 25'b10000010_00001100_10001110_0;
      patterns[33295] = 25'b10000010_00001101_10001111_0;
      patterns[33296] = 25'b10000010_00001110_10010000_0;
      patterns[33297] = 25'b10000010_00001111_10010001_0;
      patterns[33298] = 25'b10000010_00010000_10010010_0;
      patterns[33299] = 25'b10000010_00010001_10010011_0;
      patterns[33300] = 25'b10000010_00010010_10010100_0;
      patterns[33301] = 25'b10000010_00010011_10010101_0;
      patterns[33302] = 25'b10000010_00010100_10010110_0;
      patterns[33303] = 25'b10000010_00010101_10010111_0;
      patterns[33304] = 25'b10000010_00010110_10011000_0;
      patterns[33305] = 25'b10000010_00010111_10011001_0;
      patterns[33306] = 25'b10000010_00011000_10011010_0;
      patterns[33307] = 25'b10000010_00011001_10011011_0;
      patterns[33308] = 25'b10000010_00011010_10011100_0;
      patterns[33309] = 25'b10000010_00011011_10011101_0;
      patterns[33310] = 25'b10000010_00011100_10011110_0;
      patterns[33311] = 25'b10000010_00011101_10011111_0;
      patterns[33312] = 25'b10000010_00011110_10100000_0;
      patterns[33313] = 25'b10000010_00011111_10100001_0;
      patterns[33314] = 25'b10000010_00100000_10100010_0;
      patterns[33315] = 25'b10000010_00100001_10100011_0;
      patterns[33316] = 25'b10000010_00100010_10100100_0;
      patterns[33317] = 25'b10000010_00100011_10100101_0;
      patterns[33318] = 25'b10000010_00100100_10100110_0;
      patterns[33319] = 25'b10000010_00100101_10100111_0;
      patterns[33320] = 25'b10000010_00100110_10101000_0;
      patterns[33321] = 25'b10000010_00100111_10101001_0;
      patterns[33322] = 25'b10000010_00101000_10101010_0;
      patterns[33323] = 25'b10000010_00101001_10101011_0;
      patterns[33324] = 25'b10000010_00101010_10101100_0;
      patterns[33325] = 25'b10000010_00101011_10101101_0;
      patterns[33326] = 25'b10000010_00101100_10101110_0;
      patterns[33327] = 25'b10000010_00101101_10101111_0;
      patterns[33328] = 25'b10000010_00101110_10110000_0;
      patterns[33329] = 25'b10000010_00101111_10110001_0;
      patterns[33330] = 25'b10000010_00110000_10110010_0;
      patterns[33331] = 25'b10000010_00110001_10110011_0;
      patterns[33332] = 25'b10000010_00110010_10110100_0;
      patterns[33333] = 25'b10000010_00110011_10110101_0;
      patterns[33334] = 25'b10000010_00110100_10110110_0;
      patterns[33335] = 25'b10000010_00110101_10110111_0;
      patterns[33336] = 25'b10000010_00110110_10111000_0;
      patterns[33337] = 25'b10000010_00110111_10111001_0;
      patterns[33338] = 25'b10000010_00111000_10111010_0;
      patterns[33339] = 25'b10000010_00111001_10111011_0;
      patterns[33340] = 25'b10000010_00111010_10111100_0;
      patterns[33341] = 25'b10000010_00111011_10111101_0;
      patterns[33342] = 25'b10000010_00111100_10111110_0;
      patterns[33343] = 25'b10000010_00111101_10111111_0;
      patterns[33344] = 25'b10000010_00111110_11000000_0;
      patterns[33345] = 25'b10000010_00111111_11000001_0;
      patterns[33346] = 25'b10000010_01000000_11000010_0;
      patterns[33347] = 25'b10000010_01000001_11000011_0;
      patterns[33348] = 25'b10000010_01000010_11000100_0;
      patterns[33349] = 25'b10000010_01000011_11000101_0;
      patterns[33350] = 25'b10000010_01000100_11000110_0;
      patterns[33351] = 25'b10000010_01000101_11000111_0;
      patterns[33352] = 25'b10000010_01000110_11001000_0;
      patterns[33353] = 25'b10000010_01000111_11001001_0;
      patterns[33354] = 25'b10000010_01001000_11001010_0;
      patterns[33355] = 25'b10000010_01001001_11001011_0;
      patterns[33356] = 25'b10000010_01001010_11001100_0;
      patterns[33357] = 25'b10000010_01001011_11001101_0;
      patterns[33358] = 25'b10000010_01001100_11001110_0;
      patterns[33359] = 25'b10000010_01001101_11001111_0;
      patterns[33360] = 25'b10000010_01001110_11010000_0;
      patterns[33361] = 25'b10000010_01001111_11010001_0;
      patterns[33362] = 25'b10000010_01010000_11010010_0;
      patterns[33363] = 25'b10000010_01010001_11010011_0;
      patterns[33364] = 25'b10000010_01010010_11010100_0;
      patterns[33365] = 25'b10000010_01010011_11010101_0;
      patterns[33366] = 25'b10000010_01010100_11010110_0;
      patterns[33367] = 25'b10000010_01010101_11010111_0;
      patterns[33368] = 25'b10000010_01010110_11011000_0;
      patterns[33369] = 25'b10000010_01010111_11011001_0;
      patterns[33370] = 25'b10000010_01011000_11011010_0;
      patterns[33371] = 25'b10000010_01011001_11011011_0;
      patterns[33372] = 25'b10000010_01011010_11011100_0;
      patterns[33373] = 25'b10000010_01011011_11011101_0;
      patterns[33374] = 25'b10000010_01011100_11011110_0;
      patterns[33375] = 25'b10000010_01011101_11011111_0;
      patterns[33376] = 25'b10000010_01011110_11100000_0;
      patterns[33377] = 25'b10000010_01011111_11100001_0;
      patterns[33378] = 25'b10000010_01100000_11100010_0;
      patterns[33379] = 25'b10000010_01100001_11100011_0;
      patterns[33380] = 25'b10000010_01100010_11100100_0;
      patterns[33381] = 25'b10000010_01100011_11100101_0;
      patterns[33382] = 25'b10000010_01100100_11100110_0;
      patterns[33383] = 25'b10000010_01100101_11100111_0;
      patterns[33384] = 25'b10000010_01100110_11101000_0;
      patterns[33385] = 25'b10000010_01100111_11101001_0;
      patterns[33386] = 25'b10000010_01101000_11101010_0;
      patterns[33387] = 25'b10000010_01101001_11101011_0;
      patterns[33388] = 25'b10000010_01101010_11101100_0;
      patterns[33389] = 25'b10000010_01101011_11101101_0;
      patterns[33390] = 25'b10000010_01101100_11101110_0;
      patterns[33391] = 25'b10000010_01101101_11101111_0;
      patterns[33392] = 25'b10000010_01101110_11110000_0;
      patterns[33393] = 25'b10000010_01101111_11110001_0;
      patterns[33394] = 25'b10000010_01110000_11110010_0;
      patterns[33395] = 25'b10000010_01110001_11110011_0;
      patterns[33396] = 25'b10000010_01110010_11110100_0;
      patterns[33397] = 25'b10000010_01110011_11110101_0;
      patterns[33398] = 25'b10000010_01110100_11110110_0;
      patterns[33399] = 25'b10000010_01110101_11110111_0;
      patterns[33400] = 25'b10000010_01110110_11111000_0;
      patterns[33401] = 25'b10000010_01110111_11111001_0;
      patterns[33402] = 25'b10000010_01111000_11111010_0;
      patterns[33403] = 25'b10000010_01111001_11111011_0;
      patterns[33404] = 25'b10000010_01111010_11111100_0;
      patterns[33405] = 25'b10000010_01111011_11111101_0;
      patterns[33406] = 25'b10000010_01111100_11111110_0;
      patterns[33407] = 25'b10000010_01111101_11111111_0;
      patterns[33408] = 25'b10000010_01111110_00000000_1;
      patterns[33409] = 25'b10000010_01111111_00000001_1;
      patterns[33410] = 25'b10000010_10000000_00000010_1;
      patterns[33411] = 25'b10000010_10000001_00000011_1;
      patterns[33412] = 25'b10000010_10000010_00000100_1;
      patterns[33413] = 25'b10000010_10000011_00000101_1;
      patterns[33414] = 25'b10000010_10000100_00000110_1;
      patterns[33415] = 25'b10000010_10000101_00000111_1;
      patterns[33416] = 25'b10000010_10000110_00001000_1;
      patterns[33417] = 25'b10000010_10000111_00001001_1;
      patterns[33418] = 25'b10000010_10001000_00001010_1;
      patterns[33419] = 25'b10000010_10001001_00001011_1;
      patterns[33420] = 25'b10000010_10001010_00001100_1;
      patterns[33421] = 25'b10000010_10001011_00001101_1;
      patterns[33422] = 25'b10000010_10001100_00001110_1;
      patterns[33423] = 25'b10000010_10001101_00001111_1;
      patterns[33424] = 25'b10000010_10001110_00010000_1;
      patterns[33425] = 25'b10000010_10001111_00010001_1;
      patterns[33426] = 25'b10000010_10010000_00010010_1;
      patterns[33427] = 25'b10000010_10010001_00010011_1;
      patterns[33428] = 25'b10000010_10010010_00010100_1;
      patterns[33429] = 25'b10000010_10010011_00010101_1;
      patterns[33430] = 25'b10000010_10010100_00010110_1;
      patterns[33431] = 25'b10000010_10010101_00010111_1;
      patterns[33432] = 25'b10000010_10010110_00011000_1;
      patterns[33433] = 25'b10000010_10010111_00011001_1;
      patterns[33434] = 25'b10000010_10011000_00011010_1;
      patterns[33435] = 25'b10000010_10011001_00011011_1;
      patterns[33436] = 25'b10000010_10011010_00011100_1;
      patterns[33437] = 25'b10000010_10011011_00011101_1;
      patterns[33438] = 25'b10000010_10011100_00011110_1;
      patterns[33439] = 25'b10000010_10011101_00011111_1;
      patterns[33440] = 25'b10000010_10011110_00100000_1;
      patterns[33441] = 25'b10000010_10011111_00100001_1;
      patterns[33442] = 25'b10000010_10100000_00100010_1;
      patterns[33443] = 25'b10000010_10100001_00100011_1;
      patterns[33444] = 25'b10000010_10100010_00100100_1;
      patterns[33445] = 25'b10000010_10100011_00100101_1;
      patterns[33446] = 25'b10000010_10100100_00100110_1;
      patterns[33447] = 25'b10000010_10100101_00100111_1;
      patterns[33448] = 25'b10000010_10100110_00101000_1;
      patterns[33449] = 25'b10000010_10100111_00101001_1;
      patterns[33450] = 25'b10000010_10101000_00101010_1;
      patterns[33451] = 25'b10000010_10101001_00101011_1;
      patterns[33452] = 25'b10000010_10101010_00101100_1;
      patterns[33453] = 25'b10000010_10101011_00101101_1;
      patterns[33454] = 25'b10000010_10101100_00101110_1;
      patterns[33455] = 25'b10000010_10101101_00101111_1;
      patterns[33456] = 25'b10000010_10101110_00110000_1;
      patterns[33457] = 25'b10000010_10101111_00110001_1;
      patterns[33458] = 25'b10000010_10110000_00110010_1;
      patterns[33459] = 25'b10000010_10110001_00110011_1;
      patterns[33460] = 25'b10000010_10110010_00110100_1;
      patterns[33461] = 25'b10000010_10110011_00110101_1;
      patterns[33462] = 25'b10000010_10110100_00110110_1;
      patterns[33463] = 25'b10000010_10110101_00110111_1;
      patterns[33464] = 25'b10000010_10110110_00111000_1;
      patterns[33465] = 25'b10000010_10110111_00111001_1;
      patterns[33466] = 25'b10000010_10111000_00111010_1;
      patterns[33467] = 25'b10000010_10111001_00111011_1;
      patterns[33468] = 25'b10000010_10111010_00111100_1;
      patterns[33469] = 25'b10000010_10111011_00111101_1;
      patterns[33470] = 25'b10000010_10111100_00111110_1;
      patterns[33471] = 25'b10000010_10111101_00111111_1;
      patterns[33472] = 25'b10000010_10111110_01000000_1;
      patterns[33473] = 25'b10000010_10111111_01000001_1;
      patterns[33474] = 25'b10000010_11000000_01000010_1;
      patterns[33475] = 25'b10000010_11000001_01000011_1;
      patterns[33476] = 25'b10000010_11000010_01000100_1;
      patterns[33477] = 25'b10000010_11000011_01000101_1;
      patterns[33478] = 25'b10000010_11000100_01000110_1;
      patterns[33479] = 25'b10000010_11000101_01000111_1;
      patterns[33480] = 25'b10000010_11000110_01001000_1;
      patterns[33481] = 25'b10000010_11000111_01001001_1;
      patterns[33482] = 25'b10000010_11001000_01001010_1;
      patterns[33483] = 25'b10000010_11001001_01001011_1;
      patterns[33484] = 25'b10000010_11001010_01001100_1;
      patterns[33485] = 25'b10000010_11001011_01001101_1;
      patterns[33486] = 25'b10000010_11001100_01001110_1;
      patterns[33487] = 25'b10000010_11001101_01001111_1;
      patterns[33488] = 25'b10000010_11001110_01010000_1;
      patterns[33489] = 25'b10000010_11001111_01010001_1;
      patterns[33490] = 25'b10000010_11010000_01010010_1;
      patterns[33491] = 25'b10000010_11010001_01010011_1;
      patterns[33492] = 25'b10000010_11010010_01010100_1;
      patterns[33493] = 25'b10000010_11010011_01010101_1;
      patterns[33494] = 25'b10000010_11010100_01010110_1;
      patterns[33495] = 25'b10000010_11010101_01010111_1;
      patterns[33496] = 25'b10000010_11010110_01011000_1;
      patterns[33497] = 25'b10000010_11010111_01011001_1;
      patterns[33498] = 25'b10000010_11011000_01011010_1;
      patterns[33499] = 25'b10000010_11011001_01011011_1;
      patterns[33500] = 25'b10000010_11011010_01011100_1;
      patterns[33501] = 25'b10000010_11011011_01011101_1;
      patterns[33502] = 25'b10000010_11011100_01011110_1;
      patterns[33503] = 25'b10000010_11011101_01011111_1;
      patterns[33504] = 25'b10000010_11011110_01100000_1;
      patterns[33505] = 25'b10000010_11011111_01100001_1;
      patterns[33506] = 25'b10000010_11100000_01100010_1;
      patterns[33507] = 25'b10000010_11100001_01100011_1;
      patterns[33508] = 25'b10000010_11100010_01100100_1;
      patterns[33509] = 25'b10000010_11100011_01100101_1;
      patterns[33510] = 25'b10000010_11100100_01100110_1;
      patterns[33511] = 25'b10000010_11100101_01100111_1;
      patterns[33512] = 25'b10000010_11100110_01101000_1;
      patterns[33513] = 25'b10000010_11100111_01101001_1;
      patterns[33514] = 25'b10000010_11101000_01101010_1;
      patterns[33515] = 25'b10000010_11101001_01101011_1;
      patterns[33516] = 25'b10000010_11101010_01101100_1;
      patterns[33517] = 25'b10000010_11101011_01101101_1;
      patterns[33518] = 25'b10000010_11101100_01101110_1;
      patterns[33519] = 25'b10000010_11101101_01101111_1;
      patterns[33520] = 25'b10000010_11101110_01110000_1;
      patterns[33521] = 25'b10000010_11101111_01110001_1;
      patterns[33522] = 25'b10000010_11110000_01110010_1;
      patterns[33523] = 25'b10000010_11110001_01110011_1;
      patterns[33524] = 25'b10000010_11110010_01110100_1;
      patterns[33525] = 25'b10000010_11110011_01110101_1;
      patterns[33526] = 25'b10000010_11110100_01110110_1;
      patterns[33527] = 25'b10000010_11110101_01110111_1;
      patterns[33528] = 25'b10000010_11110110_01111000_1;
      patterns[33529] = 25'b10000010_11110111_01111001_1;
      patterns[33530] = 25'b10000010_11111000_01111010_1;
      patterns[33531] = 25'b10000010_11111001_01111011_1;
      patterns[33532] = 25'b10000010_11111010_01111100_1;
      patterns[33533] = 25'b10000010_11111011_01111101_1;
      patterns[33534] = 25'b10000010_11111100_01111110_1;
      patterns[33535] = 25'b10000010_11111101_01111111_1;
      patterns[33536] = 25'b10000010_11111110_10000000_1;
      patterns[33537] = 25'b10000010_11111111_10000001_1;
      patterns[33538] = 25'b10000011_00000000_10000011_0;
      patterns[33539] = 25'b10000011_00000001_10000100_0;
      patterns[33540] = 25'b10000011_00000010_10000101_0;
      patterns[33541] = 25'b10000011_00000011_10000110_0;
      patterns[33542] = 25'b10000011_00000100_10000111_0;
      patterns[33543] = 25'b10000011_00000101_10001000_0;
      patterns[33544] = 25'b10000011_00000110_10001001_0;
      patterns[33545] = 25'b10000011_00000111_10001010_0;
      patterns[33546] = 25'b10000011_00001000_10001011_0;
      patterns[33547] = 25'b10000011_00001001_10001100_0;
      patterns[33548] = 25'b10000011_00001010_10001101_0;
      patterns[33549] = 25'b10000011_00001011_10001110_0;
      patterns[33550] = 25'b10000011_00001100_10001111_0;
      patterns[33551] = 25'b10000011_00001101_10010000_0;
      patterns[33552] = 25'b10000011_00001110_10010001_0;
      patterns[33553] = 25'b10000011_00001111_10010010_0;
      patterns[33554] = 25'b10000011_00010000_10010011_0;
      patterns[33555] = 25'b10000011_00010001_10010100_0;
      patterns[33556] = 25'b10000011_00010010_10010101_0;
      patterns[33557] = 25'b10000011_00010011_10010110_0;
      patterns[33558] = 25'b10000011_00010100_10010111_0;
      patterns[33559] = 25'b10000011_00010101_10011000_0;
      patterns[33560] = 25'b10000011_00010110_10011001_0;
      patterns[33561] = 25'b10000011_00010111_10011010_0;
      patterns[33562] = 25'b10000011_00011000_10011011_0;
      patterns[33563] = 25'b10000011_00011001_10011100_0;
      patterns[33564] = 25'b10000011_00011010_10011101_0;
      patterns[33565] = 25'b10000011_00011011_10011110_0;
      patterns[33566] = 25'b10000011_00011100_10011111_0;
      patterns[33567] = 25'b10000011_00011101_10100000_0;
      patterns[33568] = 25'b10000011_00011110_10100001_0;
      patterns[33569] = 25'b10000011_00011111_10100010_0;
      patterns[33570] = 25'b10000011_00100000_10100011_0;
      patterns[33571] = 25'b10000011_00100001_10100100_0;
      patterns[33572] = 25'b10000011_00100010_10100101_0;
      patterns[33573] = 25'b10000011_00100011_10100110_0;
      patterns[33574] = 25'b10000011_00100100_10100111_0;
      patterns[33575] = 25'b10000011_00100101_10101000_0;
      patterns[33576] = 25'b10000011_00100110_10101001_0;
      patterns[33577] = 25'b10000011_00100111_10101010_0;
      patterns[33578] = 25'b10000011_00101000_10101011_0;
      patterns[33579] = 25'b10000011_00101001_10101100_0;
      patterns[33580] = 25'b10000011_00101010_10101101_0;
      patterns[33581] = 25'b10000011_00101011_10101110_0;
      patterns[33582] = 25'b10000011_00101100_10101111_0;
      patterns[33583] = 25'b10000011_00101101_10110000_0;
      patterns[33584] = 25'b10000011_00101110_10110001_0;
      patterns[33585] = 25'b10000011_00101111_10110010_0;
      patterns[33586] = 25'b10000011_00110000_10110011_0;
      patterns[33587] = 25'b10000011_00110001_10110100_0;
      patterns[33588] = 25'b10000011_00110010_10110101_0;
      patterns[33589] = 25'b10000011_00110011_10110110_0;
      patterns[33590] = 25'b10000011_00110100_10110111_0;
      patterns[33591] = 25'b10000011_00110101_10111000_0;
      patterns[33592] = 25'b10000011_00110110_10111001_0;
      patterns[33593] = 25'b10000011_00110111_10111010_0;
      patterns[33594] = 25'b10000011_00111000_10111011_0;
      patterns[33595] = 25'b10000011_00111001_10111100_0;
      patterns[33596] = 25'b10000011_00111010_10111101_0;
      patterns[33597] = 25'b10000011_00111011_10111110_0;
      patterns[33598] = 25'b10000011_00111100_10111111_0;
      patterns[33599] = 25'b10000011_00111101_11000000_0;
      patterns[33600] = 25'b10000011_00111110_11000001_0;
      patterns[33601] = 25'b10000011_00111111_11000010_0;
      patterns[33602] = 25'b10000011_01000000_11000011_0;
      patterns[33603] = 25'b10000011_01000001_11000100_0;
      patterns[33604] = 25'b10000011_01000010_11000101_0;
      patterns[33605] = 25'b10000011_01000011_11000110_0;
      patterns[33606] = 25'b10000011_01000100_11000111_0;
      patterns[33607] = 25'b10000011_01000101_11001000_0;
      patterns[33608] = 25'b10000011_01000110_11001001_0;
      patterns[33609] = 25'b10000011_01000111_11001010_0;
      patterns[33610] = 25'b10000011_01001000_11001011_0;
      patterns[33611] = 25'b10000011_01001001_11001100_0;
      patterns[33612] = 25'b10000011_01001010_11001101_0;
      patterns[33613] = 25'b10000011_01001011_11001110_0;
      patterns[33614] = 25'b10000011_01001100_11001111_0;
      patterns[33615] = 25'b10000011_01001101_11010000_0;
      patterns[33616] = 25'b10000011_01001110_11010001_0;
      patterns[33617] = 25'b10000011_01001111_11010010_0;
      patterns[33618] = 25'b10000011_01010000_11010011_0;
      patterns[33619] = 25'b10000011_01010001_11010100_0;
      patterns[33620] = 25'b10000011_01010010_11010101_0;
      patterns[33621] = 25'b10000011_01010011_11010110_0;
      patterns[33622] = 25'b10000011_01010100_11010111_0;
      patterns[33623] = 25'b10000011_01010101_11011000_0;
      patterns[33624] = 25'b10000011_01010110_11011001_0;
      patterns[33625] = 25'b10000011_01010111_11011010_0;
      patterns[33626] = 25'b10000011_01011000_11011011_0;
      patterns[33627] = 25'b10000011_01011001_11011100_0;
      patterns[33628] = 25'b10000011_01011010_11011101_0;
      patterns[33629] = 25'b10000011_01011011_11011110_0;
      patterns[33630] = 25'b10000011_01011100_11011111_0;
      patterns[33631] = 25'b10000011_01011101_11100000_0;
      patterns[33632] = 25'b10000011_01011110_11100001_0;
      patterns[33633] = 25'b10000011_01011111_11100010_0;
      patterns[33634] = 25'b10000011_01100000_11100011_0;
      patterns[33635] = 25'b10000011_01100001_11100100_0;
      patterns[33636] = 25'b10000011_01100010_11100101_0;
      patterns[33637] = 25'b10000011_01100011_11100110_0;
      patterns[33638] = 25'b10000011_01100100_11100111_0;
      patterns[33639] = 25'b10000011_01100101_11101000_0;
      patterns[33640] = 25'b10000011_01100110_11101001_0;
      patterns[33641] = 25'b10000011_01100111_11101010_0;
      patterns[33642] = 25'b10000011_01101000_11101011_0;
      patterns[33643] = 25'b10000011_01101001_11101100_0;
      patterns[33644] = 25'b10000011_01101010_11101101_0;
      patterns[33645] = 25'b10000011_01101011_11101110_0;
      patterns[33646] = 25'b10000011_01101100_11101111_0;
      patterns[33647] = 25'b10000011_01101101_11110000_0;
      patterns[33648] = 25'b10000011_01101110_11110001_0;
      patterns[33649] = 25'b10000011_01101111_11110010_0;
      patterns[33650] = 25'b10000011_01110000_11110011_0;
      patterns[33651] = 25'b10000011_01110001_11110100_0;
      patterns[33652] = 25'b10000011_01110010_11110101_0;
      patterns[33653] = 25'b10000011_01110011_11110110_0;
      patterns[33654] = 25'b10000011_01110100_11110111_0;
      patterns[33655] = 25'b10000011_01110101_11111000_0;
      patterns[33656] = 25'b10000011_01110110_11111001_0;
      patterns[33657] = 25'b10000011_01110111_11111010_0;
      patterns[33658] = 25'b10000011_01111000_11111011_0;
      patterns[33659] = 25'b10000011_01111001_11111100_0;
      patterns[33660] = 25'b10000011_01111010_11111101_0;
      patterns[33661] = 25'b10000011_01111011_11111110_0;
      patterns[33662] = 25'b10000011_01111100_11111111_0;
      patterns[33663] = 25'b10000011_01111101_00000000_1;
      patterns[33664] = 25'b10000011_01111110_00000001_1;
      patterns[33665] = 25'b10000011_01111111_00000010_1;
      patterns[33666] = 25'b10000011_10000000_00000011_1;
      patterns[33667] = 25'b10000011_10000001_00000100_1;
      patterns[33668] = 25'b10000011_10000010_00000101_1;
      patterns[33669] = 25'b10000011_10000011_00000110_1;
      patterns[33670] = 25'b10000011_10000100_00000111_1;
      patterns[33671] = 25'b10000011_10000101_00001000_1;
      patterns[33672] = 25'b10000011_10000110_00001001_1;
      patterns[33673] = 25'b10000011_10000111_00001010_1;
      patterns[33674] = 25'b10000011_10001000_00001011_1;
      patterns[33675] = 25'b10000011_10001001_00001100_1;
      patterns[33676] = 25'b10000011_10001010_00001101_1;
      patterns[33677] = 25'b10000011_10001011_00001110_1;
      patterns[33678] = 25'b10000011_10001100_00001111_1;
      patterns[33679] = 25'b10000011_10001101_00010000_1;
      patterns[33680] = 25'b10000011_10001110_00010001_1;
      patterns[33681] = 25'b10000011_10001111_00010010_1;
      patterns[33682] = 25'b10000011_10010000_00010011_1;
      patterns[33683] = 25'b10000011_10010001_00010100_1;
      patterns[33684] = 25'b10000011_10010010_00010101_1;
      patterns[33685] = 25'b10000011_10010011_00010110_1;
      patterns[33686] = 25'b10000011_10010100_00010111_1;
      patterns[33687] = 25'b10000011_10010101_00011000_1;
      patterns[33688] = 25'b10000011_10010110_00011001_1;
      patterns[33689] = 25'b10000011_10010111_00011010_1;
      patterns[33690] = 25'b10000011_10011000_00011011_1;
      patterns[33691] = 25'b10000011_10011001_00011100_1;
      patterns[33692] = 25'b10000011_10011010_00011101_1;
      patterns[33693] = 25'b10000011_10011011_00011110_1;
      patterns[33694] = 25'b10000011_10011100_00011111_1;
      patterns[33695] = 25'b10000011_10011101_00100000_1;
      patterns[33696] = 25'b10000011_10011110_00100001_1;
      patterns[33697] = 25'b10000011_10011111_00100010_1;
      patterns[33698] = 25'b10000011_10100000_00100011_1;
      patterns[33699] = 25'b10000011_10100001_00100100_1;
      patterns[33700] = 25'b10000011_10100010_00100101_1;
      patterns[33701] = 25'b10000011_10100011_00100110_1;
      patterns[33702] = 25'b10000011_10100100_00100111_1;
      patterns[33703] = 25'b10000011_10100101_00101000_1;
      patterns[33704] = 25'b10000011_10100110_00101001_1;
      patterns[33705] = 25'b10000011_10100111_00101010_1;
      patterns[33706] = 25'b10000011_10101000_00101011_1;
      patterns[33707] = 25'b10000011_10101001_00101100_1;
      patterns[33708] = 25'b10000011_10101010_00101101_1;
      patterns[33709] = 25'b10000011_10101011_00101110_1;
      patterns[33710] = 25'b10000011_10101100_00101111_1;
      patterns[33711] = 25'b10000011_10101101_00110000_1;
      patterns[33712] = 25'b10000011_10101110_00110001_1;
      patterns[33713] = 25'b10000011_10101111_00110010_1;
      patterns[33714] = 25'b10000011_10110000_00110011_1;
      patterns[33715] = 25'b10000011_10110001_00110100_1;
      patterns[33716] = 25'b10000011_10110010_00110101_1;
      patterns[33717] = 25'b10000011_10110011_00110110_1;
      patterns[33718] = 25'b10000011_10110100_00110111_1;
      patterns[33719] = 25'b10000011_10110101_00111000_1;
      patterns[33720] = 25'b10000011_10110110_00111001_1;
      patterns[33721] = 25'b10000011_10110111_00111010_1;
      patterns[33722] = 25'b10000011_10111000_00111011_1;
      patterns[33723] = 25'b10000011_10111001_00111100_1;
      patterns[33724] = 25'b10000011_10111010_00111101_1;
      patterns[33725] = 25'b10000011_10111011_00111110_1;
      patterns[33726] = 25'b10000011_10111100_00111111_1;
      patterns[33727] = 25'b10000011_10111101_01000000_1;
      patterns[33728] = 25'b10000011_10111110_01000001_1;
      patterns[33729] = 25'b10000011_10111111_01000010_1;
      patterns[33730] = 25'b10000011_11000000_01000011_1;
      patterns[33731] = 25'b10000011_11000001_01000100_1;
      patterns[33732] = 25'b10000011_11000010_01000101_1;
      patterns[33733] = 25'b10000011_11000011_01000110_1;
      patterns[33734] = 25'b10000011_11000100_01000111_1;
      patterns[33735] = 25'b10000011_11000101_01001000_1;
      patterns[33736] = 25'b10000011_11000110_01001001_1;
      patterns[33737] = 25'b10000011_11000111_01001010_1;
      patterns[33738] = 25'b10000011_11001000_01001011_1;
      patterns[33739] = 25'b10000011_11001001_01001100_1;
      patterns[33740] = 25'b10000011_11001010_01001101_1;
      patterns[33741] = 25'b10000011_11001011_01001110_1;
      patterns[33742] = 25'b10000011_11001100_01001111_1;
      patterns[33743] = 25'b10000011_11001101_01010000_1;
      patterns[33744] = 25'b10000011_11001110_01010001_1;
      patterns[33745] = 25'b10000011_11001111_01010010_1;
      patterns[33746] = 25'b10000011_11010000_01010011_1;
      patterns[33747] = 25'b10000011_11010001_01010100_1;
      patterns[33748] = 25'b10000011_11010010_01010101_1;
      patterns[33749] = 25'b10000011_11010011_01010110_1;
      patterns[33750] = 25'b10000011_11010100_01010111_1;
      patterns[33751] = 25'b10000011_11010101_01011000_1;
      patterns[33752] = 25'b10000011_11010110_01011001_1;
      patterns[33753] = 25'b10000011_11010111_01011010_1;
      patterns[33754] = 25'b10000011_11011000_01011011_1;
      patterns[33755] = 25'b10000011_11011001_01011100_1;
      patterns[33756] = 25'b10000011_11011010_01011101_1;
      patterns[33757] = 25'b10000011_11011011_01011110_1;
      patterns[33758] = 25'b10000011_11011100_01011111_1;
      patterns[33759] = 25'b10000011_11011101_01100000_1;
      patterns[33760] = 25'b10000011_11011110_01100001_1;
      patterns[33761] = 25'b10000011_11011111_01100010_1;
      patterns[33762] = 25'b10000011_11100000_01100011_1;
      patterns[33763] = 25'b10000011_11100001_01100100_1;
      patterns[33764] = 25'b10000011_11100010_01100101_1;
      patterns[33765] = 25'b10000011_11100011_01100110_1;
      patterns[33766] = 25'b10000011_11100100_01100111_1;
      patterns[33767] = 25'b10000011_11100101_01101000_1;
      patterns[33768] = 25'b10000011_11100110_01101001_1;
      patterns[33769] = 25'b10000011_11100111_01101010_1;
      patterns[33770] = 25'b10000011_11101000_01101011_1;
      patterns[33771] = 25'b10000011_11101001_01101100_1;
      patterns[33772] = 25'b10000011_11101010_01101101_1;
      patterns[33773] = 25'b10000011_11101011_01101110_1;
      patterns[33774] = 25'b10000011_11101100_01101111_1;
      patterns[33775] = 25'b10000011_11101101_01110000_1;
      patterns[33776] = 25'b10000011_11101110_01110001_1;
      patterns[33777] = 25'b10000011_11101111_01110010_1;
      patterns[33778] = 25'b10000011_11110000_01110011_1;
      patterns[33779] = 25'b10000011_11110001_01110100_1;
      patterns[33780] = 25'b10000011_11110010_01110101_1;
      patterns[33781] = 25'b10000011_11110011_01110110_1;
      patterns[33782] = 25'b10000011_11110100_01110111_1;
      patterns[33783] = 25'b10000011_11110101_01111000_1;
      patterns[33784] = 25'b10000011_11110110_01111001_1;
      patterns[33785] = 25'b10000011_11110111_01111010_1;
      patterns[33786] = 25'b10000011_11111000_01111011_1;
      patterns[33787] = 25'b10000011_11111001_01111100_1;
      patterns[33788] = 25'b10000011_11111010_01111101_1;
      patterns[33789] = 25'b10000011_11111011_01111110_1;
      patterns[33790] = 25'b10000011_11111100_01111111_1;
      patterns[33791] = 25'b10000011_11111101_10000000_1;
      patterns[33792] = 25'b10000011_11111110_10000001_1;
      patterns[33793] = 25'b10000011_11111111_10000010_1;
      patterns[33794] = 25'b10000100_00000000_10000100_0;
      patterns[33795] = 25'b10000100_00000001_10000101_0;
      patterns[33796] = 25'b10000100_00000010_10000110_0;
      patterns[33797] = 25'b10000100_00000011_10000111_0;
      patterns[33798] = 25'b10000100_00000100_10001000_0;
      patterns[33799] = 25'b10000100_00000101_10001001_0;
      patterns[33800] = 25'b10000100_00000110_10001010_0;
      patterns[33801] = 25'b10000100_00000111_10001011_0;
      patterns[33802] = 25'b10000100_00001000_10001100_0;
      patterns[33803] = 25'b10000100_00001001_10001101_0;
      patterns[33804] = 25'b10000100_00001010_10001110_0;
      patterns[33805] = 25'b10000100_00001011_10001111_0;
      patterns[33806] = 25'b10000100_00001100_10010000_0;
      patterns[33807] = 25'b10000100_00001101_10010001_0;
      patterns[33808] = 25'b10000100_00001110_10010010_0;
      patterns[33809] = 25'b10000100_00001111_10010011_0;
      patterns[33810] = 25'b10000100_00010000_10010100_0;
      patterns[33811] = 25'b10000100_00010001_10010101_0;
      patterns[33812] = 25'b10000100_00010010_10010110_0;
      patterns[33813] = 25'b10000100_00010011_10010111_0;
      patterns[33814] = 25'b10000100_00010100_10011000_0;
      patterns[33815] = 25'b10000100_00010101_10011001_0;
      patterns[33816] = 25'b10000100_00010110_10011010_0;
      patterns[33817] = 25'b10000100_00010111_10011011_0;
      patterns[33818] = 25'b10000100_00011000_10011100_0;
      patterns[33819] = 25'b10000100_00011001_10011101_0;
      patterns[33820] = 25'b10000100_00011010_10011110_0;
      patterns[33821] = 25'b10000100_00011011_10011111_0;
      patterns[33822] = 25'b10000100_00011100_10100000_0;
      patterns[33823] = 25'b10000100_00011101_10100001_0;
      patterns[33824] = 25'b10000100_00011110_10100010_0;
      patterns[33825] = 25'b10000100_00011111_10100011_0;
      patterns[33826] = 25'b10000100_00100000_10100100_0;
      patterns[33827] = 25'b10000100_00100001_10100101_0;
      patterns[33828] = 25'b10000100_00100010_10100110_0;
      patterns[33829] = 25'b10000100_00100011_10100111_0;
      patterns[33830] = 25'b10000100_00100100_10101000_0;
      patterns[33831] = 25'b10000100_00100101_10101001_0;
      patterns[33832] = 25'b10000100_00100110_10101010_0;
      patterns[33833] = 25'b10000100_00100111_10101011_0;
      patterns[33834] = 25'b10000100_00101000_10101100_0;
      patterns[33835] = 25'b10000100_00101001_10101101_0;
      patterns[33836] = 25'b10000100_00101010_10101110_0;
      patterns[33837] = 25'b10000100_00101011_10101111_0;
      patterns[33838] = 25'b10000100_00101100_10110000_0;
      patterns[33839] = 25'b10000100_00101101_10110001_0;
      patterns[33840] = 25'b10000100_00101110_10110010_0;
      patterns[33841] = 25'b10000100_00101111_10110011_0;
      patterns[33842] = 25'b10000100_00110000_10110100_0;
      patterns[33843] = 25'b10000100_00110001_10110101_0;
      patterns[33844] = 25'b10000100_00110010_10110110_0;
      patterns[33845] = 25'b10000100_00110011_10110111_0;
      patterns[33846] = 25'b10000100_00110100_10111000_0;
      patterns[33847] = 25'b10000100_00110101_10111001_0;
      patterns[33848] = 25'b10000100_00110110_10111010_0;
      patterns[33849] = 25'b10000100_00110111_10111011_0;
      patterns[33850] = 25'b10000100_00111000_10111100_0;
      patterns[33851] = 25'b10000100_00111001_10111101_0;
      patterns[33852] = 25'b10000100_00111010_10111110_0;
      patterns[33853] = 25'b10000100_00111011_10111111_0;
      patterns[33854] = 25'b10000100_00111100_11000000_0;
      patterns[33855] = 25'b10000100_00111101_11000001_0;
      patterns[33856] = 25'b10000100_00111110_11000010_0;
      patterns[33857] = 25'b10000100_00111111_11000011_0;
      patterns[33858] = 25'b10000100_01000000_11000100_0;
      patterns[33859] = 25'b10000100_01000001_11000101_0;
      patterns[33860] = 25'b10000100_01000010_11000110_0;
      patterns[33861] = 25'b10000100_01000011_11000111_0;
      patterns[33862] = 25'b10000100_01000100_11001000_0;
      patterns[33863] = 25'b10000100_01000101_11001001_0;
      patterns[33864] = 25'b10000100_01000110_11001010_0;
      patterns[33865] = 25'b10000100_01000111_11001011_0;
      patterns[33866] = 25'b10000100_01001000_11001100_0;
      patterns[33867] = 25'b10000100_01001001_11001101_0;
      patterns[33868] = 25'b10000100_01001010_11001110_0;
      patterns[33869] = 25'b10000100_01001011_11001111_0;
      patterns[33870] = 25'b10000100_01001100_11010000_0;
      patterns[33871] = 25'b10000100_01001101_11010001_0;
      patterns[33872] = 25'b10000100_01001110_11010010_0;
      patterns[33873] = 25'b10000100_01001111_11010011_0;
      patterns[33874] = 25'b10000100_01010000_11010100_0;
      patterns[33875] = 25'b10000100_01010001_11010101_0;
      patterns[33876] = 25'b10000100_01010010_11010110_0;
      patterns[33877] = 25'b10000100_01010011_11010111_0;
      patterns[33878] = 25'b10000100_01010100_11011000_0;
      patterns[33879] = 25'b10000100_01010101_11011001_0;
      patterns[33880] = 25'b10000100_01010110_11011010_0;
      patterns[33881] = 25'b10000100_01010111_11011011_0;
      patterns[33882] = 25'b10000100_01011000_11011100_0;
      patterns[33883] = 25'b10000100_01011001_11011101_0;
      patterns[33884] = 25'b10000100_01011010_11011110_0;
      patterns[33885] = 25'b10000100_01011011_11011111_0;
      patterns[33886] = 25'b10000100_01011100_11100000_0;
      patterns[33887] = 25'b10000100_01011101_11100001_0;
      patterns[33888] = 25'b10000100_01011110_11100010_0;
      patterns[33889] = 25'b10000100_01011111_11100011_0;
      patterns[33890] = 25'b10000100_01100000_11100100_0;
      patterns[33891] = 25'b10000100_01100001_11100101_0;
      patterns[33892] = 25'b10000100_01100010_11100110_0;
      patterns[33893] = 25'b10000100_01100011_11100111_0;
      patterns[33894] = 25'b10000100_01100100_11101000_0;
      patterns[33895] = 25'b10000100_01100101_11101001_0;
      patterns[33896] = 25'b10000100_01100110_11101010_0;
      patterns[33897] = 25'b10000100_01100111_11101011_0;
      patterns[33898] = 25'b10000100_01101000_11101100_0;
      patterns[33899] = 25'b10000100_01101001_11101101_0;
      patterns[33900] = 25'b10000100_01101010_11101110_0;
      patterns[33901] = 25'b10000100_01101011_11101111_0;
      patterns[33902] = 25'b10000100_01101100_11110000_0;
      patterns[33903] = 25'b10000100_01101101_11110001_0;
      patterns[33904] = 25'b10000100_01101110_11110010_0;
      patterns[33905] = 25'b10000100_01101111_11110011_0;
      patterns[33906] = 25'b10000100_01110000_11110100_0;
      patterns[33907] = 25'b10000100_01110001_11110101_0;
      patterns[33908] = 25'b10000100_01110010_11110110_0;
      patterns[33909] = 25'b10000100_01110011_11110111_0;
      patterns[33910] = 25'b10000100_01110100_11111000_0;
      patterns[33911] = 25'b10000100_01110101_11111001_0;
      patterns[33912] = 25'b10000100_01110110_11111010_0;
      patterns[33913] = 25'b10000100_01110111_11111011_0;
      patterns[33914] = 25'b10000100_01111000_11111100_0;
      patterns[33915] = 25'b10000100_01111001_11111101_0;
      patterns[33916] = 25'b10000100_01111010_11111110_0;
      patterns[33917] = 25'b10000100_01111011_11111111_0;
      patterns[33918] = 25'b10000100_01111100_00000000_1;
      patterns[33919] = 25'b10000100_01111101_00000001_1;
      patterns[33920] = 25'b10000100_01111110_00000010_1;
      patterns[33921] = 25'b10000100_01111111_00000011_1;
      patterns[33922] = 25'b10000100_10000000_00000100_1;
      patterns[33923] = 25'b10000100_10000001_00000101_1;
      patterns[33924] = 25'b10000100_10000010_00000110_1;
      patterns[33925] = 25'b10000100_10000011_00000111_1;
      patterns[33926] = 25'b10000100_10000100_00001000_1;
      patterns[33927] = 25'b10000100_10000101_00001001_1;
      patterns[33928] = 25'b10000100_10000110_00001010_1;
      patterns[33929] = 25'b10000100_10000111_00001011_1;
      patterns[33930] = 25'b10000100_10001000_00001100_1;
      patterns[33931] = 25'b10000100_10001001_00001101_1;
      patterns[33932] = 25'b10000100_10001010_00001110_1;
      patterns[33933] = 25'b10000100_10001011_00001111_1;
      patterns[33934] = 25'b10000100_10001100_00010000_1;
      patterns[33935] = 25'b10000100_10001101_00010001_1;
      patterns[33936] = 25'b10000100_10001110_00010010_1;
      patterns[33937] = 25'b10000100_10001111_00010011_1;
      patterns[33938] = 25'b10000100_10010000_00010100_1;
      patterns[33939] = 25'b10000100_10010001_00010101_1;
      patterns[33940] = 25'b10000100_10010010_00010110_1;
      patterns[33941] = 25'b10000100_10010011_00010111_1;
      patterns[33942] = 25'b10000100_10010100_00011000_1;
      patterns[33943] = 25'b10000100_10010101_00011001_1;
      patterns[33944] = 25'b10000100_10010110_00011010_1;
      patterns[33945] = 25'b10000100_10010111_00011011_1;
      patterns[33946] = 25'b10000100_10011000_00011100_1;
      patterns[33947] = 25'b10000100_10011001_00011101_1;
      patterns[33948] = 25'b10000100_10011010_00011110_1;
      patterns[33949] = 25'b10000100_10011011_00011111_1;
      patterns[33950] = 25'b10000100_10011100_00100000_1;
      patterns[33951] = 25'b10000100_10011101_00100001_1;
      patterns[33952] = 25'b10000100_10011110_00100010_1;
      patterns[33953] = 25'b10000100_10011111_00100011_1;
      patterns[33954] = 25'b10000100_10100000_00100100_1;
      patterns[33955] = 25'b10000100_10100001_00100101_1;
      patterns[33956] = 25'b10000100_10100010_00100110_1;
      patterns[33957] = 25'b10000100_10100011_00100111_1;
      patterns[33958] = 25'b10000100_10100100_00101000_1;
      patterns[33959] = 25'b10000100_10100101_00101001_1;
      patterns[33960] = 25'b10000100_10100110_00101010_1;
      patterns[33961] = 25'b10000100_10100111_00101011_1;
      patterns[33962] = 25'b10000100_10101000_00101100_1;
      patterns[33963] = 25'b10000100_10101001_00101101_1;
      patterns[33964] = 25'b10000100_10101010_00101110_1;
      patterns[33965] = 25'b10000100_10101011_00101111_1;
      patterns[33966] = 25'b10000100_10101100_00110000_1;
      patterns[33967] = 25'b10000100_10101101_00110001_1;
      patterns[33968] = 25'b10000100_10101110_00110010_1;
      patterns[33969] = 25'b10000100_10101111_00110011_1;
      patterns[33970] = 25'b10000100_10110000_00110100_1;
      patterns[33971] = 25'b10000100_10110001_00110101_1;
      patterns[33972] = 25'b10000100_10110010_00110110_1;
      patterns[33973] = 25'b10000100_10110011_00110111_1;
      patterns[33974] = 25'b10000100_10110100_00111000_1;
      patterns[33975] = 25'b10000100_10110101_00111001_1;
      patterns[33976] = 25'b10000100_10110110_00111010_1;
      patterns[33977] = 25'b10000100_10110111_00111011_1;
      patterns[33978] = 25'b10000100_10111000_00111100_1;
      patterns[33979] = 25'b10000100_10111001_00111101_1;
      patterns[33980] = 25'b10000100_10111010_00111110_1;
      patterns[33981] = 25'b10000100_10111011_00111111_1;
      patterns[33982] = 25'b10000100_10111100_01000000_1;
      patterns[33983] = 25'b10000100_10111101_01000001_1;
      patterns[33984] = 25'b10000100_10111110_01000010_1;
      patterns[33985] = 25'b10000100_10111111_01000011_1;
      patterns[33986] = 25'b10000100_11000000_01000100_1;
      patterns[33987] = 25'b10000100_11000001_01000101_1;
      patterns[33988] = 25'b10000100_11000010_01000110_1;
      patterns[33989] = 25'b10000100_11000011_01000111_1;
      patterns[33990] = 25'b10000100_11000100_01001000_1;
      patterns[33991] = 25'b10000100_11000101_01001001_1;
      patterns[33992] = 25'b10000100_11000110_01001010_1;
      patterns[33993] = 25'b10000100_11000111_01001011_1;
      patterns[33994] = 25'b10000100_11001000_01001100_1;
      patterns[33995] = 25'b10000100_11001001_01001101_1;
      patterns[33996] = 25'b10000100_11001010_01001110_1;
      patterns[33997] = 25'b10000100_11001011_01001111_1;
      patterns[33998] = 25'b10000100_11001100_01010000_1;
      patterns[33999] = 25'b10000100_11001101_01010001_1;
      patterns[34000] = 25'b10000100_11001110_01010010_1;
      patterns[34001] = 25'b10000100_11001111_01010011_1;
      patterns[34002] = 25'b10000100_11010000_01010100_1;
      patterns[34003] = 25'b10000100_11010001_01010101_1;
      patterns[34004] = 25'b10000100_11010010_01010110_1;
      patterns[34005] = 25'b10000100_11010011_01010111_1;
      patterns[34006] = 25'b10000100_11010100_01011000_1;
      patterns[34007] = 25'b10000100_11010101_01011001_1;
      patterns[34008] = 25'b10000100_11010110_01011010_1;
      patterns[34009] = 25'b10000100_11010111_01011011_1;
      patterns[34010] = 25'b10000100_11011000_01011100_1;
      patterns[34011] = 25'b10000100_11011001_01011101_1;
      patterns[34012] = 25'b10000100_11011010_01011110_1;
      patterns[34013] = 25'b10000100_11011011_01011111_1;
      patterns[34014] = 25'b10000100_11011100_01100000_1;
      patterns[34015] = 25'b10000100_11011101_01100001_1;
      patterns[34016] = 25'b10000100_11011110_01100010_1;
      patterns[34017] = 25'b10000100_11011111_01100011_1;
      patterns[34018] = 25'b10000100_11100000_01100100_1;
      patterns[34019] = 25'b10000100_11100001_01100101_1;
      patterns[34020] = 25'b10000100_11100010_01100110_1;
      patterns[34021] = 25'b10000100_11100011_01100111_1;
      patterns[34022] = 25'b10000100_11100100_01101000_1;
      patterns[34023] = 25'b10000100_11100101_01101001_1;
      patterns[34024] = 25'b10000100_11100110_01101010_1;
      patterns[34025] = 25'b10000100_11100111_01101011_1;
      patterns[34026] = 25'b10000100_11101000_01101100_1;
      patterns[34027] = 25'b10000100_11101001_01101101_1;
      patterns[34028] = 25'b10000100_11101010_01101110_1;
      patterns[34029] = 25'b10000100_11101011_01101111_1;
      patterns[34030] = 25'b10000100_11101100_01110000_1;
      patterns[34031] = 25'b10000100_11101101_01110001_1;
      patterns[34032] = 25'b10000100_11101110_01110010_1;
      patterns[34033] = 25'b10000100_11101111_01110011_1;
      patterns[34034] = 25'b10000100_11110000_01110100_1;
      patterns[34035] = 25'b10000100_11110001_01110101_1;
      patterns[34036] = 25'b10000100_11110010_01110110_1;
      patterns[34037] = 25'b10000100_11110011_01110111_1;
      patterns[34038] = 25'b10000100_11110100_01111000_1;
      patterns[34039] = 25'b10000100_11110101_01111001_1;
      patterns[34040] = 25'b10000100_11110110_01111010_1;
      patterns[34041] = 25'b10000100_11110111_01111011_1;
      patterns[34042] = 25'b10000100_11111000_01111100_1;
      patterns[34043] = 25'b10000100_11111001_01111101_1;
      patterns[34044] = 25'b10000100_11111010_01111110_1;
      patterns[34045] = 25'b10000100_11111011_01111111_1;
      patterns[34046] = 25'b10000100_11111100_10000000_1;
      patterns[34047] = 25'b10000100_11111101_10000001_1;
      patterns[34048] = 25'b10000100_11111110_10000010_1;
      patterns[34049] = 25'b10000100_11111111_10000011_1;
      patterns[34050] = 25'b10000101_00000000_10000101_0;
      patterns[34051] = 25'b10000101_00000001_10000110_0;
      patterns[34052] = 25'b10000101_00000010_10000111_0;
      patterns[34053] = 25'b10000101_00000011_10001000_0;
      patterns[34054] = 25'b10000101_00000100_10001001_0;
      patterns[34055] = 25'b10000101_00000101_10001010_0;
      patterns[34056] = 25'b10000101_00000110_10001011_0;
      patterns[34057] = 25'b10000101_00000111_10001100_0;
      patterns[34058] = 25'b10000101_00001000_10001101_0;
      patterns[34059] = 25'b10000101_00001001_10001110_0;
      patterns[34060] = 25'b10000101_00001010_10001111_0;
      patterns[34061] = 25'b10000101_00001011_10010000_0;
      patterns[34062] = 25'b10000101_00001100_10010001_0;
      patterns[34063] = 25'b10000101_00001101_10010010_0;
      patterns[34064] = 25'b10000101_00001110_10010011_0;
      patterns[34065] = 25'b10000101_00001111_10010100_0;
      patterns[34066] = 25'b10000101_00010000_10010101_0;
      patterns[34067] = 25'b10000101_00010001_10010110_0;
      patterns[34068] = 25'b10000101_00010010_10010111_0;
      patterns[34069] = 25'b10000101_00010011_10011000_0;
      patterns[34070] = 25'b10000101_00010100_10011001_0;
      patterns[34071] = 25'b10000101_00010101_10011010_0;
      patterns[34072] = 25'b10000101_00010110_10011011_0;
      patterns[34073] = 25'b10000101_00010111_10011100_0;
      patterns[34074] = 25'b10000101_00011000_10011101_0;
      patterns[34075] = 25'b10000101_00011001_10011110_0;
      patterns[34076] = 25'b10000101_00011010_10011111_0;
      patterns[34077] = 25'b10000101_00011011_10100000_0;
      patterns[34078] = 25'b10000101_00011100_10100001_0;
      patterns[34079] = 25'b10000101_00011101_10100010_0;
      patterns[34080] = 25'b10000101_00011110_10100011_0;
      patterns[34081] = 25'b10000101_00011111_10100100_0;
      patterns[34082] = 25'b10000101_00100000_10100101_0;
      patterns[34083] = 25'b10000101_00100001_10100110_0;
      patterns[34084] = 25'b10000101_00100010_10100111_0;
      patterns[34085] = 25'b10000101_00100011_10101000_0;
      patterns[34086] = 25'b10000101_00100100_10101001_0;
      patterns[34087] = 25'b10000101_00100101_10101010_0;
      patterns[34088] = 25'b10000101_00100110_10101011_0;
      patterns[34089] = 25'b10000101_00100111_10101100_0;
      patterns[34090] = 25'b10000101_00101000_10101101_0;
      patterns[34091] = 25'b10000101_00101001_10101110_0;
      patterns[34092] = 25'b10000101_00101010_10101111_0;
      patterns[34093] = 25'b10000101_00101011_10110000_0;
      patterns[34094] = 25'b10000101_00101100_10110001_0;
      patterns[34095] = 25'b10000101_00101101_10110010_0;
      patterns[34096] = 25'b10000101_00101110_10110011_0;
      patterns[34097] = 25'b10000101_00101111_10110100_0;
      patterns[34098] = 25'b10000101_00110000_10110101_0;
      patterns[34099] = 25'b10000101_00110001_10110110_0;
      patterns[34100] = 25'b10000101_00110010_10110111_0;
      patterns[34101] = 25'b10000101_00110011_10111000_0;
      patterns[34102] = 25'b10000101_00110100_10111001_0;
      patterns[34103] = 25'b10000101_00110101_10111010_0;
      patterns[34104] = 25'b10000101_00110110_10111011_0;
      patterns[34105] = 25'b10000101_00110111_10111100_0;
      patterns[34106] = 25'b10000101_00111000_10111101_0;
      patterns[34107] = 25'b10000101_00111001_10111110_0;
      patterns[34108] = 25'b10000101_00111010_10111111_0;
      patterns[34109] = 25'b10000101_00111011_11000000_0;
      patterns[34110] = 25'b10000101_00111100_11000001_0;
      patterns[34111] = 25'b10000101_00111101_11000010_0;
      patterns[34112] = 25'b10000101_00111110_11000011_0;
      patterns[34113] = 25'b10000101_00111111_11000100_0;
      patterns[34114] = 25'b10000101_01000000_11000101_0;
      patterns[34115] = 25'b10000101_01000001_11000110_0;
      patterns[34116] = 25'b10000101_01000010_11000111_0;
      patterns[34117] = 25'b10000101_01000011_11001000_0;
      patterns[34118] = 25'b10000101_01000100_11001001_0;
      patterns[34119] = 25'b10000101_01000101_11001010_0;
      patterns[34120] = 25'b10000101_01000110_11001011_0;
      patterns[34121] = 25'b10000101_01000111_11001100_0;
      patterns[34122] = 25'b10000101_01001000_11001101_0;
      patterns[34123] = 25'b10000101_01001001_11001110_0;
      patterns[34124] = 25'b10000101_01001010_11001111_0;
      patterns[34125] = 25'b10000101_01001011_11010000_0;
      patterns[34126] = 25'b10000101_01001100_11010001_0;
      patterns[34127] = 25'b10000101_01001101_11010010_0;
      patterns[34128] = 25'b10000101_01001110_11010011_0;
      patterns[34129] = 25'b10000101_01001111_11010100_0;
      patterns[34130] = 25'b10000101_01010000_11010101_0;
      patterns[34131] = 25'b10000101_01010001_11010110_0;
      patterns[34132] = 25'b10000101_01010010_11010111_0;
      patterns[34133] = 25'b10000101_01010011_11011000_0;
      patterns[34134] = 25'b10000101_01010100_11011001_0;
      patterns[34135] = 25'b10000101_01010101_11011010_0;
      patterns[34136] = 25'b10000101_01010110_11011011_0;
      patterns[34137] = 25'b10000101_01010111_11011100_0;
      patterns[34138] = 25'b10000101_01011000_11011101_0;
      patterns[34139] = 25'b10000101_01011001_11011110_0;
      patterns[34140] = 25'b10000101_01011010_11011111_0;
      patterns[34141] = 25'b10000101_01011011_11100000_0;
      patterns[34142] = 25'b10000101_01011100_11100001_0;
      patterns[34143] = 25'b10000101_01011101_11100010_0;
      patterns[34144] = 25'b10000101_01011110_11100011_0;
      patterns[34145] = 25'b10000101_01011111_11100100_0;
      patterns[34146] = 25'b10000101_01100000_11100101_0;
      patterns[34147] = 25'b10000101_01100001_11100110_0;
      patterns[34148] = 25'b10000101_01100010_11100111_0;
      patterns[34149] = 25'b10000101_01100011_11101000_0;
      patterns[34150] = 25'b10000101_01100100_11101001_0;
      patterns[34151] = 25'b10000101_01100101_11101010_0;
      patterns[34152] = 25'b10000101_01100110_11101011_0;
      patterns[34153] = 25'b10000101_01100111_11101100_0;
      patterns[34154] = 25'b10000101_01101000_11101101_0;
      patterns[34155] = 25'b10000101_01101001_11101110_0;
      patterns[34156] = 25'b10000101_01101010_11101111_0;
      patterns[34157] = 25'b10000101_01101011_11110000_0;
      patterns[34158] = 25'b10000101_01101100_11110001_0;
      patterns[34159] = 25'b10000101_01101101_11110010_0;
      patterns[34160] = 25'b10000101_01101110_11110011_0;
      patterns[34161] = 25'b10000101_01101111_11110100_0;
      patterns[34162] = 25'b10000101_01110000_11110101_0;
      patterns[34163] = 25'b10000101_01110001_11110110_0;
      patterns[34164] = 25'b10000101_01110010_11110111_0;
      patterns[34165] = 25'b10000101_01110011_11111000_0;
      patterns[34166] = 25'b10000101_01110100_11111001_0;
      patterns[34167] = 25'b10000101_01110101_11111010_0;
      patterns[34168] = 25'b10000101_01110110_11111011_0;
      patterns[34169] = 25'b10000101_01110111_11111100_0;
      patterns[34170] = 25'b10000101_01111000_11111101_0;
      patterns[34171] = 25'b10000101_01111001_11111110_0;
      patterns[34172] = 25'b10000101_01111010_11111111_0;
      patterns[34173] = 25'b10000101_01111011_00000000_1;
      patterns[34174] = 25'b10000101_01111100_00000001_1;
      patterns[34175] = 25'b10000101_01111101_00000010_1;
      patterns[34176] = 25'b10000101_01111110_00000011_1;
      patterns[34177] = 25'b10000101_01111111_00000100_1;
      patterns[34178] = 25'b10000101_10000000_00000101_1;
      patterns[34179] = 25'b10000101_10000001_00000110_1;
      patterns[34180] = 25'b10000101_10000010_00000111_1;
      patterns[34181] = 25'b10000101_10000011_00001000_1;
      patterns[34182] = 25'b10000101_10000100_00001001_1;
      patterns[34183] = 25'b10000101_10000101_00001010_1;
      patterns[34184] = 25'b10000101_10000110_00001011_1;
      patterns[34185] = 25'b10000101_10000111_00001100_1;
      patterns[34186] = 25'b10000101_10001000_00001101_1;
      patterns[34187] = 25'b10000101_10001001_00001110_1;
      patterns[34188] = 25'b10000101_10001010_00001111_1;
      patterns[34189] = 25'b10000101_10001011_00010000_1;
      patterns[34190] = 25'b10000101_10001100_00010001_1;
      patterns[34191] = 25'b10000101_10001101_00010010_1;
      patterns[34192] = 25'b10000101_10001110_00010011_1;
      patterns[34193] = 25'b10000101_10001111_00010100_1;
      patterns[34194] = 25'b10000101_10010000_00010101_1;
      patterns[34195] = 25'b10000101_10010001_00010110_1;
      patterns[34196] = 25'b10000101_10010010_00010111_1;
      patterns[34197] = 25'b10000101_10010011_00011000_1;
      patterns[34198] = 25'b10000101_10010100_00011001_1;
      patterns[34199] = 25'b10000101_10010101_00011010_1;
      patterns[34200] = 25'b10000101_10010110_00011011_1;
      patterns[34201] = 25'b10000101_10010111_00011100_1;
      patterns[34202] = 25'b10000101_10011000_00011101_1;
      patterns[34203] = 25'b10000101_10011001_00011110_1;
      patterns[34204] = 25'b10000101_10011010_00011111_1;
      patterns[34205] = 25'b10000101_10011011_00100000_1;
      patterns[34206] = 25'b10000101_10011100_00100001_1;
      patterns[34207] = 25'b10000101_10011101_00100010_1;
      patterns[34208] = 25'b10000101_10011110_00100011_1;
      patterns[34209] = 25'b10000101_10011111_00100100_1;
      patterns[34210] = 25'b10000101_10100000_00100101_1;
      patterns[34211] = 25'b10000101_10100001_00100110_1;
      patterns[34212] = 25'b10000101_10100010_00100111_1;
      patterns[34213] = 25'b10000101_10100011_00101000_1;
      patterns[34214] = 25'b10000101_10100100_00101001_1;
      patterns[34215] = 25'b10000101_10100101_00101010_1;
      patterns[34216] = 25'b10000101_10100110_00101011_1;
      patterns[34217] = 25'b10000101_10100111_00101100_1;
      patterns[34218] = 25'b10000101_10101000_00101101_1;
      patterns[34219] = 25'b10000101_10101001_00101110_1;
      patterns[34220] = 25'b10000101_10101010_00101111_1;
      patterns[34221] = 25'b10000101_10101011_00110000_1;
      patterns[34222] = 25'b10000101_10101100_00110001_1;
      patterns[34223] = 25'b10000101_10101101_00110010_1;
      patterns[34224] = 25'b10000101_10101110_00110011_1;
      patterns[34225] = 25'b10000101_10101111_00110100_1;
      patterns[34226] = 25'b10000101_10110000_00110101_1;
      patterns[34227] = 25'b10000101_10110001_00110110_1;
      patterns[34228] = 25'b10000101_10110010_00110111_1;
      patterns[34229] = 25'b10000101_10110011_00111000_1;
      patterns[34230] = 25'b10000101_10110100_00111001_1;
      patterns[34231] = 25'b10000101_10110101_00111010_1;
      patterns[34232] = 25'b10000101_10110110_00111011_1;
      patterns[34233] = 25'b10000101_10110111_00111100_1;
      patterns[34234] = 25'b10000101_10111000_00111101_1;
      patterns[34235] = 25'b10000101_10111001_00111110_1;
      patterns[34236] = 25'b10000101_10111010_00111111_1;
      patterns[34237] = 25'b10000101_10111011_01000000_1;
      patterns[34238] = 25'b10000101_10111100_01000001_1;
      patterns[34239] = 25'b10000101_10111101_01000010_1;
      patterns[34240] = 25'b10000101_10111110_01000011_1;
      patterns[34241] = 25'b10000101_10111111_01000100_1;
      patterns[34242] = 25'b10000101_11000000_01000101_1;
      patterns[34243] = 25'b10000101_11000001_01000110_1;
      patterns[34244] = 25'b10000101_11000010_01000111_1;
      patterns[34245] = 25'b10000101_11000011_01001000_1;
      patterns[34246] = 25'b10000101_11000100_01001001_1;
      patterns[34247] = 25'b10000101_11000101_01001010_1;
      patterns[34248] = 25'b10000101_11000110_01001011_1;
      patterns[34249] = 25'b10000101_11000111_01001100_1;
      patterns[34250] = 25'b10000101_11001000_01001101_1;
      patterns[34251] = 25'b10000101_11001001_01001110_1;
      patterns[34252] = 25'b10000101_11001010_01001111_1;
      patterns[34253] = 25'b10000101_11001011_01010000_1;
      patterns[34254] = 25'b10000101_11001100_01010001_1;
      patterns[34255] = 25'b10000101_11001101_01010010_1;
      patterns[34256] = 25'b10000101_11001110_01010011_1;
      patterns[34257] = 25'b10000101_11001111_01010100_1;
      patterns[34258] = 25'b10000101_11010000_01010101_1;
      patterns[34259] = 25'b10000101_11010001_01010110_1;
      patterns[34260] = 25'b10000101_11010010_01010111_1;
      patterns[34261] = 25'b10000101_11010011_01011000_1;
      patterns[34262] = 25'b10000101_11010100_01011001_1;
      patterns[34263] = 25'b10000101_11010101_01011010_1;
      patterns[34264] = 25'b10000101_11010110_01011011_1;
      patterns[34265] = 25'b10000101_11010111_01011100_1;
      patterns[34266] = 25'b10000101_11011000_01011101_1;
      patterns[34267] = 25'b10000101_11011001_01011110_1;
      patterns[34268] = 25'b10000101_11011010_01011111_1;
      patterns[34269] = 25'b10000101_11011011_01100000_1;
      patterns[34270] = 25'b10000101_11011100_01100001_1;
      patterns[34271] = 25'b10000101_11011101_01100010_1;
      patterns[34272] = 25'b10000101_11011110_01100011_1;
      patterns[34273] = 25'b10000101_11011111_01100100_1;
      patterns[34274] = 25'b10000101_11100000_01100101_1;
      patterns[34275] = 25'b10000101_11100001_01100110_1;
      patterns[34276] = 25'b10000101_11100010_01100111_1;
      patterns[34277] = 25'b10000101_11100011_01101000_1;
      patterns[34278] = 25'b10000101_11100100_01101001_1;
      patterns[34279] = 25'b10000101_11100101_01101010_1;
      patterns[34280] = 25'b10000101_11100110_01101011_1;
      patterns[34281] = 25'b10000101_11100111_01101100_1;
      patterns[34282] = 25'b10000101_11101000_01101101_1;
      patterns[34283] = 25'b10000101_11101001_01101110_1;
      patterns[34284] = 25'b10000101_11101010_01101111_1;
      patterns[34285] = 25'b10000101_11101011_01110000_1;
      patterns[34286] = 25'b10000101_11101100_01110001_1;
      patterns[34287] = 25'b10000101_11101101_01110010_1;
      patterns[34288] = 25'b10000101_11101110_01110011_1;
      patterns[34289] = 25'b10000101_11101111_01110100_1;
      patterns[34290] = 25'b10000101_11110000_01110101_1;
      patterns[34291] = 25'b10000101_11110001_01110110_1;
      patterns[34292] = 25'b10000101_11110010_01110111_1;
      patterns[34293] = 25'b10000101_11110011_01111000_1;
      patterns[34294] = 25'b10000101_11110100_01111001_1;
      patterns[34295] = 25'b10000101_11110101_01111010_1;
      patterns[34296] = 25'b10000101_11110110_01111011_1;
      patterns[34297] = 25'b10000101_11110111_01111100_1;
      patterns[34298] = 25'b10000101_11111000_01111101_1;
      patterns[34299] = 25'b10000101_11111001_01111110_1;
      patterns[34300] = 25'b10000101_11111010_01111111_1;
      patterns[34301] = 25'b10000101_11111011_10000000_1;
      patterns[34302] = 25'b10000101_11111100_10000001_1;
      patterns[34303] = 25'b10000101_11111101_10000010_1;
      patterns[34304] = 25'b10000101_11111110_10000011_1;
      patterns[34305] = 25'b10000101_11111111_10000100_1;
      patterns[34306] = 25'b10000110_00000000_10000110_0;
      patterns[34307] = 25'b10000110_00000001_10000111_0;
      patterns[34308] = 25'b10000110_00000010_10001000_0;
      patterns[34309] = 25'b10000110_00000011_10001001_0;
      patterns[34310] = 25'b10000110_00000100_10001010_0;
      patterns[34311] = 25'b10000110_00000101_10001011_0;
      patterns[34312] = 25'b10000110_00000110_10001100_0;
      patterns[34313] = 25'b10000110_00000111_10001101_0;
      patterns[34314] = 25'b10000110_00001000_10001110_0;
      patterns[34315] = 25'b10000110_00001001_10001111_0;
      patterns[34316] = 25'b10000110_00001010_10010000_0;
      patterns[34317] = 25'b10000110_00001011_10010001_0;
      patterns[34318] = 25'b10000110_00001100_10010010_0;
      patterns[34319] = 25'b10000110_00001101_10010011_0;
      patterns[34320] = 25'b10000110_00001110_10010100_0;
      patterns[34321] = 25'b10000110_00001111_10010101_0;
      patterns[34322] = 25'b10000110_00010000_10010110_0;
      patterns[34323] = 25'b10000110_00010001_10010111_0;
      patterns[34324] = 25'b10000110_00010010_10011000_0;
      patterns[34325] = 25'b10000110_00010011_10011001_0;
      patterns[34326] = 25'b10000110_00010100_10011010_0;
      patterns[34327] = 25'b10000110_00010101_10011011_0;
      patterns[34328] = 25'b10000110_00010110_10011100_0;
      patterns[34329] = 25'b10000110_00010111_10011101_0;
      patterns[34330] = 25'b10000110_00011000_10011110_0;
      patterns[34331] = 25'b10000110_00011001_10011111_0;
      patterns[34332] = 25'b10000110_00011010_10100000_0;
      patterns[34333] = 25'b10000110_00011011_10100001_0;
      patterns[34334] = 25'b10000110_00011100_10100010_0;
      patterns[34335] = 25'b10000110_00011101_10100011_0;
      patterns[34336] = 25'b10000110_00011110_10100100_0;
      patterns[34337] = 25'b10000110_00011111_10100101_0;
      patterns[34338] = 25'b10000110_00100000_10100110_0;
      patterns[34339] = 25'b10000110_00100001_10100111_0;
      patterns[34340] = 25'b10000110_00100010_10101000_0;
      patterns[34341] = 25'b10000110_00100011_10101001_0;
      patterns[34342] = 25'b10000110_00100100_10101010_0;
      patterns[34343] = 25'b10000110_00100101_10101011_0;
      patterns[34344] = 25'b10000110_00100110_10101100_0;
      patterns[34345] = 25'b10000110_00100111_10101101_0;
      patterns[34346] = 25'b10000110_00101000_10101110_0;
      patterns[34347] = 25'b10000110_00101001_10101111_0;
      patterns[34348] = 25'b10000110_00101010_10110000_0;
      patterns[34349] = 25'b10000110_00101011_10110001_0;
      patterns[34350] = 25'b10000110_00101100_10110010_0;
      patterns[34351] = 25'b10000110_00101101_10110011_0;
      patterns[34352] = 25'b10000110_00101110_10110100_0;
      patterns[34353] = 25'b10000110_00101111_10110101_0;
      patterns[34354] = 25'b10000110_00110000_10110110_0;
      patterns[34355] = 25'b10000110_00110001_10110111_0;
      patterns[34356] = 25'b10000110_00110010_10111000_0;
      patterns[34357] = 25'b10000110_00110011_10111001_0;
      patterns[34358] = 25'b10000110_00110100_10111010_0;
      patterns[34359] = 25'b10000110_00110101_10111011_0;
      patterns[34360] = 25'b10000110_00110110_10111100_0;
      patterns[34361] = 25'b10000110_00110111_10111101_0;
      patterns[34362] = 25'b10000110_00111000_10111110_0;
      patterns[34363] = 25'b10000110_00111001_10111111_0;
      patterns[34364] = 25'b10000110_00111010_11000000_0;
      patterns[34365] = 25'b10000110_00111011_11000001_0;
      patterns[34366] = 25'b10000110_00111100_11000010_0;
      patterns[34367] = 25'b10000110_00111101_11000011_0;
      patterns[34368] = 25'b10000110_00111110_11000100_0;
      patterns[34369] = 25'b10000110_00111111_11000101_0;
      patterns[34370] = 25'b10000110_01000000_11000110_0;
      patterns[34371] = 25'b10000110_01000001_11000111_0;
      patterns[34372] = 25'b10000110_01000010_11001000_0;
      patterns[34373] = 25'b10000110_01000011_11001001_0;
      patterns[34374] = 25'b10000110_01000100_11001010_0;
      patterns[34375] = 25'b10000110_01000101_11001011_0;
      patterns[34376] = 25'b10000110_01000110_11001100_0;
      patterns[34377] = 25'b10000110_01000111_11001101_0;
      patterns[34378] = 25'b10000110_01001000_11001110_0;
      patterns[34379] = 25'b10000110_01001001_11001111_0;
      patterns[34380] = 25'b10000110_01001010_11010000_0;
      patterns[34381] = 25'b10000110_01001011_11010001_0;
      patterns[34382] = 25'b10000110_01001100_11010010_0;
      patterns[34383] = 25'b10000110_01001101_11010011_0;
      patterns[34384] = 25'b10000110_01001110_11010100_0;
      patterns[34385] = 25'b10000110_01001111_11010101_0;
      patterns[34386] = 25'b10000110_01010000_11010110_0;
      patterns[34387] = 25'b10000110_01010001_11010111_0;
      patterns[34388] = 25'b10000110_01010010_11011000_0;
      patterns[34389] = 25'b10000110_01010011_11011001_0;
      patterns[34390] = 25'b10000110_01010100_11011010_0;
      patterns[34391] = 25'b10000110_01010101_11011011_0;
      patterns[34392] = 25'b10000110_01010110_11011100_0;
      patterns[34393] = 25'b10000110_01010111_11011101_0;
      patterns[34394] = 25'b10000110_01011000_11011110_0;
      patterns[34395] = 25'b10000110_01011001_11011111_0;
      patterns[34396] = 25'b10000110_01011010_11100000_0;
      patterns[34397] = 25'b10000110_01011011_11100001_0;
      patterns[34398] = 25'b10000110_01011100_11100010_0;
      patterns[34399] = 25'b10000110_01011101_11100011_0;
      patterns[34400] = 25'b10000110_01011110_11100100_0;
      patterns[34401] = 25'b10000110_01011111_11100101_0;
      patterns[34402] = 25'b10000110_01100000_11100110_0;
      patterns[34403] = 25'b10000110_01100001_11100111_0;
      patterns[34404] = 25'b10000110_01100010_11101000_0;
      patterns[34405] = 25'b10000110_01100011_11101001_0;
      patterns[34406] = 25'b10000110_01100100_11101010_0;
      patterns[34407] = 25'b10000110_01100101_11101011_0;
      patterns[34408] = 25'b10000110_01100110_11101100_0;
      patterns[34409] = 25'b10000110_01100111_11101101_0;
      patterns[34410] = 25'b10000110_01101000_11101110_0;
      patterns[34411] = 25'b10000110_01101001_11101111_0;
      patterns[34412] = 25'b10000110_01101010_11110000_0;
      patterns[34413] = 25'b10000110_01101011_11110001_0;
      patterns[34414] = 25'b10000110_01101100_11110010_0;
      patterns[34415] = 25'b10000110_01101101_11110011_0;
      patterns[34416] = 25'b10000110_01101110_11110100_0;
      patterns[34417] = 25'b10000110_01101111_11110101_0;
      patterns[34418] = 25'b10000110_01110000_11110110_0;
      patterns[34419] = 25'b10000110_01110001_11110111_0;
      patterns[34420] = 25'b10000110_01110010_11111000_0;
      patterns[34421] = 25'b10000110_01110011_11111001_0;
      patterns[34422] = 25'b10000110_01110100_11111010_0;
      patterns[34423] = 25'b10000110_01110101_11111011_0;
      patterns[34424] = 25'b10000110_01110110_11111100_0;
      patterns[34425] = 25'b10000110_01110111_11111101_0;
      patterns[34426] = 25'b10000110_01111000_11111110_0;
      patterns[34427] = 25'b10000110_01111001_11111111_0;
      patterns[34428] = 25'b10000110_01111010_00000000_1;
      patterns[34429] = 25'b10000110_01111011_00000001_1;
      patterns[34430] = 25'b10000110_01111100_00000010_1;
      patterns[34431] = 25'b10000110_01111101_00000011_1;
      patterns[34432] = 25'b10000110_01111110_00000100_1;
      patterns[34433] = 25'b10000110_01111111_00000101_1;
      patterns[34434] = 25'b10000110_10000000_00000110_1;
      patterns[34435] = 25'b10000110_10000001_00000111_1;
      patterns[34436] = 25'b10000110_10000010_00001000_1;
      patterns[34437] = 25'b10000110_10000011_00001001_1;
      patterns[34438] = 25'b10000110_10000100_00001010_1;
      patterns[34439] = 25'b10000110_10000101_00001011_1;
      patterns[34440] = 25'b10000110_10000110_00001100_1;
      patterns[34441] = 25'b10000110_10000111_00001101_1;
      patterns[34442] = 25'b10000110_10001000_00001110_1;
      patterns[34443] = 25'b10000110_10001001_00001111_1;
      patterns[34444] = 25'b10000110_10001010_00010000_1;
      patterns[34445] = 25'b10000110_10001011_00010001_1;
      patterns[34446] = 25'b10000110_10001100_00010010_1;
      patterns[34447] = 25'b10000110_10001101_00010011_1;
      patterns[34448] = 25'b10000110_10001110_00010100_1;
      patterns[34449] = 25'b10000110_10001111_00010101_1;
      patterns[34450] = 25'b10000110_10010000_00010110_1;
      patterns[34451] = 25'b10000110_10010001_00010111_1;
      patterns[34452] = 25'b10000110_10010010_00011000_1;
      patterns[34453] = 25'b10000110_10010011_00011001_1;
      patterns[34454] = 25'b10000110_10010100_00011010_1;
      patterns[34455] = 25'b10000110_10010101_00011011_1;
      patterns[34456] = 25'b10000110_10010110_00011100_1;
      patterns[34457] = 25'b10000110_10010111_00011101_1;
      patterns[34458] = 25'b10000110_10011000_00011110_1;
      patterns[34459] = 25'b10000110_10011001_00011111_1;
      patterns[34460] = 25'b10000110_10011010_00100000_1;
      patterns[34461] = 25'b10000110_10011011_00100001_1;
      patterns[34462] = 25'b10000110_10011100_00100010_1;
      patterns[34463] = 25'b10000110_10011101_00100011_1;
      patterns[34464] = 25'b10000110_10011110_00100100_1;
      patterns[34465] = 25'b10000110_10011111_00100101_1;
      patterns[34466] = 25'b10000110_10100000_00100110_1;
      patterns[34467] = 25'b10000110_10100001_00100111_1;
      patterns[34468] = 25'b10000110_10100010_00101000_1;
      patterns[34469] = 25'b10000110_10100011_00101001_1;
      patterns[34470] = 25'b10000110_10100100_00101010_1;
      patterns[34471] = 25'b10000110_10100101_00101011_1;
      patterns[34472] = 25'b10000110_10100110_00101100_1;
      patterns[34473] = 25'b10000110_10100111_00101101_1;
      patterns[34474] = 25'b10000110_10101000_00101110_1;
      patterns[34475] = 25'b10000110_10101001_00101111_1;
      patterns[34476] = 25'b10000110_10101010_00110000_1;
      patterns[34477] = 25'b10000110_10101011_00110001_1;
      patterns[34478] = 25'b10000110_10101100_00110010_1;
      patterns[34479] = 25'b10000110_10101101_00110011_1;
      patterns[34480] = 25'b10000110_10101110_00110100_1;
      patterns[34481] = 25'b10000110_10101111_00110101_1;
      patterns[34482] = 25'b10000110_10110000_00110110_1;
      patterns[34483] = 25'b10000110_10110001_00110111_1;
      patterns[34484] = 25'b10000110_10110010_00111000_1;
      patterns[34485] = 25'b10000110_10110011_00111001_1;
      patterns[34486] = 25'b10000110_10110100_00111010_1;
      patterns[34487] = 25'b10000110_10110101_00111011_1;
      patterns[34488] = 25'b10000110_10110110_00111100_1;
      patterns[34489] = 25'b10000110_10110111_00111101_1;
      patterns[34490] = 25'b10000110_10111000_00111110_1;
      patterns[34491] = 25'b10000110_10111001_00111111_1;
      patterns[34492] = 25'b10000110_10111010_01000000_1;
      patterns[34493] = 25'b10000110_10111011_01000001_1;
      patterns[34494] = 25'b10000110_10111100_01000010_1;
      patterns[34495] = 25'b10000110_10111101_01000011_1;
      patterns[34496] = 25'b10000110_10111110_01000100_1;
      patterns[34497] = 25'b10000110_10111111_01000101_1;
      patterns[34498] = 25'b10000110_11000000_01000110_1;
      patterns[34499] = 25'b10000110_11000001_01000111_1;
      patterns[34500] = 25'b10000110_11000010_01001000_1;
      patterns[34501] = 25'b10000110_11000011_01001001_1;
      patterns[34502] = 25'b10000110_11000100_01001010_1;
      patterns[34503] = 25'b10000110_11000101_01001011_1;
      patterns[34504] = 25'b10000110_11000110_01001100_1;
      patterns[34505] = 25'b10000110_11000111_01001101_1;
      patterns[34506] = 25'b10000110_11001000_01001110_1;
      patterns[34507] = 25'b10000110_11001001_01001111_1;
      patterns[34508] = 25'b10000110_11001010_01010000_1;
      patterns[34509] = 25'b10000110_11001011_01010001_1;
      patterns[34510] = 25'b10000110_11001100_01010010_1;
      patterns[34511] = 25'b10000110_11001101_01010011_1;
      patterns[34512] = 25'b10000110_11001110_01010100_1;
      patterns[34513] = 25'b10000110_11001111_01010101_1;
      patterns[34514] = 25'b10000110_11010000_01010110_1;
      patterns[34515] = 25'b10000110_11010001_01010111_1;
      patterns[34516] = 25'b10000110_11010010_01011000_1;
      patterns[34517] = 25'b10000110_11010011_01011001_1;
      patterns[34518] = 25'b10000110_11010100_01011010_1;
      patterns[34519] = 25'b10000110_11010101_01011011_1;
      patterns[34520] = 25'b10000110_11010110_01011100_1;
      patterns[34521] = 25'b10000110_11010111_01011101_1;
      patterns[34522] = 25'b10000110_11011000_01011110_1;
      patterns[34523] = 25'b10000110_11011001_01011111_1;
      patterns[34524] = 25'b10000110_11011010_01100000_1;
      patterns[34525] = 25'b10000110_11011011_01100001_1;
      patterns[34526] = 25'b10000110_11011100_01100010_1;
      patterns[34527] = 25'b10000110_11011101_01100011_1;
      patterns[34528] = 25'b10000110_11011110_01100100_1;
      patterns[34529] = 25'b10000110_11011111_01100101_1;
      patterns[34530] = 25'b10000110_11100000_01100110_1;
      patterns[34531] = 25'b10000110_11100001_01100111_1;
      patterns[34532] = 25'b10000110_11100010_01101000_1;
      patterns[34533] = 25'b10000110_11100011_01101001_1;
      patterns[34534] = 25'b10000110_11100100_01101010_1;
      patterns[34535] = 25'b10000110_11100101_01101011_1;
      patterns[34536] = 25'b10000110_11100110_01101100_1;
      patterns[34537] = 25'b10000110_11100111_01101101_1;
      patterns[34538] = 25'b10000110_11101000_01101110_1;
      patterns[34539] = 25'b10000110_11101001_01101111_1;
      patterns[34540] = 25'b10000110_11101010_01110000_1;
      patterns[34541] = 25'b10000110_11101011_01110001_1;
      patterns[34542] = 25'b10000110_11101100_01110010_1;
      patterns[34543] = 25'b10000110_11101101_01110011_1;
      patterns[34544] = 25'b10000110_11101110_01110100_1;
      patterns[34545] = 25'b10000110_11101111_01110101_1;
      patterns[34546] = 25'b10000110_11110000_01110110_1;
      patterns[34547] = 25'b10000110_11110001_01110111_1;
      patterns[34548] = 25'b10000110_11110010_01111000_1;
      patterns[34549] = 25'b10000110_11110011_01111001_1;
      patterns[34550] = 25'b10000110_11110100_01111010_1;
      patterns[34551] = 25'b10000110_11110101_01111011_1;
      patterns[34552] = 25'b10000110_11110110_01111100_1;
      patterns[34553] = 25'b10000110_11110111_01111101_1;
      patterns[34554] = 25'b10000110_11111000_01111110_1;
      patterns[34555] = 25'b10000110_11111001_01111111_1;
      patterns[34556] = 25'b10000110_11111010_10000000_1;
      patterns[34557] = 25'b10000110_11111011_10000001_1;
      patterns[34558] = 25'b10000110_11111100_10000010_1;
      patterns[34559] = 25'b10000110_11111101_10000011_1;
      patterns[34560] = 25'b10000110_11111110_10000100_1;
      patterns[34561] = 25'b10000110_11111111_10000101_1;
      patterns[34562] = 25'b10000111_00000000_10000111_0;
      patterns[34563] = 25'b10000111_00000001_10001000_0;
      patterns[34564] = 25'b10000111_00000010_10001001_0;
      patterns[34565] = 25'b10000111_00000011_10001010_0;
      patterns[34566] = 25'b10000111_00000100_10001011_0;
      patterns[34567] = 25'b10000111_00000101_10001100_0;
      patterns[34568] = 25'b10000111_00000110_10001101_0;
      patterns[34569] = 25'b10000111_00000111_10001110_0;
      patterns[34570] = 25'b10000111_00001000_10001111_0;
      patterns[34571] = 25'b10000111_00001001_10010000_0;
      patterns[34572] = 25'b10000111_00001010_10010001_0;
      patterns[34573] = 25'b10000111_00001011_10010010_0;
      patterns[34574] = 25'b10000111_00001100_10010011_0;
      patterns[34575] = 25'b10000111_00001101_10010100_0;
      patterns[34576] = 25'b10000111_00001110_10010101_0;
      patterns[34577] = 25'b10000111_00001111_10010110_0;
      patterns[34578] = 25'b10000111_00010000_10010111_0;
      patterns[34579] = 25'b10000111_00010001_10011000_0;
      patterns[34580] = 25'b10000111_00010010_10011001_0;
      patterns[34581] = 25'b10000111_00010011_10011010_0;
      patterns[34582] = 25'b10000111_00010100_10011011_0;
      patterns[34583] = 25'b10000111_00010101_10011100_0;
      patterns[34584] = 25'b10000111_00010110_10011101_0;
      patterns[34585] = 25'b10000111_00010111_10011110_0;
      patterns[34586] = 25'b10000111_00011000_10011111_0;
      patterns[34587] = 25'b10000111_00011001_10100000_0;
      patterns[34588] = 25'b10000111_00011010_10100001_0;
      patterns[34589] = 25'b10000111_00011011_10100010_0;
      patterns[34590] = 25'b10000111_00011100_10100011_0;
      patterns[34591] = 25'b10000111_00011101_10100100_0;
      patterns[34592] = 25'b10000111_00011110_10100101_0;
      patterns[34593] = 25'b10000111_00011111_10100110_0;
      patterns[34594] = 25'b10000111_00100000_10100111_0;
      patterns[34595] = 25'b10000111_00100001_10101000_0;
      patterns[34596] = 25'b10000111_00100010_10101001_0;
      patterns[34597] = 25'b10000111_00100011_10101010_0;
      patterns[34598] = 25'b10000111_00100100_10101011_0;
      patterns[34599] = 25'b10000111_00100101_10101100_0;
      patterns[34600] = 25'b10000111_00100110_10101101_0;
      patterns[34601] = 25'b10000111_00100111_10101110_0;
      patterns[34602] = 25'b10000111_00101000_10101111_0;
      patterns[34603] = 25'b10000111_00101001_10110000_0;
      patterns[34604] = 25'b10000111_00101010_10110001_0;
      patterns[34605] = 25'b10000111_00101011_10110010_0;
      patterns[34606] = 25'b10000111_00101100_10110011_0;
      patterns[34607] = 25'b10000111_00101101_10110100_0;
      patterns[34608] = 25'b10000111_00101110_10110101_0;
      patterns[34609] = 25'b10000111_00101111_10110110_0;
      patterns[34610] = 25'b10000111_00110000_10110111_0;
      patterns[34611] = 25'b10000111_00110001_10111000_0;
      patterns[34612] = 25'b10000111_00110010_10111001_0;
      patterns[34613] = 25'b10000111_00110011_10111010_0;
      patterns[34614] = 25'b10000111_00110100_10111011_0;
      patterns[34615] = 25'b10000111_00110101_10111100_0;
      patterns[34616] = 25'b10000111_00110110_10111101_0;
      patterns[34617] = 25'b10000111_00110111_10111110_0;
      patterns[34618] = 25'b10000111_00111000_10111111_0;
      patterns[34619] = 25'b10000111_00111001_11000000_0;
      patterns[34620] = 25'b10000111_00111010_11000001_0;
      patterns[34621] = 25'b10000111_00111011_11000010_0;
      patterns[34622] = 25'b10000111_00111100_11000011_0;
      patterns[34623] = 25'b10000111_00111101_11000100_0;
      patterns[34624] = 25'b10000111_00111110_11000101_0;
      patterns[34625] = 25'b10000111_00111111_11000110_0;
      patterns[34626] = 25'b10000111_01000000_11000111_0;
      patterns[34627] = 25'b10000111_01000001_11001000_0;
      patterns[34628] = 25'b10000111_01000010_11001001_0;
      patterns[34629] = 25'b10000111_01000011_11001010_0;
      patterns[34630] = 25'b10000111_01000100_11001011_0;
      patterns[34631] = 25'b10000111_01000101_11001100_0;
      patterns[34632] = 25'b10000111_01000110_11001101_0;
      patterns[34633] = 25'b10000111_01000111_11001110_0;
      patterns[34634] = 25'b10000111_01001000_11001111_0;
      patterns[34635] = 25'b10000111_01001001_11010000_0;
      patterns[34636] = 25'b10000111_01001010_11010001_0;
      patterns[34637] = 25'b10000111_01001011_11010010_0;
      patterns[34638] = 25'b10000111_01001100_11010011_0;
      patterns[34639] = 25'b10000111_01001101_11010100_0;
      patterns[34640] = 25'b10000111_01001110_11010101_0;
      patterns[34641] = 25'b10000111_01001111_11010110_0;
      patterns[34642] = 25'b10000111_01010000_11010111_0;
      patterns[34643] = 25'b10000111_01010001_11011000_0;
      patterns[34644] = 25'b10000111_01010010_11011001_0;
      patterns[34645] = 25'b10000111_01010011_11011010_0;
      patterns[34646] = 25'b10000111_01010100_11011011_0;
      patterns[34647] = 25'b10000111_01010101_11011100_0;
      patterns[34648] = 25'b10000111_01010110_11011101_0;
      patterns[34649] = 25'b10000111_01010111_11011110_0;
      patterns[34650] = 25'b10000111_01011000_11011111_0;
      patterns[34651] = 25'b10000111_01011001_11100000_0;
      patterns[34652] = 25'b10000111_01011010_11100001_0;
      patterns[34653] = 25'b10000111_01011011_11100010_0;
      patterns[34654] = 25'b10000111_01011100_11100011_0;
      patterns[34655] = 25'b10000111_01011101_11100100_0;
      patterns[34656] = 25'b10000111_01011110_11100101_0;
      patterns[34657] = 25'b10000111_01011111_11100110_0;
      patterns[34658] = 25'b10000111_01100000_11100111_0;
      patterns[34659] = 25'b10000111_01100001_11101000_0;
      patterns[34660] = 25'b10000111_01100010_11101001_0;
      patterns[34661] = 25'b10000111_01100011_11101010_0;
      patterns[34662] = 25'b10000111_01100100_11101011_0;
      patterns[34663] = 25'b10000111_01100101_11101100_0;
      patterns[34664] = 25'b10000111_01100110_11101101_0;
      patterns[34665] = 25'b10000111_01100111_11101110_0;
      patterns[34666] = 25'b10000111_01101000_11101111_0;
      patterns[34667] = 25'b10000111_01101001_11110000_0;
      patterns[34668] = 25'b10000111_01101010_11110001_0;
      patterns[34669] = 25'b10000111_01101011_11110010_0;
      patterns[34670] = 25'b10000111_01101100_11110011_0;
      patterns[34671] = 25'b10000111_01101101_11110100_0;
      patterns[34672] = 25'b10000111_01101110_11110101_0;
      patterns[34673] = 25'b10000111_01101111_11110110_0;
      patterns[34674] = 25'b10000111_01110000_11110111_0;
      patterns[34675] = 25'b10000111_01110001_11111000_0;
      patterns[34676] = 25'b10000111_01110010_11111001_0;
      patterns[34677] = 25'b10000111_01110011_11111010_0;
      patterns[34678] = 25'b10000111_01110100_11111011_0;
      patterns[34679] = 25'b10000111_01110101_11111100_0;
      patterns[34680] = 25'b10000111_01110110_11111101_0;
      patterns[34681] = 25'b10000111_01110111_11111110_0;
      patterns[34682] = 25'b10000111_01111000_11111111_0;
      patterns[34683] = 25'b10000111_01111001_00000000_1;
      patterns[34684] = 25'b10000111_01111010_00000001_1;
      patterns[34685] = 25'b10000111_01111011_00000010_1;
      patterns[34686] = 25'b10000111_01111100_00000011_1;
      patterns[34687] = 25'b10000111_01111101_00000100_1;
      patterns[34688] = 25'b10000111_01111110_00000101_1;
      patterns[34689] = 25'b10000111_01111111_00000110_1;
      patterns[34690] = 25'b10000111_10000000_00000111_1;
      patterns[34691] = 25'b10000111_10000001_00001000_1;
      patterns[34692] = 25'b10000111_10000010_00001001_1;
      patterns[34693] = 25'b10000111_10000011_00001010_1;
      patterns[34694] = 25'b10000111_10000100_00001011_1;
      patterns[34695] = 25'b10000111_10000101_00001100_1;
      patterns[34696] = 25'b10000111_10000110_00001101_1;
      patterns[34697] = 25'b10000111_10000111_00001110_1;
      patterns[34698] = 25'b10000111_10001000_00001111_1;
      patterns[34699] = 25'b10000111_10001001_00010000_1;
      patterns[34700] = 25'b10000111_10001010_00010001_1;
      patterns[34701] = 25'b10000111_10001011_00010010_1;
      patterns[34702] = 25'b10000111_10001100_00010011_1;
      patterns[34703] = 25'b10000111_10001101_00010100_1;
      patterns[34704] = 25'b10000111_10001110_00010101_1;
      patterns[34705] = 25'b10000111_10001111_00010110_1;
      patterns[34706] = 25'b10000111_10010000_00010111_1;
      patterns[34707] = 25'b10000111_10010001_00011000_1;
      patterns[34708] = 25'b10000111_10010010_00011001_1;
      patterns[34709] = 25'b10000111_10010011_00011010_1;
      patterns[34710] = 25'b10000111_10010100_00011011_1;
      patterns[34711] = 25'b10000111_10010101_00011100_1;
      patterns[34712] = 25'b10000111_10010110_00011101_1;
      patterns[34713] = 25'b10000111_10010111_00011110_1;
      patterns[34714] = 25'b10000111_10011000_00011111_1;
      patterns[34715] = 25'b10000111_10011001_00100000_1;
      patterns[34716] = 25'b10000111_10011010_00100001_1;
      patterns[34717] = 25'b10000111_10011011_00100010_1;
      patterns[34718] = 25'b10000111_10011100_00100011_1;
      patterns[34719] = 25'b10000111_10011101_00100100_1;
      patterns[34720] = 25'b10000111_10011110_00100101_1;
      patterns[34721] = 25'b10000111_10011111_00100110_1;
      patterns[34722] = 25'b10000111_10100000_00100111_1;
      patterns[34723] = 25'b10000111_10100001_00101000_1;
      patterns[34724] = 25'b10000111_10100010_00101001_1;
      patterns[34725] = 25'b10000111_10100011_00101010_1;
      patterns[34726] = 25'b10000111_10100100_00101011_1;
      patterns[34727] = 25'b10000111_10100101_00101100_1;
      patterns[34728] = 25'b10000111_10100110_00101101_1;
      patterns[34729] = 25'b10000111_10100111_00101110_1;
      patterns[34730] = 25'b10000111_10101000_00101111_1;
      patterns[34731] = 25'b10000111_10101001_00110000_1;
      patterns[34732] = 25'b10000111_10101010_00110001_1;
      patterns[34733] = 25'b10000111_10101011_00110010_1;
      patterns[34734] = 25'b10000111_10101100_00110011_1;
      patterns[34735] = 25'b10000111_10101101_00110100_1;
      patterns[34736] = 25'b10000111_10101110_00110101_1;
      patterns[34737] = 25'b10000111_10101111_00110110_1;
      patterns[34738] = 25'b10000111_10110000_00110111_1;
      patterns[34739] = 25'b10000111_10110001_00111000_1;
      patterns[34740] = 25'b10000111_10110010_00111001_1;
      patterns[34741] = 25'b10000111_10110011_00111010_1;
      patterns[34742] = 25'b10000111_10110100_00111011_1;
      patterns[34743] = 25'b10000111_10110101_00111100_1;
      patterns[34744] = 25'b10000111_10110110_00111101_1;
      patterns[34745] = 25'b10000111_10110111_00111110_1;
      patterns[34746] = 25'b10000111_10111000_00111111_1;
      patterns[34747] = 25'b10000111_10111001_01000000_1;
      patterns[34748] = 25'b10000111_10111010_01000001_1;
      patterns[34749] = 25'b10000111_10111011_01000010_1;
      patterns[34750] = 25'b10000111_10111100_01000011_1;
      patterns[34751] = 25'b10000111_10111101_01000100_1;
      patterns[34752] = 25'b10000111_10111110_01000101_1;
      patterns[34753] = 25'b10000111_10111111_01000110_1;
      patterns[34754] = 25'b10000111_11000000_01000111_1;
      patterns[34755] = 25'b10000111_11000001_01001000_1;
      patterns[34756] = 25'b10000111_11000010_01001001_1;
      patterns[34757] = 25'b10000111_11000011_01001010_1;
      patterns[34758] = 25'b10000111_11000100_01001011_1;
      patterns[34759] = 25'b10000111_11000101_01001100_1;
      patterns[34760] = 25'b10000111_11000110_01001101_1;
      patterns[34761] = 25'b10000111_11000111_01001110_1;
      patterns[34762] = 25'b10000111_11001000_01001111_1;
      patterns[34763] = 25'b10000111_11001001_01010000_1;
      patterns[34764] = 25'b10000111_11001010_01010001_1;
      patterns[34765] = 25'b10000111_11001011_01010010_1;
      patterns[34766] = 25'b10000111_11001100_01010011_1;
      patterns[34767] = 25'b10000111_11001101_01010100_1;
      patterns[34768] = 25'b10000111_11001110_01010101_1;
      patterns[34769] = 25'b10000111_11001111_01010110_1;
      patterns[34770] = 25'b10000111_11010000_01010111_1;
      patterns[34771] = 25'b10000111_11010001_01011000_1;
      patterns[34772] = 25'b10000111_11010010_01011001_1;
      patterns[34773] = 25'b10000111_11010011_01011010_1;
      patterns[34774] = 25'b10000111_11010100_01011011_1;
      patterns[34775] = 25'b10000111_11010101_01011100_1;
      patterns[34776] = 25'b10000111_11010110_01011101_1;
      patterns[34777] = 25'b10000111_11010111_01011110_1;
      patterns[34778] = 25'b10000111_11011000_01011111_1;
      patterns[34779] = 25'b10000111_11011001_01100000_1;
      patterns[34780] = 25'b10000111_11011010_01100001_1;
      patterns[34781] = 25'b10000111_11011011_01100010_1;
      patterns[34782] = 25'b10000111_11011100_01100011_1;
      patterns[34783] = 25'b10000111_11011101_01100100_1;
      patterns[34784] = 25'b10000111_11011110_01100101_1;
      patterns[34785] = 25'b10000111_11011111_01100110_1;
      patterns[34786] = 25'b10000111_11100000_01100111_1;
      patterns[34787] = 25'b10000111_11100001_01101000_1;
      patterns[34788] = 25'b10000111_11100010_01101001_1;
      patterns[34789] = 25'b10000111_11100011_01101010_1;
      patterns[34790] = 25'b10000111_11100100_01101011_1;
      patterns[34791] = 25'b10000111_11100101_01101100_1;
      patterns[34792] = 25'b10000111_11100110_01101101_1;
      patterns[34793] = 25'b10000111_11100111_01101110_1;
      patterns[34794] = 25'b10000111_11101000_01101111_1;
      patterns[34795] = 25'b10000111_11101001_01110000_1;
      patterns[34796] = 25'b10000111_11101010_01110001_1;
      patterns[34797] = 25'b10000111_11101011_01110010_1;
      patterns[34798] = 25'b10000111_11101100_01110011_1;
      patterns[34799] = 25'b10000111_11101101_01110100_1;
      patterns[34800] = 25'b10000111_11101110_01110101_1;
      patterns[34801] = 25'b10000111_11101111_01110110_1;
      patterns[34802] = 25'b10000111_11110000_01110111_1;
      patterns[34803] = 25'b10000111_11110001_01111000_1;
      patterns[34804] = 25'b10000111_11110010_01111001_1;
      patterns[34805] = 25'b10000111_11110011_01111010_1;
      patterns[34806] = 25'b10000111_11110100_01111011_1;
      patterns[34807] = 25'b10000111_11110101_01111100_1;
      patterns[34808] = 25'b10000111_11110110_01111101_1;
      patterns[34809] = 25'b10000111_11110111_01111110_1;
      patterns[34810] = 25'b10000111_11111000_01111111_1;
      patterns[34811] = 25'b10000111_11111001_10000000_1;
      patterns[34812] = 25'b10000111_11111010_10000001_1;
      patterns[34813] = 25'b10000111_11111011_10000010_1;
      patterns[34814] = 25'b10000111_11111100_10000011_1;
      patterns[34815] = 25'b10000111_11111101_10000100_1;
      patterns[34816] = 25'b10000111_11111110_10000101_1;
      patterns[34817] = 25'b10000111_11111111_10000110_1;
      patterns[34818] = 25'b10001000_00000000_10001000_0;
      patterns[34819] = 25'b10001000_00000001_10001001_0;
      patterns[34820] = 25'b10001000_00000010_10001010_0;
      patterns[34821] = 25'b10001000_00000011_10001011_0;
      patterns[34822] = 25'b10001000_00000100_10001100_0;
      patterns[34823] = 25'b10001000_00000101_10001101_0;
      patterns[34824] = 25'b10001000_00000110_10001110_0;
      patterns[34825] = 25'b10001000_00000111_10001111_0;
      patterns[34826] = 25'b10001000_00001000_10010000_0;
      patterns[34827] = 25'b10001000_00001001_10010001_0;
      patterns[34828] = 25'b10001000_00001010_10010010_0;
      patterns[34829] = 25'b10001000_00001011_10010011_0;
      patterns[34830] = 25'b10001000_00001100_10010100_0;
      patterns[34831] = 25'b10001000_00001101_10010101_0;
      patterns[34832] = 25'b10001000_00001110_10010110_0;
      patterns[34833] = 25'b10001000_00001111_10010111_0;
      patterns[34834] = 25'b10001000_00010000_10011000_0;
      patterns[34835] = 25'b10001000_00010001_10011001_0;
      patterns[34836] = 25'b10001000_00010010_10011010_0;
      patterns[34837] = 25'b10001000_00010011_10011011_0;
      patterns[34838] = 25'b10001000_00010100_10011100_0;
      patterns[34839] = 25'b10001000_00010101_10011101_0;
      patterns[34840] = 25'b10001000_00010110_10011110_0;
      patterns[34841] = 25'b10001000_00010111_10011111_0;
      patterns[34842] = 25'b10001000_00011000_10100000_0;
      patterns[34843] = 25'b10001000_00011001_10100001_0;
      patterns[34844] = 25'b10001000_00011010_10100010_0;
      patterns[34845] = 25'b10001000_00011011_10100011_0;
      patterns[34846] = 25'b10001000_00011100_10100100_0;
      patterns[34847] = 25'b10001000_00011101_10100101_0;
      patterns[34848] = 25'b10001000_00011110_10100110_0;
      patterns[34849] = 25'b10001000_00011111_10100111_0;
      patterns[34850] = 25'b10001000_00100000_10101000_0;
      patterns[34851] = 25'b10001000_00100001_10101001_0;
      patterns[34852] = 25'b10001000_00100010_10101010_0;
      patterns[34853] = 25'b10001000_00100011_10101011_0;
      patterns[34854] = 25'b10001000_00100100_10101100_0;
      patterns[34855] = 25'b10001000_00100101_10101101_0;
      patterns[34856] = 25'b10001000_00100110_10101110_0;
      patterns[34857] = 25'b10001000_00100111_10101111_0;
      patterns[34858] = 25'b10001000_00101000_10110000_0;
      patterns[34859] = 25'b10001000_00101001_10110001_0;
      patterns[34860] = 25'b10001000_00101010_10110010_0;
      patterns[34861] = 25'b10001000_00101011_10110011_0;
      patterns[34862] = 25'b10001000_00101100_10110100_0;
      patterns[34863] = 25'b10001000_00101101_10110101_0;
      patterns[34864] = 25'b10001000_00101110_10110110_0;
      patterns[34865] = 25'b10001000_00101111_10110111_0;
      patterns[34866] = 25'b10001000_00110000_10111000_0;
      patterns[34867] = 25'b10001000_00110001_10111001_0;
      patterns[34868] = 25'b10001000_00110010_10111010_0;
      patterns[34869] = 25'b10001000_00110011_10111011_0;
      patterns[34870] = 25'b10001000_00110100_10111100_0;
      patterns[34871] = 25'b10001000_00110101_10111101_0;
      patterns[34872] = 25'b10001000_00110110_10111110_0;
      patterns[34873] = 25'b10001000_00110111_10111111_0;
      patterns[34874] = 25'b10001000_00111000_11000000_0;
      patterns[34875] = 25'b10001000_00111001_11000001_0;
      patterns[34876] = 25'b10001000_00111010_11000010_0;
      patterns[34877] = 25'b10001000_00111011_11000011_0;
      patterns[34878] = 25'b10001000_00111100_11000100_0;
      patterns[34879] = 25'b10001000_00111101_11000101_0;
      patterns[34880] = 25'b10001000_00111110_11000110_0;
      patterns[34881] = 25'b10001000_00111111_11000111_0;
      patterns[34882] = 25'b10001000_01000000_11001000_0;
      patterns[34883] = 25'b10001000_01000001_11001001_0;
      patterns[34884] = 25'b10001000_01000010_11001010_0;
      patterns[34885] = 25'b10001000_01000011_11001011_0;
      patterns[34886] = 25'b10001000_01000100_11001100_0;
      patterns[34887] = 25'b10001000_01000101_11001101_0;
      patterns[34888] = 25'b10001000_01000110_11001110_0;
      patterns[34889] = 25'b10001000_01000111_11001111_0;
      patterns[34890] = 25'b10001000_01001000_11010000_0;
      patterns[34891] = 25'b10001000_01001001_11010001_0;
      patterns[34892] = 25'b10001000_01001010_11010010_0;
      patterns[34893] = 25'b10001000_01001011_11010011_0;
      patterns[34894] = 25'b10001000_01001100_11010100_0;
      patterns[34895] = 25'b10001000_01001101_11010101_0;
      patterns[34896] = 25'b10001000_01001110_11010110_0;
      patterns[34897] = 25'b10001000_01001111_11010111_0;
      patterns[34898] = 25'b10001000_01010000_11011000_0;
      patterns[34899] = 25'b10001000_01010001_11011001_0;
      patterns[34900] = 25'b10001000_01010010_11011010_0;
      patterns[34901] = 25'b10001000_01010011_11011011_0;
      patterns[34902] = 25'b10001000_01010100_11011100_0;
      patterns[34903] = 25'b10001000_01010101_11011101_0;
      patterns[34904] = 25'b10001000_01010110_11011110_0;
      patterns[34905] = 25'b10001000_01010111_11011111_0;
      patterns[34906] = 25'b10001000_01011000_11100000_0;
      patterns[34907] = 25'b10001000_01011001_11100001_0;
      patterns[34908] = 25'b10001000_01011010_11100010_0;
      patterns[34909] = 25'b10001000_01011011_11100011_0;
      patterns[34910] = 25'b10001000_01011100_11100100_0;
      patterns[34911] = 25'b10001000_01011101_11100101_0;
      patterns[34912] = 25'b10001000_01011110_11100110_0;
      patterns[34913] = 25'b10001000_01011111_11100111_0;
      patterns[34914] = 25'b10001000_01100000_11101000_0;
      patterns[34915] = 25'b10001000_01100001_11101001_0;
      patterns[34916] = 25'b10001000_01100010_11101010_0;
      patterns[34917] = 25'b10001000_01100011_11101011_0;
      patterns[34918] = 25'b10001000_01100100_11101100_0;
      patterns[34919] = 25'b10001000_01100101_11101101_0;
      patterns[34920] = 25'b10001000_01100110_11101110_0;
      patterns[34921] = 25'b10001000_01100111_11101111_0;
      patterns[34922] = 25'b10001000_01101000_11110000_0;
      patterns[34923] = 25'b10001000_01101001_11110001_0;
      patterns[34924] = 25'b10001000_01101010_11110010_0;
      patterns[34925] = 25'b10001000_01101011_11110011_0;
      patterns[34926] = 25'b10001000_01101100_11110100_0;
      patterns[34927] = 25'b10001000_01101101_11110101_0;
      patterns[34928] = 25'b10001000_01101110_11110110_0;
      patterns[34929] = 25'b10001000_01101111_11110111_0;
      patterns[34930] = 25'b10001000_01110000_11111000_0;
      patterns[34931] = 25'b10001000_01110001_11111001_0;
      patterns[34932] = 25'b10001000_01110010_11111010_0;
      patterns[34933] = 25'b10001000_01110011_11111011_0;
      patterns[34934] = 25'b10001000_01110100_11111100_0;
      patterns[34935] = 25'b10001000_01110101_11111101_0;
      patterns[34936] = 25'b10001000_01110110_11111110_0;
      patterns[34937] = 25'b10001000_01110111_11111111_0;
      patterns[34938] = 25'b10001000_01111000_00000000_1;
      patterns[34939] = 25'b10001000_01111001_00000001_1;
      patterns[34940] = 25'b10001000_01111010_00000010_1;
      patterns[34941] = 25'b10001000_01111011_00000011_1;
      patterns[34942] = 25'b10001000_01111100_00000100_1;
      patterns[34943] = 25'b10001000_01111101_00000101_1;
      patterns[34944] = 25'b10001000_01111110_00000110_1;
      patterns[34945] = 25'b10001000_01111111_00000111_1;
      patterns[34946] = 25'b10001000_10000000_00001000_1;
      patterns[34947] = 25'b10001000_10000001_00001001_1;
      patterns[34948] = 25'b10001000_10000010_00001010_1;
      patterns[34949] = 25'b10001000_10000011_00001011_1;
      patterns[34950] = 25'b10001000_10000100_00001100_1;
      patterns[34951] = 25'b10001000_10000101_00001101_1;
      patterns[34952] = 25'b10001000_10000110_00001110_1;
      patterns[34953] = 25'b10001000_10000111_00001111_1;
      patterns[34954] = 25'b10001000_10001000_00010000_1;
      patterns[34955] = 25'b10001000_10001001_00010001_1;
      patterns[34956] = 25'b10001000_10001010_00010010_1;
      patterns[34957] = 25'b10001000_10001011_00010011_1;
      patterns[34958] = 25'b10001000_10001100_00010100_1;
      patterns[34959] = 25'b10001000_10001101_00010101_1;
      patterns[34960] = 25'b10001000_10001110_00010110_1;
      patterns[34961] = 25'b10001000_10001111_00010111_1;
      patterns[34962] = 25'b10001000_10010000_00011000_1;
      patterns[34963] = 25'b10001000_10010001_00011001_1;
      patterns[34964] = 25'b10001000_10010010_00011010_1;
      patterns[34965] = 25'b10001000_10010011_00011011_1;
      patterns[34966] = 25'b10001000_10010100_00011100_1;
      patterns[34967] = 25'b10001000_10010101_00011101_1;
      patterns[34968] = 25'b10001000_10010110_00011110_1;
      patterns[34969] = 25'b10001000_10010111_00011111_1;
      patterns[34970] = 25'b10001000_10011000_00100000_1;
      patterns[34971] = 25'b10001000_10011001_00100001_1;
      patterns[34972] = 25'b10001000_10011010_00100010_1;
      patterns[34973] = 25'b10001000_10011011_00100011_1;
      patterns[34974] = 25'b10001000_10011100_00100100_1;
      patterns[34975] = 25'b10001000_10011101_00100101_1;
      patterns[34976] = 25'b10001000_10011110_00100110_1;
      patterns[34977] = 25'b10001000_10011111_00100111_1;
      patterns[34978] = 25'b10001000_10100000_00101000_1;
      patterns[34979] = 25'b10001000_10100001_00101001_1;
      patterns[34980] = 25'b10001000_10100010_00101010_1;
      patterns[34981] = 25'b10001000_10100011_00101011_1;
      patterns[34982] = 25'b10001000_10100100_00101100_1;
      patterns[34983] = 25'b10001000_10100101_00101101_1;
      patterns[34984] = 25'b10001000_10100110_00101110_1;
      patterns[34985] = 25'b10001000_10100111_00101111_1;
      patterns[34986] = 25'b10001000_10101000_00110000_1;
      patterns[34987] = 25'b10001000_10101001_00110001_1;
      patterns[34988] = 25'b10001000_10101010_00110010_1;
      patterns[34989] = 25'b10001000_10101011_00110011_1;
      patterns[34990] = 25'b10001000_10101100_00110100_1;
      patterns[34991] = 25'b10001000_10101101_00110101_1;
      patterns[34992] = 25'b10001000_10101110_00110110_1;
      patterns[34993] = 25'b10001000_10101111_00110111_1;
      patterns[34994] = 25'b10001000_10110000_00111000_1;
      patterns[34995] = 25'b10001000_10110001_00111001_1;
      patterns[34996] = 25'b10001000_10110010_00111010_1;
      patterns[34997] = 25'b10001000_10110011_00111011_1;
      patterns[34998] = 25'b10001000_10110100_00111100_1;
      patterns[34999] = 25'b10001000_10110101_00111101_1;
      patterns[35000] = 25'b10001000_10110110_00111110_1;
      patterns[35001] = 25'b10001000_10110111_00111111_1;
      patterns[35002] = 25'b10001000_10111000_01000000_1;
      patterns[35003] = 25'b10001000_10111001_01000001_1;
      patterns[35004] = 25'b10001000_10111010_01000010_1;
      patterns[35005] = 25'b10001000_10111011_01000011_1;
      patterns[35006] = 25'b10001000_10111100_01000100_1;
      patterns[35007] = 25'b10001000_10111101_01000101_1;
      patterns[35008] = 25'b10001000_10111110_01000110_1;
      patterns[35009] = 25'b10001000_10111111_01000111_1;
      patterns[35010] = 25'b10001000_11000000_01001000_1;
      patterns[35011] = 25'b10001000_11000001_01001001_1;
      patterns[35012] = 25'b10001000_11000010_01001010_1;
      patterns[35013] = 25'b10001000_11000011_01001011_1;
      patterns[35014] = 25'b10001000_11000100_01001100_1;
      patterns[35015] = 25'b10001000_11000101_01001101_1;
      patterns[35016] = 25'b10001000_11000110_01001110_1;
      patterns[35017] = 25'b10001000_11000111_01001111_1;
      patterns[35018] = 25'b10001000_11001000_01010000_1;
      patterns[35019] = 25'b10001000_11001001_01010001_1;
      patterns[35020] = 25'b10001000_11001010_01010010_1;
      patterns[35021] = 25'b10001000_11001011_01010011_1;
      patterns[35022] = 25'b10001000_11001100_01010100_1;
      patterns[35023] = 25'b10001000_11001101_01010101_1;
      patterns[35024] = 25'b10001000_11001110_01010110_1;
      patterns[35025] = 25'b10001000_11001111_01010111_1;
      patterns[35026] = 25'b10001000_11010000_01011000_1;
      patterns[35027] = 25'b10001000_11010001_01011001_1;
      patterns[35028] = 25'b10001000_11010010_01011010_1;
      patterns[35029] = 25'b10001000_11010011_01011011_1;
      patterns[35030] = 25'b10001000_11010100_01011100_1;
      patterns[35031] = 25'b10001000_11010101_01011101_1;
      patterns[35032] = 25'b10001000_11010110_01011110_1;
      patterns[35033] = 25'b10001000_11010111_01011111_1;
      patterns[35034] = 25'b10001000_11011000_01100000_1;
      patterns[35035] = 25'b10001000_11011001_01100001_1;
      patterns[35036] = 25'b10001000_11011010_01100010_1;
      patterns[35037] = 25'b10001000_11011011_01100011_1;
      patterns[35038] = 25'b10001000_11011100_01100100_1;
      patterns[35039] = 25'b10001000_11011101_01100101_1;
      patterns[35040] = 25'b10001000_11011110_01100110_1;
      patterns[35041] = 25'b10001000_11011111_01100111_1;
      patterns[35042] = 25'b10001000_11100000_01101000_1;
      patterns[35043] = 25'b10001000_11100001_01101001_1;
      patterns[35044] = 25'b10001000_11100010_01101010_1;
      patterns[35045] = 25'b10001000_11100011_01101011_1;
      patterns[35046] = 25'b10001000_11100100_01101100_1;
      patterns[35047] = 25'b10001000_11100101_01101101_1;
      patterns[35048] = 25'b10001000_11100110_01101110_1;
      patterns[35049] = 25'b10001000_11100111_01101111_1;
      patterns[35050] = 25'b10001000_11101000_01110000_1;
      patterns[35051] = 25'b10001000_11101001_01110001_1;
      patterns[35052] = 25'b10001000_11101010_01110010_1;
      patterns[35053] = 25'b10001000_11101011_01110011_1;
      patterns[35054] = 25'b10001000_11101100_01110100_1;
      patterns[35055] = 25'b10001000_11101101_01110101_1;
      patterns[35056] = 25'b10001000_11101110_01110110_1;
      patterns[35057] = 25'b10001000_11101111_01110111_1;
      patterns[35058] = 25'b10001000_11110000_01111000_1;
      patterns[35059] = 25'b10001000_11110001_01111001_1;
      patterns[35060] = 25'b10001000_11110010_01111010_1;
      patterns[35061] = 25'b10001000_11110011_01111011_1;
      patterns[35062] = 25'b10001000_11110100_01111100_1;
      patterns[35063] = 25'b10001000_11110101_01111101_1;
      patterns[35064] = 25'b10001000_11110110_01111110_1;
      patterns[35065] = 25'b10001000_11110111_01111111_1;
      patterns[35066] = 25'b10001000_11111000_10000000_1;
      patterns[35067] = 25'b10001000_11111001_10000001_1;
      patterns[35068] = 25'b10001000_11111010_10000010_1;
      patterns[35069] = 25'b10001000_11111011_10000011_1;
      patterns[35070] = 25'b10001000_11111100_10000100_1;
      patterns[35071] = 25'b10001000_11111101_10000101_1;
      patterns[35072] = 25'b10001000_11111110_10000110_1;
      patterns[35073] = 25'b10001000_11111111_10000111_1;
      patterns[35074] = 25'b10001001_00000000_10001001_0;
      patterns[35075] = 25'b10001001_00000001_10001010_0;
      patterns[35076] = 25'b10001001_00000010_10001011_0;
      patterns[35077] = 25'b10001001_00000011_10001100_0;
      patterns[35078] = 25'b10001001_00000100_10001101_0;
      patterns[35079] = 25'b10001001_00000101_10001110_0;
      patterns[35080] = 25'b10001001_00000110_10001111_0;
      patterns[35081] = 25'b10001001_00000111_10010000_0;
      patterns[35082] = 25'b10001001_00001000_10010001_0;
      patterns[35083] = 25'b10001001_00001001_10010010_0;
      patterns[35084] = 25'b10001001_00001010_10010011_0;
      patterns[35085] = 25'b10001001_00001011_10010100_0;
      patterns[35086] = 25'b10001001_00001100_10010101_0;
      patterns[35087] = 25'b10001001_00001101_10010110_0;
      patterns[35088] = 25'b10001001_00001110_10010111_0;
      patterns[35089] = 25'b10001001_00001111_10011000_0;
      patterns[35090] = 25'b10001001_00010000_10011001_0;
      patterns[35091] = 25'b10001001_00010001_10011010_0;
      patterns[35092] = 25'b10001001_00010010_10011011_0;
      patterns[35093] = 25'b10001001_00010011_10011100_0;
      patterns[35094] = 25'b10001001_00010100_10011101_0;
      patterns[35095] = 25'b10001001_00010101_10011110_0;
      patterns[35096] = 25'b10001001_00010110_10011111_0;
      patterns[35097] = 25'b10001001_00010111_10100000_0;
      patterns[35098] = 25'b10001001_00011000_10100001_0;
      patterns[35099] = 25'b10001001_00011001_10100010_0;
      patterns[35100] = 25'b10001001_00011010_10100011_0;
      patterns[35101] = 25'b10001001_00011011_10100100_0;
      patterns[35102] = 25'b10001001_00011100_10100101_0;
      patterns[35103] = 25'b10001001_00011101_10100110_0;
      patterns[35104] = 25'b10001001_00011110_10100111_0;
      patterns[35105] = 25'b10001001_00011111_10101000_0;
      patterns[35106] = 25'b10001001_00100000_10101001_0;
      patterns[35107] = 25'b10001001_00100001_10101010_0;
      patterns[35108] = 25'b10001001_00100010_10101011_0;
      patterns[35109] = 25'b10001001_00100011_10101100_0;
      patterns[35110] = 25'b10001001_00100100_10101101_0;
      patterns[35111] = 25'b10001001_00100101_10101110_0;
      patterns[35112] = 25'b10001001_00100110_10101111_0;
      patterns[35113] = 25'b10001001_00100111_10110000_0;
      patterns[35114] = 25'b10001001_00101000_10110001_0;
      patterns[35115] = 25'b10001001_00101001_10110010_0;
      patterns[35116] = 25'b10001001_00101010_10110011_0;
      patterns[35117] = 25'b10001001_00101011_10110100_0;
      patterns[35118] = 25'b10001001_00101100_10110101_0;
      patterns[35119] = 25'b10001001_00101101_10110110_0;
      patterns[35120] = 25'b10001001_00101110_10110111_0;
      patterns[35121] = 25'b10001001_00101111_10111000_0;
      patterns[35122] = 25'b10001001_00110000_10111001_0;
      patterns[35123] = 25'b10001001_00110001_10111010_0;
      patterns[35124] = 25'b10001001_00110010_10111011_0;
      patterns[35125] = 25'b10001001_00110011_10111100_0;
      patterns[35126] = 25'b10001001_00110100_10111101_0;
      patterns[35127] = 25'b10001001_00110101_10111110_0;
      patterns[35128] = 25'b10001001_00110110_10111111_0;
      patterns[35129] = 25'b10001001_00110111_11000000_0;
      patterns[35130] = 25'b10001001_00111000_11000001_0;
      patterns[35131] = 25'b10001001_00111001_11000010_0;
      patterns[35132] = 25'b10001001_00111010_11000011_0;
      patterns[35133] = 25'b10001001_00111011_11000100_0;
      patterns[35134] = 25'b10001001_00111100_11000101_0;
      patterns[35135] = 25'b10001001_00111101_11000110_0;
      patterns[35136] = 25'b10001001_00111110_11000111_0;
      patterns[35137] = 25'b10001001_00111111_11001000_0;
      patterns[35138] = 25'b10001001_01000000_11001001_0;
      patterns[35139] = 25'b10001001_01000001_11001010_0;
      patterns[35140] = 25'b10001001_01000010_11001011_0;
      patterns[35141] = 25'b10001001_01000011_11001100_0;
      patterns[35142] = 25'b10001001_01000100_11001101_0;
      patterns[35143] = 25'b10001001_01000101_11001110_0;
      patterns[35144] = 25'b10001001_01000110_11001111_0;
      patterns[35145] = 25'b10001001_01000111_11010000_0;
      patterns[35146] = 25'b10001001_01001000_11010001_0;
      patterns[35147] = 25'b10001001_01001001_11010010_0;
      patterns[35148] = 25'b10001001_01001010_11010011_0;
      patterns[35149] = 25'b10001001_01001011_11010100_0;
      patterns[35150] = 25'b10001001_01001100_11010101_0;
      patterns[35151] = 25'b10001001_01001101_11010110_0;
      patterns[35152] = 25'b10001001_01001110_11010111_0;
      patterns[35153] = 25'b10001001_01001111_11011000_0;
      patterns[35154] = 25'b10001001_01010000_11011001_0;
      patterns[35155] = 25'b10001001_01010001_11011010_0;
      patterns[35156] = 25'b10001001_01010010_11011011_0;
      patterns[35157] = 25'b10001001_01010011_11011100_0;
      patterns[35158] = 25'b10001001_01010100_11011101_0;
      patterns[35159] = 25'b10001001_01010101_11011110_0;
      patterns[35160] = 25'b10001001_01010110_11011111_0;
      patterns[35161] = 25'b10001001_01010111_11100000_0;
      patterns[35162] = 25'b10001001_01011000_11100001_0;
      patterns[35163] = 25'b10001001_01011001_11100010_0;
      patterns[35164] = 25'b10001001_01011010_11100011_0;
      patterns[35165] = 25'b10001001_01011011_11100100_0;
      patterns[35166] = 25'b10001001_01011100_11100101_0;
      patterns[35167] = 25'b10001001_01011101_11100110_0;
      patterns[35168] = 25'b10001001_01011110_11100111_0;
      patterns[35169] = 25'b10001001_01011111_11101000_0;
      patterns[35170] = 25'b10001001_01100000_11101001_0;
      patterns[35171] = 25'b10001001_01100001_11101010_0;
      patterns[35172] = 25'b10001001_01100010_11101011_0;
      patterns[35173] = 25'b10001001_01100011_11101100_0;
      patterns[35174] = 25'b10001001_01100100_11101101_0;
      patterns[35175] = 25'b10001001_01100101_11101110_0;
      patterns[35176] = 25'b10001001_01100110_11101111_0;
      patterns[35177] = 25'b10001001_01100111_11110000_0;
      patterns[35178] = 25'b10001001_01101000_11110001_0;
      patterns[35179] = 25'b10001001_01101001_11110010_0;
      patterns[35180] = 25'b10001001_01101010_11110011_0;
      patterns[35181] = 25'b10001001_01101011_11110100_0;
      patterns[35182] = 25'b10001001_01101100_11110101_0;
      patterns[35183] = 25'b10001001_01101101_11110110_0;
      patterns[35184] = 25'b10001001_01101110_11110111_0;
      patterns[35185] = 25'b10001001_01101111_11111000_0;
      patterns[35186] = 25'b10001001_01110000_11111001_0;
      patterns[35187] = 25'b10001001_01110001_11111010_0;
      patterns[35188] = 25'b10001001_01110010_11111011_0;
      patterns[35189] = 25'b10001001_01110011_11111100_0;
      patterns[35190] = 25'b10001001_01110100_11111101_0;
      patterns[35191] = 25'b10001001_01110101_11111110_0;
      patterns[35192] = 25'b10001001_01110110_11111111_0;
      patterns[35193] = 25'b10001001_01110111_00000000_1;
      patterns[35194] = 25'b10001001_01111000_00000001_1;
      patterns[35195] = 25'b10001001_01111001_00000010_1;
      patterns[35196] = 25'b10001001_01111010_00000011_1;
      patterns[35197] = 25'b10001001_01111011_00000100_1;
      patterns[35198] = 25'b10001001_01111100_00000101_1;
      patterns[35199] = 25'b10001001_01111101_00000110_1;
      patterns[35200] = 25'b10001001_01111110_00000111_1;
      patterns[35201] = 25'b10001001_01111111_00001000_1;
      patterns[35202] = 25'b10001001_10000000_00001001_1;
      patterns[35203] = 25'b10001001_10000001_00001010_1;
      patterns[35204] = 25'b10001001_10000010_00001011_1;
      patterns[35205] = 25'b10001001_10000011_00001100_1;
      patterns[35206] = 25'b10001001_10000100_00001101_1;
      patterns[35207] = 25'b10001001_10000101_00001110_1;
      patterns[35208] = 25'b10001001_10000110_00001111_1;
      patterns[35209] = 25'b10001001_10000111_00010000_1;
      patterns[35210] = 25'b10001001_10001000_00010001_1;
      patterns[35211] = 25'b10001001_10001001_00010010_1;
      patterns[35212] = 25'b10001001_10001010_00010011_1;
      patterns[35213] = 25'b10001001_10001011_00010100_1;
      patterns[35214] = 25'b10001001_10001100_00010101_1;
      patterns[35215] = 25'b10001001_10001101_00010110_1;
      patterns[35216] = 25'b10001001_10001110_00010111_1;
      patterns[35217] = 25'b10001001_10001111_00011000_1;
      patterns[35218] = 25'b10001001_10010000_00011001_1;
      patterns[35219] = 25'b10001001_10010001_00011010_1;
      patterns[35220] = 25'b10001001_10010010_00011011_1;
      patterns[35221] = 25'b10001001_10010011_00011100_1;
      patterns[35222] = 25'b10001001_10010100_00011101_1;
      patterns[35223] = 25'b10001001_10010101_00011110_1;
      patterns[35224] = 25'b10001001_10010110_00011111_1;
      patterns[35225] = 25'b10001001_10010111_00100000_1;
      patterns[35226] = 25'b10001001_10011000_00100001_1;
      patterns[35227] = 25'b10001001_10011001_00100010_1;
      patterns[35228] = 25'b10001001_10011010_00100011_1;
      patterns[35229] = 25'b10001001_10011011_00100100_1;
      patterns[35230] = 25'b10001001_10011100_00100101_1;
      patterns[35231] = 25'b10001001_10011101_00100110_1;
      patterns[35232] = 25'b10001001_10011110_00100111_1;
      patterns[35233] = 25'b10001001_10011111_00101000_1;
      patterns[35234] = 25'b10001001_10100000_00101001_1;
      patterns[35235] = 25'b10001001_10100001_00101010_1;
      patterns[35236] = 25'b10001001_10100010_00101011_1;
      patterns[35237] = 25'b10001001_10100011_00101100_1;
      patterns[35238] = 25'b10001001_10100100_00101101_1;
      patterns[35239] = 25'b10001001_10100101_00101110_1;
      patterns[35240] = 25'b10001001_10100110_00101111_1;
      patterns[35241] = 25'b10001001_10100111_00110000_1;
      patterns[35242] = 25'b10001001_10101000_00110001_1;
      patterns[35243] = 25'b10001001_10101001_00110010_1;
      patterns[35244] = 25'b10001001_10101010_00110011_1;
      patterns[35245] = 25'b10001001_10101011_00110100_1;
      patterns[35246] = 25'b10001001_10101100_00110101_1;
      patterns[35247] = 25'b10001001_10101101_00110110_1;
      patterns[35248] = 25'b10001001_10101110_00110111_1;
      patterns[35249] = 25'b10001001_10101111_00111000_1;
      patterns[35250] = 25'b10001001_10110000_00111001_1;
      patterns[35251] = 25'b10001001_10110001_00111010_1;
      patterns[35252] = 25'b10001001_10110010_00111011_1;
      patterns[35253] = 25'b10001001_10110011_00111100_1;
      patterns[35254] = 25'b10001001_10110100_00111101_1;
      patterns[35255] = 25'b10001001_10110101_00111110_1;
      patterns[35256] = 25'b10001001_10110110_00111111_1;
      patterns[35257] = 25'b10001001_10110111_01000000_1;
      patterns[35258] = 25'b10001001_10111000_01000001_1;
      patterns[35259] = 25'b10001001_10111001_01000010_1;
      patterns[35260] = 25'b10001001_10111010_01000011_1;
      patterns[35261] = 25'b10001001_10111011_01000100_1;
      patterns[35262] = 25'b10001001_10111100_01000101_1;
      patterns[35263] = 25'b10001001_10111101_01000110_1;
      patterns[35264] = 25'b10001001_10111110_01000111_1;
      patterns[35265] = 25'b10001001_10111111_01001000_1;
      patterns[35266] = 25'b10001001_11000000_01001001_1;
      patterns[35267] = 25'b10001001_11000001_01001010_1;
      patterns[35268] = 25'b10001001_11000010_01001011_1;
      patterns[35269] = 25'b10001001_11000011_01001100_1;
      patterns[35270] = 25'b10001001_11000100_01001101_1;
      patterns[35271] = 25'b10001001_11000101_01001110_1;
      patterns[35272] = 25'b10001001_11000110_01001111_1;
      patterns[35273] = 25'b10001001_11000111_01010000_1;
      patterns[35274] = 25'b10001001_11001000_01010001_1;
      patterns[35275] = 25'b10001001_11001001_01010010_1;
      patterns[35276] = 25'b10001001_11001010_01010011_1;
      patterns[35277] = 25'b10001001_11001011_01010100_1;
      patterns[35278] = 25'b10001001_11001100_01010101_1;
      patterns[35279] = 25'b10001001_11001101_01010110_1;
      patterns[35280] = 25'b10001001_11001110_01010111_1;
      patterns[35281] = 25'b10001001_11001111_01011000_1;
      patterns[35282] = 25'b10001001_11010000_01011001_1;
      patterns[35283] = 25'b10001001_11010001_01011010_1;
      patterns[35284] = 25'b10001001_11010010_01011011_1;
      patterns[35285] = 25'b10001001_11010011_01011100_1;
      patterns[35286] = 25'b10001001_11010100_01011101_1;
      patterns[35287] = 25'b10001001_11010101_01011110_1;
      patterns[35288] = 25'b10001001_11010110_01011111_1;
      patterns[35289] = 25'b10001001_11010111_01100000_1;
      patterns[35290] = 25'b10001001_11011000_01100001_1;
      patterns[35291] = 25'b10001001_11011001_01100010_1;
      patterns[35292] = 25'b10001001_11011010_01100011_1;
      patterns[35293] = 25'b10001001_11011011_01100100_1;
      patterns[35294] = 25'b10001001_11011100_01100101_1;
      patterns[35295] = 25'b10001001_11011101_01100110_1;
      patterns[35296] = 25'b10001001_11011110_01100111_1;
      patterns[35297] = 25'b10001001_11011111_01101000_1;
      patterns[35298] = 25'b10001001_11100000_01101001_1;
      patterns[35299] = 25'b10001001_11100001_01101010_1;
      patterns[35300] = 25'b10001001_11100010_01101011_1;
      patterns[35301] = 25'b10001001_11100011_01101100_1;
      patterns[35302] = 25'b10001001_11100100_01101101_1;
      patterns[35303] = 25'b10001001_11100101_01101110_1;
      patterns[35304] = 25'b10001001_11100110_01101111_1;
      patterns[35305] = 25'b10001001_11100111_01110000_1;
      patterns[35306] = 25'b10001001_11101000_01110001_1;
      patterns[35307] = 25'b10001001_11101001_01110010_1;
      patterns[35308] = 25'b10001001_11101010_01110011_1;
      patterns[35309] = 25'b10001001_11101011_01110100_1;
      patterns[35310] = 25'b10001001_11101100_01110101_1;
      patterns[35311] = 25'b10001001_11101101_01110110_1;
      patterns[35312] = 25'b10001001_11101110_01110111_1;
      patterns[35313] = 25'b10001001_11101111_01111000_1;
      patterns[35314] = 25'b10001001_11110000_01111001_1;
      patterns[35315] = 25'b10001001_11110001_01111010_1;
      patterns[35316] = 25'b10001001_11110010_01111011_1;
      patterns[35317] = 25'b10001001_11110011_01111100_1;
      patterns[35318] = 25'b10001001_11110100_01111101_1;
      patterns[35319] = 25'b10001001_11110101_01111110_1;
      patterns[35320] = 25'b10001001_11110110_01111111_1;
      patterns[35321] = 25'b10001001_11110111_10000000_1;
      patterns[35322] = 25'b10001001_11111000_10000001_1;
      patterns[35323] = 25'b10001001_11111001_10000010_1;
      patterns[35324] = 25'b10001001_11111010_10000011_1;
      patterns[35325] = 25'b10001001_11111011_10000100_1;
      patterns[35326] = 25'b10001001_11111100_10000101_1;
      patterns[35327] = 25'b10001001_11111101_10000110_1;
      patterns[35328] = 25'b10001001_11111110_10000111_1;
      patterns[35329] = 25'b10001001_11111111_10001000_1;
      patterns[35330] = 25'b10001010_00000000_10001010_0;
      patterns[35331] = 25'b10001010_00000001_10001011_0;
      patterns[35332] = 25'b10001010_00000010_10001100_0;
      patterns[35333] = 25'b10001010_00000011_10001101_0;
      patterns[35334] = 25'b10001010_00000100_10001110_0;
      patterns[35335] = 25'b10001010_00000101_10001111_0;
      patterns[35336] = 25'b10001010_00000110_10010000_0;
      patterns[35337] = 25'b10001010_00000111_10010001_0;
      patterns[35338] = 25'b10001010_00001000_10010010_0;
      patterns[35339] = 25'b10001010_00001001_10010011_0;
      patterns[35340] = 25'b10001010_00001010_10010100_0;
      patterns[35341] = 25'b10001010_00001011_10010101_0;
      patterns[35342] = 25'b10001010_00001100_10010110_0;
      patterns[35343] = 25'b10001010_00001101_10010111_0;
      patterns[35344] = 25'b10001010_00001110_10011000_0;
      patterns[35345] = 25'b10001010_00001111_10011001_0;
      patterns[35346] = 25'b10001010_00010000_10011010_0;
      patterns[35347] = 25'b10001010_00010001_10011011_0;
      patterns[35348] = 25'b10001010_00010010_10011100_0;
      patterns[35349] = 25'b10001010_00010011_10011101_0;
      patterns[35350] = 25'b10001010_00010100_10011110_0;
      patterns[35351] = 25'b10001010_00010101_10011111_0;
      patterns[35352] = 25'b10001010_00010110_10100000_0;
      patterns[35353] = 25'b10001010_00010111_10100001_0;
      patterns[35354] = 25'b10001010_00011000_10100010_0;
      patterns[35355] = 25'b10001010_00011001_10100011_0;
      patterns[35356] = 25'b10001010_00011010_10100100_0;
      patterns[35357] = 25'b10001010_00011011_10100101_0;
      patterns[35358] = 25'b10001010_00011100_10100110_0;
      patterns[35359] = 25'b10001010_00011101_10100111_0;
      patterns[35360] = 25'b10001010_00011110_10101000_0;
      patterns[35361] = 25'b10001010_00011111_10101001_0;
      patterns[35362] = 25'b10001010_00100000_10101010_0;
      patterns[35363] = 25'b10001010_00100001_10101011_0;
      patterns[35364] = 25'b10001010_00100010_10101100_0;
      patterns[35365] = 25'b10001010_00100011_10101101_0;
      patterns[35366] = 25'b10001010_00100100_10101110_0;
      patterns[35367] = 25'b10001010_00100101_10101111_0;
      patterns[35368] = 25'b10001010_00100110_10110000_0;
      patterns[35369] = 25'b10001010_00100111_10110001_0;
      patterns[35370] = 25'b10001010_00101000_10110010_0;
      patterns[35371] = 25'b10001010_00101001_10110011_0;
      patterns[35372] = 25'b10001010_00101010_10110100_0;
      patterns[35373] = 25'b10001010_00101011_10110101_0;
      patterns[35374] = 25'b10001010_00101100_10110110_0;
      patterns[35375] = 25'b10001010_00101101_10110111_0;
      patterns[35376] = 25'b10001010_00101110_10111000_0;
      patterns[35377] = 25'b10001010_00101111_10111001_0;
      patterns[35378] = 25'b10001010_00110000_10111010_0;
      patterns[35379] = 25'b10001010_00110001_10111011_0;
      patterns[35380] = 25'b10001010_00110010_10111100_0;
      patterns[35381] = 25'b10001010_00110011_10111101_0;
      patterns[35382] = 25'b10001010_00110100_10111110_0;
      patterns[35383] = 25'b10001010_00110101_10111111_0;
      patterns[35384] = 25'b10001010_00110110_11000000_0;
      patterns[35385] = 25'b10001010_00110111_11000001_0;
      patterns[35386] = 25'b10001010_00111000_11000010_0;
      patterns[35387] = 25'b10001010_00111001_11000011_0;
      patterns[35388] = 25'b10001010_00111010_11000100_0;
      patterns[35389] = 25'b10001010_00111011_11000101_0;
      patterns[35390] = 25'b10001010_00111100_11000110_0;
      patterns[35391] = 25'b10001010_00111101_11000111_0;
      patterns[35392] = 25'b10001010_00111110_11001000_0;
      patterns[35393] = 25'b10001010_00111111_11001001_0;
      patterns[35394] = 25'b10001010_01000000_11001010_0;
      patterns[35395] = 25'b10001010_01000001_11001011_0;
      patterns[35396] = 25'b10001010_01000010_11001100_0;
      patterns[35397] = 25'b10001010_01000011_11001101_0;
      patterns[35398] = 25'b10001010_01000100_11001110_0;
      patterns[35399] = 25'b10001010_01000101_11001111_0;
      patterns[35400] = 25'b10001010_01000110_11010000_0;
      patterns[35401] = 25'b10001010_01000111_11010001_0;
      patterns[35402] = 25'b10001010_01001000_11010010_0;
      patterns[35403] = 25'b10001010_01001001_11010011_0;
      patterns[35404] = 25'b10001010_01001010_11010100_0;
      patterns[35405] = 25'b10001010_01001011_11010101_0;
      patterns[35406] = 25'b10001010_01001100_11010110_0;
      patterns[35407] = 25'b10001010_01001101_11010111_0;
      patterns[35408] = 25'b10001010_01001110_11011000_0;
      patterns[35409] = 25'b10001010_01001111_11011001_0;
      patterns[35410] = 25'b10001010_01010000_11011010_0;
      patterns[35411] = 25'b10001010_01010001_11011011_0;
      patterns[35412] = 25'b10001010_01010010_11011100_0;
      patterns[35413] = 25'b10001010_01010011_11011101_0;
      patterns[35414] = 25'b10001010_01010100_11011110_0;
      patterns[35415] = 25'b10001010_01010101_11011111_0;
      patterns[35416] = 25'b10001010_01010110_11100000_0;
      patterns[35417] = 25'b10001010_01010111_11100001_0;
      patterns[35418] = 25'b10001010_01011000_11100010_0;
      patterns[35419] = 25'b10001010_01011001_11100011_0;
      patterns[35420] = 25'b10001010_01011010_11100100_0;
      patterns[35421] = 25'b10001010_01011011_11100101_0;
      patterns[35422] = 25'b10001010_01011100_11100110_0;
      patterns[35423] = 25'b10001010_01011101_11100111_0;
      patterns[35424] = 25'b10001010_01011110_11101000_0;
      patterns[35425] = 25'b10001010_01011111_11101001_0;
      patterns[35426] = 25'b10001010_01100000_11101010_0;
      patterns[35427] = 25'b10001010_01100001_11101011_0;
      patterns[35428] = 25'b10001010_01100010_11101100_0;
      patterns[35429] = 25'b10001010_01100011_11101101_0;
      patterns[35430] = 25'b10001010_01100100_11101110_0;
      patterns[35431] = 25'b10001010_01100101_11101111_0;
      patterns[35432] = 25'b10001010_01100110_11110000_0;
      patterns[35433] = 25'b10001010_01100111_11110001_0;
      patterns[35434] = 25'b10001010_01101000_11110010_0;
      patterns[35435] = 25'b10001010_01101001_11110011_0;
      patterns[35436] = 25'b10001010_01101010_11110100_0;
      patterns[35437] = 25'b10001010_01101011_11110101_0;
      patterns[35438] = 25'b10001010_01101100_11110110_0;
      patterns[35439] = 25'b10001010_01101101_11110111_0;
      patterns[35440] = 25'b10001010_01101110_11111000_0;
      patterns[35441] = 25'b10001010_01101111_11111001_0;
      patterns[35442] = 25'b10001010_01110000_11111010_0;
      patterns[35443] = 25'b10001010_01110001_11111011_0;
      patterns[35444] = 25'b10001010_01110010_11111100_0;
      patterns[35445] = 25'b10001010_01110011_11111101_0;
      patterns[35446] = 25'b10001010_01110100_11111110_0;
      patterns[35447] = 25'b10001010_01110101_11111111_0;
      patterns[35448] = 25'b10001010_01110110_00000000_1;
      patterns[35449] = 25'b10001010_01110111_00000001_1;
      patterns[35450] = 25'b10001010_01111000_00000010_1;
      patterns[35451] = 25'b10001010_01111001_00000011_1;
      patterns[35452] = 25'b10001010_01111010_00000100_1;
      patterns[35453] = 25'b10001010_01111011_00000101_1;
      patterns[35454] = 25'b10001010_01111100_00000110_1;
      patterns[35455] = 25'b10001010_01111101_00000111_1;
      patterns[35456] = 25'b10001010_01111110_00001000_1;
      patterns[35457] = 25'b10001010_01111111_00001001_1;
      patterns[35458] = 25'b10001010_10000000_00001010_1;
      patterns[35459] = 25'b10001010_10000001_00001011_1;
      patterns[35460] = 25'b10001010_10000010_00001100_1;
      patterns[35461] = 25'b10001010_10000011_00001101_1;
      patterns[35462] = 25'b10001010_10000100_00001110_1;
      patterns[35463] = 25'b10001010_10000101_00001111_1;
      patterns[35464] = 25'b10001010_10000110_00010000_1;
      patterns[35465] = 25'b10001010_10000111_00010001_1;
      patterns[35466] = 25'b10001010_10001000_00010010_1;
      patterns[35467] = 25'b10001010_10001001_00010011_1;
      patterns[35468] = 25'b10001010_10001010_00010100_1;
      patterns[35469] = 25'b10001010_10001011_00010101_1;
      patterns[35470] = 25'b10001010_10001100_00010110_1;
      patterns[35471] = 25'b10001010_10001101_00010111_1;
      patterns[35472] = 25'b10001010_10001110_00011000_1;
      patterns[35473] = 25'b10001010_10001111_00011001_1;
      patterns[35474] = 25'b10001010_10010000_00011010_1;
      patterns[35475] = 25'b10001010_10010001_00011011_1;
      patterns[35476] = 25'b10001010_10010010_00011100_1;
      patterns[35477] = 25'b10001010_10010011_00011101_1;
      patterns[35478] = 25'b10001010_10010100_00011110_1;
      patterns[35479] = 25'b10001010_10010101_00011111_1;
      patterns[35480] = 25'b10001010_10010110_00100000_1;
      patterns[35481] = 25'b10001010_10010111_00100001_1;
      patterns[35482] = 25'b10001010_10011000_00100010_1;
      patterns[35483] = 25'b10001010_10011001_00100011_1;
      patterns[35484] = 25'b10001010_10011010_00100100_1;
      patterns[35485] = 25'b10001010_10011011_00100101_1;
      patterns[35486] = 25'b10001010_10011100_00100110_1;
      patterns[35487] = 25'b10001010_10011101_00100111_1;
      patterns[35488] = 25'b10001010_10011110_00101000_1;
      patterns[35489] = 25'b10001010_10011111_00101001_1;
      patterns[35490] = 25'b10001010_10100000_00101010_1;
      patterns[35491] = 25'b10001010_10100001_00101011_1;
      patterns[35492] = 25'b10001010_10100010_00101100_1;
      patterns[35493] = 25'b10001010_10100011_00101101_1;
      patterns[35494] = 25'b10001010_10100100_00101110_1;
      patterns[35495] = 25'b10001010_10100101_00101111_1;
      patterns[35496] = 25'b10001010_10100110_00110000_1;
      patterns[35497] = 25'b10001010_10100111_00110001_1;
      patterns[35498] = 25'b10001010_10101000_00110010_1;
      patterns[35499] = 25'b10001010_10101001_00110011_1;
      patterns[35500] = 25'b10001010_10101010_00110100_1;
      patterns[35501] = 25'b10001010_10101011_00110101_1;
      patterns[35502] = 25'b10001010_10101100_00110110_1;
      patterns[35503] = 25'b10001010_10101101_00110111_1;
      patterns[35504] = 25'b10001010_10101110_00111000_1;
      patterns[35505] = 25'b10001010_10101111_00111001_1;
      patterns[35506] = 25'b10001010_10110000_00111010_1;
      patterns[35507] = 25'b10001010_10110001_00111011_1;
      patterns[35508] = 25'b10001010_10110010_00111100_1;
      patterns[35509] = 25'b10001010_10110011_00111101_1;
      patterns[35510] = 25'b10001010_10110100_00111110_1;
      patterns[35511] = 25'b10001010_10110101_00111111_1;
      patterns[35512] = 25'b10001010_10110110_01000000_1;
      patterns[35513] = 25'b10001010_10110111_01000001_1;
      patterns[35514] = 25'b10001010_10111000_01000010_1;
      patterns[35515] = 25'b10001010_10111001_01000011_1;
      patterns[35516] = 25'b10001010_10111010_01000100_1;
      patterns[35517] = 25'b10001010_10111011_01000101_1;
      patterns[35518] = 25'b10001010_10111100_01000110_1;
      patterns[35519] = 25'b10001010_10111101_01000111_1;
      patterns[35520] = 25'b10001010_10111110_01001000_1;
      patterns[35521] = 25'b10001010_10111111_01001001_1;
      patterns[35522] = 25'b10001010_11000000_01001010_1;
      patterns[35523] = 25'b10001010_11000001_01001011_1;
      patterns[35524] = 25'b10001010_11000010_01001100_1;
      patterns[35525] = 25'b10001010_11000011_01001101_1;
      patterns[35526] = 25'b10001010_11000100_01001110_1;
      patterns[35527] = 25'b10001010_11000101_01001111_1;
      patterns[35528] = 25'b10001010_11000110_01010000_1;
      patterns[35529] = 25'b10001010_11000111_01010001_1;
      patterns[35530] = 25'b10001010_11001000_01010010_1;
      patterns[35531] = 25'b10001010_11001001_01010011_1;
      patterns[35532] = 25'b10001010_11001010_01010100_1;
      patterns[35533] = 25'b10001010_11001011_01010101_1;
      patterns[35534] = 25'b10001010_11001100_01010110_1;
      patterns[35535] = 25'b10001010_11001101_01010111_1;
      patterns[35536] = 25'b10001010_11001110_01011000_1;
      patterns[35537] = 25'b10001010_11001111_01011001_1;
      patterns[35538] = 25'b10001010_11010000_01011010_1;
      patterns[35539] = 25'b10001010_11010001_01011011_1;
      patterns[35540] = 25'b10001010_11010010_01011100_1;
      patterns[35541] = 25'b10001010_11010011_01011101_1;
      patterns[35542] = 25'b10001010_11010100_01011110_1;
      patterns[35543] = 25'b10001010_11010101_01011111_1;
      patterns[35544] = 25'b10001010_11010110_01100000_1;
      patterns[35545] = 25'b10001010_11010111_01100001_1;
      patterns[35546] = 25'b10001010_11011000_01100010_1;
      patterns[35547] = 25'b10001010_11011001_01100011_1;
      patterns[35548] = 25'b10001010_11011010_01100100_1;
      patterns[35549] = 25'b10001010_11011011_01100101_1;
      patterns[35550] = 25'b10001010_11011100_01100110_1;
      patterns[35551] = 25'b10001010_11011101_01100111_1;
      patterns[35552] = 25'b10001010_11011110_01101000_1;
      patterns[35553] = 25'b10001010_11011111_01101001_1;
      patterns[35554] = 25'b10001010_11100000_01101010_1;
      patterns[35555] = 25'b10001010_11100001_01101011_1;
      patterns[35556] = 25'b10001010_11100010_01101100_1;
      patterns[35557] = 25'b10001010_11100011_01101101_1;
      patterns[35558] = 25'b10001010_11100100_01101110_1;
      patterns[35559] = 25'b10001010_11100101_01101111_1;
      patterns[35560] = 25'b10001010_11100110_01110000_1;
      patterns[35561] = 25'b10001010_11100111_01110001_1;
      patterns[35562] = 25'b10001010_11101000_01110010_1;
      patterns[35563] = 25'b10001010_11101001_01110011_1;
      patterns[35564] = 25'b10001010_11101010_01110100_1;
      patterns[35565] = 25'b10001010_11101011_01110101_1;
      patterns[35566] = 25'b10001010_11101100_01110110_1;
      patterns[35567] = 25'b10001010_11101101_01110111_1;
      patterns[35568] = 25'b10001010_11101110_01111000_1;
      patterns[35569] = 25'b10001010_11101111_01111001_1;
      patterns[35570] = 25'b10001010_11110000_01111010_1;
      patterns[35571] = 25'b10001010_11110001_01111011_1;
      patterns[35572] = 25'b10001010_11110010_01111100_1;
      patterns[35573] = 25'b10001010_11110011_01111101_1;
      patterns[35574] = 25'b10001010_11110100_01111110_1;
      patterns[35575] = 25'b10001010_11110101_01111111_1;
      patterns[35576] = 25'b10001010_11110110_10000000_1;
      patterns[35577] = 25'b10001010_11110111_10000001_1;
      patterns[35578] = 25'b10001010_11111000_10000010_1;
      patterns[35579] = 25'b10001010_11111001_10000011_1;
      patterns[35580] = 25'b10001010_11111010_10000100_1;
      patterns[35581] = 25'b10001010_11111011_10000101_1;
      patterns[35582] = 25'b10001010_11111100_10000110_1;
      patterns[35583] = 25'b10001010_11111101_10000111_1;
      patterns[35584] = 25'b10001010_11111110_10001000_1;
      patterns[35585] = 25'b10001010_11111111_10001001_1;
      patterns[35586] = 25'b10001011_00000000_10001011_0;
      patterns[35587] = 25'b10001011_00000001_10001100_0;
      patterns[35588] = 25'b10001011_00000010_10001101_0;
      patterns[35589] = 25'b10001011_00000011_10001110_0;
      patterns[35590] = 25'b10001011_00000100_10001111_0;
      patterns[35591] = 25'b10001011_00000101_10010000_0;
      patterns[35592] = 25'b10001011_00000110_10010001_0;
      patterns[35593] = 25'b10001011_00000111_10010010_0;
      patterns[35594] = 25'b10001011_00001000_10010011_0;
      patterns[35595] = 25'b10001011_00001001_10010100_0;
      patterns[35596] = 25'b10001011_00001010_10010101_0;
      patterns[35597] = 25'b10001011_00001011_10010110_0;
      patterns[35598] = 25'b10001011_00001100_10010111_0;
      patterns[35599] = 25'b10001011_00001101_10011000_0;
      patterns[35600] = 25'b10001011_00001110_10011001_0;
      patterns[35601] = 25'b10001011_00001111_10011010_0;
      patterns[35602] = 25'b10001011_00010000_10011011_0;
      patterns[35603] = 25'b10001011_00010001_10011100_0;
      patterns[35604] = 25'b10001011_00010010_10011101_0;
      patterns[35605] = 25'b10001011_00010011_10011110_0;
      patterns[35606] = 25'b10001011_00010100_10011111_0;
      patterns[35607] = 25'b10001011_00010101_10100000_0;
      patterns[35608] = 25'b10001011_00010110_10100001_0;
      patterns[35609] = 25'b10001011_00010111_10100010_0;
      patterns[35610] = 25'b10001011_00011000_10100011_0;
      patterns[35611] = 25'b10001011_00011001_10100100_0;
      patterns[35612] = 25'b10001011_00011010_10100101_0;
      patterns[35613] = 25'b10001011_00011011_10100110_0;
      patterns[35614] = 25'b10001011_00011100_10100111_0;
      patterns[35615] = 25'b10001011_00011101_10101000_0;
      patterns[35616] = 25'b10001011_00011110_10101001_0;
      patterns[35617] = 25'b10001011_00011111_10101010_0;
      patterns[35618] = 25'b10001011_00100000_10101011_0;
      patterns[35619] = 25'b10001011_00100001_10101100_0;
      patterns[35620] = 25'b10001011_00100010_10101101_0;
      patterns[35621] = 25'b10001011_00100011_10101110_0;
      patterns[35622] = 25'b10001011_00100100_10101111_0;
      patterns[35623] = 25'b10001011_00100101_10110000_0;
      patterns[35624] = 25'b10001011_00100110_10110001_0;
      patterns[35625] = 25'b10001011_00100111_10110010_0;
      patterns[35626] = 25'b10001011_00101000_10110011_0;
      patterns[35627] = 25'b10001011_00101001_10110100_0;
      patterns[35628] = 25'b10001011_00101010_10110101_0;
      patterns[35629] = 25'b10001011_00101011_10110110_0;
      patterns[35630] = 25'b10001011_00101100_10110111_0;
      patterns[35631] = 25'b10001011_00101101_10111000_0;
      patterns[35632] = 25'b10001011_00101110_10111001_0;
      patterns[35633] = 25'b10001011_00101111_10111010_0;
      patterns[35634] = 25'b10001011_00110000_10111011_0;
      patterns[35635] = 25'b10001011_00110001_10111100_0;
      patterns[35636] = 25'b10001011_00110010_10111101_0;
      patterns[35637] = 25'b10001011_00110011_10111110_0;
      patterns[35638] = 25'b10001011_00110100_10111111_0;
      patterns[35639] = 25'b10001011_00110101_11000000_0;
      patterns[35640] = 25'b10001011_00110110_11000001_0;
      patterns[35641] = 25'b10001011_00110111_11000010_0;
      patterns[35642] = 25'b10001011_00111000_11000011_0;
      patterns[35643] = 25'b10001011_00111001_11000100_0;
      patterns[35644] = 25'b10001011_00111010_11000101_0;
      patterns[35645] = 25'b10001011_00111011_11000110_0;
      patterns[35646] = 25'b10001011_00111100_11000111_0;
      patterns[35647] = 25'b10001011_00111101_11001000_0;
      patterns[35648] = 25'b10001011_00111110_11001001_0;
      patterns[35649] = 25'b10001011_00111111_11001010_0;
      patterns[35650] = 25'b10001011_01000000_11001011_0;
      patterns[35651] = 25'b10001011_01000001_11001100_0;
      patterns[35652] = 25'b10001011_01000010_11001101_0;
      patterns[35653] = 25'b10001011_01000011_11001110_0;
      patterns[35654] = 25'b10001011_01000100_11001111_0;
      patterns[35655] = 25'b10001011_01000101_11010000_0;
      patterns[35656] = 25'b10001011_01000110_11010001_0;
      patterns[35657] = 25'b10001011_01000111_11010010_0;
      patterns[35658] = 25'b10001011_01001000_11010011_0;
      patterns[35659] = 25'b10001011_01001001_11010100_0;
      patterns[35660] = 25'b10001011_01001010_11010101_0;
      patterns[35661] = 25'b10001011_01001011_11010110_0;
      patterns[35662] = 25'b10001011_01001100_11010111_0;
      patterns[35663] = 25'b10001011_01001101_11011000_0;
      patterns[35664] = 25'b10001011_01001110_11011001_0;
      patterns[35665] = 25'b10001011_01001111_11011010_0;
      patterns[35666] = 25'b10001011_01010000_11011011_0;
      patterns[35667] = 25'b10001011_01010001_11011100_0;
      patterns[35668] = 25'b10001011_01010010_11011101_0;
      patterns[35669] = 25'b10001011_01010011_11011110_0;
      patterns[35670] = 25'b10001011_01010100_11011111_0;
      patterns[35671] = 25'b10001011_01010101_11100000_0;
      patterns[35672] = 25'b10001011_01010110_11100001_0;
      patterns[35673] = 25'b10001011_01010111_11100010_0;
      patterns[35674] = 25'b10001011_01011000_11100011_0;
      patterns[35675] = 25'b10001011_01011001_11100100_0;
      patterns[35676] = 25'b10001011_01011010_11100101_0;
      patterns[35677] = 25'b10001011_01011011_11100110_0;
      patterns[35678] = 25'b10001011_01011100_11100111_0;
      patterns[35679] = 25'b10001011_01011101_11101000_0;
      patterns[35680] = 25'b10001011_01011110_11101001_0;
      patterns[35681] = 25'b10001011_01011111_11101010_0;
      patterns[35682] = 25'b10001011_01100000_11101011_0;
      patterns[35683] = 25'b10001011_01100001_11101100_0;
      patterns[35684] = 25'b10001011_01100010_11101101_0;
      patterns[35685] = 25'b10001011_01100011_11101110_0;
      patterns[35686] = 25'b10001011_01100100_11101111_0;
      patterns[35687] = 25'b10001011_01100101_11110000_0;
      patterns[35688] = 25'b10001011_01100110_11110001_0;
      patterns[35689] = 25'b10001011_01100111_11110010_0;
      patterns[35690] = 25'b10001011_01101000_11110011_0;
      patterns[35691] = 25'b10001011_01101001_11110100_0;
      patterns[35692] = 25'b10001011_01101010_11110101_0;
      patterns[35693] = 25'b10001011_01101011_11110110_0;
      patterns[35694] = 25'b10001011_01101100_11110111_0;
      patterns[35695] = 25'b10001011_01101101_11111000_0;
      patterns[35696] = 25'b10001011_01101110_11111001_0;
      patterns[35697] = 25'b10001011_01101111_11111010_0;
      patterns[35698] = 25'b10001011_01110000_11111011_0;
      patterns[35699] = 25'b10001011_01110001_11111100_0;
      patterns[35700] = 25'b10001011_01110010_11111101_0;
      patterns[35701] = 25'b10001011_01110011_11111110_0;
      patterns[35702] = 25'b10001011_01110100_11111111_0;
      patterns[35703] = 25'b10001011_01110101_00000000_1;
      patterns[35704] = 25'b10001011_01110110_00000001_1;
      patterns[35705] = 25'b10001011_01110111_00000010_1;
      patterns[35706] = 25'b10001011_01111000_00000011_1;
      patterns[35707] = 25'b10001011_01111001_00000100_1;
      patterns[35708] = 25'b10001011_01111010_00000101_1;
      patterns[35709] = 25'b10001011_01111011_00000110_1;
      patterns[35710] = 25'b10001011_01111100_00000111_1;
      patterns[35711] = 25'b10001011_01111101_00001000_1;
      patterns[35712] = 25'b10001011_01111110_00001001_1;
      patterns[35713] = 25'b10001011_01111111_00001010_1;
      patterns[35714] = 25'b10001011_10000000_00001011_1;
      patterns[35715] = 25'b10001011_10000001_00001100_1;
      patterns[35716] = 25'b10001011_10000010_00001101_1;
      patterns[35717] = 25'b10001011_10000011_00001110_1;
      patterns[35718] = 25'b10001011_10000100_00001111_1;
      patterns[35719] = 25'b10001011_10000101_00010000_1;
      patterns[35720] = 25'b10001011_10000110_00010001_1;
      patterns[35721] = 25'b10001011_10000111_00010010_1;
      patterns[35722] = 25'b10001011_10001000_00010011_1;
      patterns[35723] = 25'b10001011_10001001_00010100_1;
      patterns[35724] = 25'b10001011_10001010_00010101_1;
      patterns[35725] = 25'b10001011_10001011_00010110_1;
      patterns[35726] = 25'b10001011_10001100_00010111_1;
      patterns[35727] = 25'b10001011_10001101_00011000_1;
      patterns[35728] = 25'b10001011_10001110_00011001_1;
      patterns[35729] = 25'b10001011_10001111_00011010_1;
      patterns[35730] = 25'b10001011_10010000_00011011_1;
      patterns[35731] = 25'b10001011_10010001_00011100_1;
      patterns[35732] = 25'b10001011_10010010_00011101_1;
      patterns[35733] = 25'b10001011_10010011_00011110_1;
      patterns[35734] = 25'b10001011_10010100_00011111_1;
      patterns[35735] = 25'b10001011_10010101_00100000_1;
      patterns[35736] = 25'b10001011_10010110_00100001_1;
      patterns[35737] = 25'b10001011_10010111_00100010_1;
      patterns[35738] = 25'b10001011_10011000_00100011_1;
      patterns[35739] = 25'b10001011_10011001_00100100_1;
      patterns[35740] = 25'b10001011_10011010_00100101_1;
      patterns[35741] = 25'b10001011_10011011_00100110_1;
      patterns[35742] = 25'b10001011_10011100_00100111_1;
      patterns[35743] = 25'b10001011_10011101_00101000_1;
      patterns[35744] = 25'b10001011_10011110_00101001_1;
      patterns[35745] = 25'b10001011_10011111_00101010_1;
      patterns[35746] = 25'b10001011_10100000_00101011_1;
      patterns[35747] = 25'b10001011_10100001_00101100_1;
      patterns[35748] = 25'b10001011_10100010_00101101_1;
      patterns[35749] = 25'b10001011_10100011_00101110_1;
      patterns[35750] = 25'b10001011_10100100_00101111_1;
      patterns[35751] = 25'b10001011_10100101_00110000_1;
      patterns[35752] = 25'b10001011_10100110_00110001_1;
      patterns[35753] = 25'b10001011_10100111_00110010_1;
      patterns[35754] = 25'b10001011_10101000_00110011_1;
      patterns[35755] = 25'b10001011_10101001_00110100_1;
      patterns[35756] = 25'b10001011_10101010_00110101_1;
      patterns[35757] = 25'b10001011_10101011_00110110_1;
      patterns[35758] = 25'b10001011_10101100_00110111_1;
      patterns[35759] = 25'b10001011_10101101_00111000_1;
      patterns[35760] = 25'b10001011_10101110_00111001_1;
      patterns[35761] = 25'b10001011_10101111_00111010_1;
      patterns[35762] = 25'b10001011_10110000_00111011_1;
      patterns[35763] = 25'b10001011_10110001_00111100_1;
      patterns[35764] = 25'b10001011_10110010_00111101_1;
      patterns[35765] = 25'b10001011_10110011_00111110_1;
      patterns[35766] = 25'b10001011_10110100_00111111_1;
      patterns[35767] = 25'b10001011_10110101_01000000_1;
      patterns[35768] = 25'b10001011_10110110_01000001_1;
      patterns[35769] = 25'b10001011_10110111_01000010_1;
      patterns[35770] = 25'b10001011_10111000_01000011_1;
      patterns[35771] = 25'b10001011_10111001_01000100_1;
      patterns[35772] = 25'b10001011_10111010_01000101_1;
      patterns[35773] = 25'b10001011_10111011_01000110_1;
      patterns[35774] = 25'b10001011_10111100_01000111_1;
      patterns[35775] = 25'b10001011_10111101_01001000_1;
      patterns[35776] = 25'b10001011_10111110_01001001_1;
      patterns[35777] = 25'b10001011_10111111_01001010_1;
      patterns[35778] = 25'b10001011_11000000_01001011_1;
      patterns[35779] = 25'b10001011_11000001_01001100_1;
      patterns[35780] = 25'b10001011_11000010_01001101_1;
      patterns[35781] = 25'b10001011_11000011_01001110_1;
      patterns[35782] = 25'b10001011_11000100_01001111_1;
      patterns[35783] = 25'b10001011_11000101_01010000_1;
      patterns[35784] = 25'b10001011_11000110_01010001_1;
      patterns[35785] = 25'b10001011_11000111_01010010_1;
      patterns[35786] = 25'b10001011_11001000_01010011_1;
      patterns[35787] = 25'b10001011_11001001_01010100_1;
      patterns[35788] = 25'b10001011_11001010_01010101_1;
      patterns[35789] = 25'b10001011_11001011_01010110_1;
      patterns[35790] = 25'b10001011_11001100_01010111_1;
      patterns[35791] = 25'b10001011_11001101_01011000_1;
      patterns[35792] = 25'b10001011_11001110_01011001_1;
      patterns[35793] = 25'b10001011_11001111_01011010_1;
      patterns[35794] = 25'b10001011_11010000_01011011_1;
      patterns[35795] = 25'b10001011_11010001_01011100_1;
      patterns[35796] = 25'b10001011_11010010_01011101_1;
      patterns[35797] = 25'b10001011_11010011_01011110_1;
      patterns[35798] = 25'b10001011_11010100_01011111_1;
      patterns[35799] = 25'b10001011_11010101_01100000_1;
      patterns[35800] = 25'b10001011_11010110_01100001_1;
      patterns[35801] = 25'b10001011_11010111_01100010_1;
      patterns[35802] = 25'b10001011_11011000_01100011_1;
      patterns[35803] = 25'b10001011_11011001_01100100_1;
      patterns[35804] = 25'b10001011_11011010_01100101_1;
      patterns[35805] = 25'b10001011_11011011_01100110_1;
      patterns[35806] = 25'b10001011_11011100_01100111_1;
      patterns[35807] = 25'b10001011_11011101_01101000_1;
      patterns[35808] = 25'b10001011_11011110_01101001_1;
      patterns[35809] = 25'b10001011_11011111_01101010_1;
      patterns[35810] = 25'b10001011_11100000_01101011_1;
      patterns[35811] = 25'b10001011_11100001_01101100_1;
      patterns[35812] = 25'b10001011_11100010_01101101_1;
      patterns[35813] = 25'b10001011_11100011_01101110_1;
      patterns[35814] = 25'b10001011_11100100_01101111_1;
      patterns[35815] = 25'b10001011_11100101_01110000_1;
      patterns[35816] = 25'b10001011_11100110_01110001_1;
      patterns[35817] = 25'b10001011_11100111_01110010_1;
      patterns[35818] = 25'b10001011_11101000_01110011_1;
      patterns[35819] = 25'b10001011_11101001_01110100_1;
      patterns[35820] = 25'b10001011_11101010_01110101_1;
      patterns[35821] = 25'b10001011_11101011_01110110_1;
      patterns[35822] = 25'b10001011_11101100_01110111_1;
      patterns[35823] = 25'b10001011_11101101_01111000_1;
      patterns[35824] = 25'b10001011_11101110_01111001_1;
      patterns[35825] = 25'b10001011_11101111_01111010_1;
      patterns[35826] = 25'b10001011_11110000_01111011_1;
      patterns[35827] = 25'b10001011_11110001_01111100_1;
      patterns[35828] = 25'b10001011_11110010_01111101_1;
      patterns[35829] = 25'b10001011_11110011_01111110_1;
      patterns[35830] = 25'b10001011_11110100_01111111_1;
      patterns[35831] = 25'b10001011_11110101_10000000_1;
      patterns[35832] = 25'b10001011_11110110_10000001_1;
      patterns[35833] = 25'b10001011_11110111_10000010_1;
      patterns[35834] = 25'b10001011_11111000_10000011_1;
      patterns[35835] = 25'b10001011_11111001_10000100_1;
      patterns[35836] = 25'b10001011_11111010_10000101_1;
      patterns[35837] = 25'b10001011_11111011_10000110_1;
      patterns[35838] = 25'b10001011_11111100_10000111_1;
      patterns[35839] = 25'b10001011_11111101_10001000_1;
      patterns[35840] = 25'b10001011_11111110_10001001_1;
      patterns[35841] = 25'b10001011_11111111_10001010_1;
      patterns[35842] = 25'b10001100_00000000_10001100_0;
      patterns[35843] = 25'b10001100_00000001_10001101_0;
      patterns[35844] = 25'b10001100_00000010_10001110_0;
      patterns[35845] = 25'b10001100_00000011_10001111_0;
      patterns[35846] = 25'b10001100_00000100_10010000_0;
      patterns[35847] = 25'b10001100_00000101_10010001_0;
      patterns[35848] = 25'b10001100_00000110_10010010_0;
      patterns[35849] = 25'b10001100_00000111_10010011_0;
      patterns[35850] = 25'b10001100_00001000_10010100_0;
      patterns[35851] = 25'b10001100_00001001_10010101_0;
      patterns[35852] = 25'b10001100_00001010_10010110_0;
      patterns[35853] = 25'b10001100_00001011_10010111_0;
      patterns[35854] = 25'b10001100_00001100_10011000_0;
      patterns[35855] = 25'b10001100_00001101_10011001_0;
      patterns[35856] = 25'b10001100_00001110_10011010_0;
      patterns[35857] = 25'b10001100_00001111_10011011_0;
      patterns[35858] = 25'b10001100_00010000_10011100_0;
      patterns[35859] = 25'b10001100_00010001_10011101_0;
      patterns[35860] = 25'b10001100_00010010_10011110_0;
      patterns[35861] = 25'b10001100_00010011_10011111_0;
      patterns[35862] = 25'b10001100_00010100_10100000_0;
      patterns[35863] = 25'b10001100_00010101_10100001_0;
      patterns[35864] = 25'b10001100_00010110_10100010_0;
      patterns[35865] = 25'b10001100_00010111_10100011_0;
      patterns[35866] = 25'b10001100_00011000_10100100_0;
      patterns[35867] = 25'b10001100_00011001_10100101_0;
      patterns[35868] = 25'b10001100_00011010_10100110_0;
      patterns[35869] = 25'b10001100_00011011_10100111_0;
      patterns[35870] = 25'b10001100_00011100_10101000_0;
      patterns[35871] = 25'b10001100_00011101_10101001_0;
      patterns[35872] = 25'b10001100_00011110_10101010_0;
      patterns[35873] = 25'b10001100_00011111_10101011_0;
      patterns[35874] = 25'b10001100_00100000_10101100_0;
      patterns[35875] = 25'b10001100_00100001_10101101_0;
      patterns[35876] = 25'b10001100_00100010_10101110_0;
      patterns[35877] = 25'b10001100_00100011_10101111_0;
      patterns[35878] = 25'b10001100_00100100_10110000_0;
      patterns[35879] = 25'b10001100_00100101_10110001_0;
      patterns[35880] = 25'b10001100_00100110_10110010_0;
      patterns[35881] = 25'b10001100_00100111_10110011_0;
      patterns[35882] = 25'b10001100_00101000_10110100_0;
      patterns[35883] = 25'b10001100_00101001_10110101_0;
      patterns[35884] = 25'b10001100_00101010_10110110_0;
      patterns[35885] = 25'b10001100_00101011_10110111_0;
      patterns[35886] = 25'b10001100_00101100_10111000_0;
      patterns[35887] = 25'b10001100_00101101_10111001_0;
      patterns[35888] = 25'b10001100_00101110_10111010_0;
      patterns[35889] = 25'b10001100_00101111_10111011_0;
      patterns[35890] = 25'b10001100_00110000_10111100_0;
      patterns[35891] = 25'b10001100_00110001_10111101_0;
      patterns[35892] = 25'b10001100_00110010_10111110_0;
      patterns[35893] = 25'b10001100_00110011_10111111_0;
      patterns[35894] = 25'b10001100_00110100_11000000_0;
      patterns[35895] = 25'b10001100_00110101_11000001_0;
      patterns[35896] = 25'b10001100_00110110_11000010_0;
      patterns[35897] = 25'b10001100_00110111_11000011_0;
      patterns[35898] = 25'b10001100_00111000_11000100_0;
      patterns[35899] = 25'b10001100_00111001_11000101_0;
      patterns[35900] = 25'b10001100_00111010_11000110_0;
      patterns[35901] = 25'b10001100_00111011_11000111_0;
      patterns[35902] = 25'b10001100_00111100_11001000_0;
      patterns[35903] = 25'b10001100_00111101_11001001_0;
      patterns[35904] = 25'b10001100_00111110_11001010_0;
      patterns[35905] = 25'b10001100_00111111_11001011_0;
      patterns[35906] = 25'b10001100_01000000_11001100_0;
      patterns[35907] = 25'b10001100_01000001_11001101_0;
      patterns[35908] = 25'b10001100_01000010_11001110_0;
      patterns[35909] = 25'b10001100_01000011_11001111_0;
      patterns[35910] = 25'b10001100_01000100_11010000_0;
      patterns[35911] = 25'b10001100_01000101_11010001_0;
      patterns[35912] = 25'b10001100_01000110_11010010_0;
      patterns[35913] = 25'b10001100_01000111_11010011_0;
      patterns[35914] = 25'b10001100_01001000_11010100_0;
      patterns[35915] = 25'b10001100_01001001_11010101_0;
      patterns[35916] = 25'b10001100_01001010_11010110_0;
      patterns[35917] = 25'b10001100_01001011_11010111_0;
      patterns[35918] = 25'b10001100_01001100_11011000_0;
      patterns[35919] = 25'b10001100_01001101_11011001_0;
      patterns[35920] = 25'b10001100_01001110_11011010_0;
      patterns[35921] = 25'b10001100_01001111_11011011_0;
      patterns[35922] = 25'b10001100_01010000_11011100_0;
      patterns[35923] = 25'b10001100_01010001_11011101_0;
      patterns[35924] = 25'b10001100_01010010_11011110_0;
      patterns[35925] = 25'b10001100_01010011_11011111_0;
      patterns[35926] = 25'b10001100_01010100_11100000_0;
      patterns[35927] = 25'b10001100_01010101_11100001_0;
      patterns[35928] = 25'b10001100_01010110_11100010_0;
      patterns[35929] = 25'b10001100_01010111_11100011_0;
      patterns[35930] = 25'b10001100_01011000_11100100_0;
      patterns[35931] = 25'b10001100_01011001_11100101_0;
      patterns[35932] = 25'b10001100_01011010_11100110_0;
      patterns[35933] = 25'b10001100_01011011_11100111_0;
      patterns[35934] = 25'b10001100_01011100_11101000_0;
      patterns[35935] = 25'b10001100_01011101_11101001_0;
      patterns[35936] = 25'b10001100_01011110_11101010_0;
      patterns[35937] = 25'b10001100_01011111_11101011_0;
      patterns[35938] = 25'b10001100_01100000_11101100_0;
      patterns[35939] = 25'b10001100_01100001_11101101_0;
      patterns[35940] = 25'b10001100_01100010_11101110_0;
      patterns[35941] = 25'b10001100_01100011_11101111_0;
      patterns[35942] = 25'b10001100_01100100_11110000_0;
      patterns[35943] = 25'b10001100_01100101_11110001_0;
      patterns[35944] = 25'b10001100_01100110_11110010_0;
      patterns[35945] = 25'b10001100_01100111_11110011_0;
      patterns[35946] = 25'b10001100_01101000_11110100_0;
      patterns[35947] = 25'b10001100_01101001_11110101_0;
      patterns[35948] = 25'b10001100_01101010_11110110_0;
      patterns[35949] = 25'b10001100_01101011_11110111_0;
      patterns[35950] = 25'b10001100_01101100_11111000_0;
      patterns[35951] = 25'b10001100_01101101_11111001_0;
      patterns[35952] = 25'b10001100_01101110_11111010_0;
      patterns[35953] = 25'b10001100_01101111_11111011_0;
      patterns[35954] = 25'b10001100_01110000_11111100_0;
      patterns[35955] = 25'b10001100_01110001_11111101_0;
      patterns[35956] = 25'b10001100_01110010_11111110_0;
      patterns[35957] = 25'b10001100_01110011_11111111_0;
      patterns[35958] = 25'b10001100_01110100_00000000_1;
      patterns[35959] = 25'b10001100_01110101_00000001_1;
      patterns[35960] = 25'b10001100_01110110_00000010_1;
      patterns[35961] = 25'b10001100_01110111_00000011_1;
      patterns[35962] = 25'b10001100_01111000_00000100_1;
      patterns[35963] = 25'b10001100_01111001_00000101_1;
      patterns[35964] = 25'b10001100_01111010_00000110_1;
      patterns[35965] = 25'b10001100_01111011_00000111_1;
      patterns[35966] = 25'b10001100_01111100_00001000_1;
      patterns[35967] = 25'b10001100_01111101_00001001_1;
      patterns[35968] = 25'b10001100_01111110_00001010_1;
      patterns[35969] = 25'b10001100_01111111_00001011_1;
      patterns[35970] = 25'b10001100_10000000_00001100_1;
      patterns[35971] = 25'b10001100_10000001_00001101_1;
      patterns[35972] = 25'b10001100_10000010_00001110_1;
      patterns[35973] = 25'b10001100_10000011_00001111_1;
      patterns[35974] = 25'b10001100_10000100_00010000_1;
      patterns[35975] = 25'b10001100_10000101_00010001_1;
      patterns[35976] = 25'b10001100_10000110_00010010_1;
      patterns[35977] = 25'b10001100_10000111_00010011_1;
      patterns[35978] = 25'b10001100_10001000_00010100_1;
      patterns[35979] = 25'b10001100_10001001_00010101_1;
      patterns[35980] = 25'b10001100_10001010_00010110_1;
      patterns[35981] = 25'b10001100_10001011_00010111_1;
      patterns[35982] = 25'b10001100_10001100_00011000_1;
      patterns[35983] = 25'b10001100_10001101_00011001_1;
      patterns[35984] = 25'b10001100_10001110_00011010_1;
      patterns[35985] = 25'b10001100_10001111_00011011_1;
      patterns[35986] = 25'b10001100_10010000_00011100_1;
      patterns[35987] = 25'b10001100_10010001_00011101_1;
      patterns[35988] = 25'b10001100_10010010_00011110_1;
      patterns[35989] = 25'b10001100_10010011_00011111_1;
      patterns[35990] = 25'b10001100_10010100_00100000_1;
      patterns[35991] = 25'b10001100_10010101_00100001_1;
      patterns[35992] = 25'b10001100_10010110_00100010_1;
      patterns[35993] = 25'b10001100_10010111_00100011_1;
      patterns[35994] = 25'b10001100_10011000_00100100_1;
      patterns[35995] = 25'b10001100_10011001_00100101_1;
      patterns[35996] = 25'b10001100_10011010_00100110_1;
      patterns[35997] = 25'b10001100_10011011_00100111_1;
      patterns[35998] = 25'b10001100_10011100_00101000_1;
      patterns[35999] = 25'b10001100_10011101_00101001_1;
      patterns[36000] = 25'b10001100_10011110_00101010_1;
      patterns[36001] = 25'b10001100_10011111_00101011_1;
      patterns[36002] = 25'b10001100_10100000_00101100_1;
      patterns[36003] = 25'b10001100_10100001_00101101_1;
      patterns[36004] = 25'b10001100_10100010_00101110_1;
      patterns[36005] = 25'b10001100_10100011_00101111_1;
      patterns[36006] = 25'b10001100_10100100_00110000_1;
      patterns[36007] = 25'b10001100_10100101_00110001_1;
      patterns[36008] = 25'b10001100_10100110_00110010_1;
      patterns[36009] = 25'b10001100_10100111_00110011_1;
      patterns[36010] = 25'b10001100_10101000_00110100_1;
      patterns[36011] = 25'b10001100_10101001_00110101_1;
      patterns[36012] = 25'b10001100_10101010_00110110_1;
      patterns[36013] = 25'b10001100_10101011_00110111_1;
      patterns[36014] = 25'b10001100_10101100_00111000_1;
      patterns[36015] = 25'b10001100_10101101_00111001_1;
      patterns[36016] = 25'b10001100_10101110_00111010_1;
      patterns[36017] = 25'b10001100_10101111_00111011_1;
      patterns[36018] = 25'b10001100_10110000_00111100_1;
      patterns[36019] = 25'b10001100_10110001_00111101_1;
      patterns[36020] = 25'b10001100_10110010_00111110_1;
      patterns[36021] = 25'b10001100_10110011_00111111_1;
      patterns[36022] = 25'b10001100_10110100_01000000_1;
      patterns[36023] = 25'b10001100_10110101_01000001_1;
      patterns[36024] = 25'b10001100_10110110_01000010_1;
      patterns[36025] = 25'b10001100_10110111_01000011_1;
      patterns[36026] = 25'b10001100_10111000_01000100_1;
      patterns[36027] = 25'b10001100_10111001_01000101_1;
      patterns[36028] = 25'b10001100_10111010_01000110_1;
      patterns[36029] = 25'b10001100_10111011_01000111_1;
      patterns[36030] = 25'b10001100_10111100_01001000_1;
      patterns[36031] = 25'b10001100_10111101_01001001_1;
      patterns[36032] = 25'b10001100_10111110_01001010_1;
      patterns[36033] = 25'b10001100_10111111_01001011_1;
      patterns[36034] = 25'b10001100_11000000_01001100_1;
      patterns[36035] = 25'b10001100_11000001_01001101_1;
      patterns[36036] = 25'b10001100_11000010_01001110_1;
      patterns[36037] = 25'b10001100_11000011_01001111_1;
      patterns[36038] = 25'b10001100_11000100_01010000_1;
      patterns[36039] = 25'b10001100_11000101_01010001_1;
      patterns[36040] = 25'b10001100_11000110_01010010_1;
      patterns[36041] = 25'b10001100_11000111_01010011_1;
      patterns[36042] = 25'b10001100_11001000_01010100_1;
      patterns[36043] = 25'b10001100_11001001_01010101_1;
      patterns[36044] = 25'b10001100_11001010_01010110_1;
      patterns[36045] = 25'b10001100_11001011_01010111_1;
      patterns[36046] = 25'b10001100_11001100_01011000_1;
      patterns[36047] = 25'b10001100_11001101_01011001_1;
      patterns[36048] = 25'b10001100_11001110_01011010_1;
      patterns[36049] = 25'b10001100_11001111_01011011_1;
      patterns[36050] = 25'b10001100_11010000_01011100_1;
      patterns[36051] = 25'b10001100_11010001_01011101_1;
      patterns[36052] = 25'b10001100_11010010_01011110_1;
      patterns[36053] = 25'b10001100_11010011_01011111_1;
      patterns[36054] = 25'b10001100_11010100_01100000_1;
      patterns[36055] = 25'b10001100_11010101_01100001_1;
      patterns[36056] = 25'b10001100_11010110_01100010_1;
      patterns[36057] = 25'b10001100_11010111_01100011_1;
      patterns[36058] = 25'b10001100_11011000_01100100_1;
      patterns[36059] = 25'b10001100_11011001_01100101_1;
      patterns[36060] = 25'b10001100_11011010_01100110_1;
      patterns[36061] = 25'b10001100_11011011_01100111_1;
      patterns[36062] = 25'b10001100_11011100_01101000_1;
      patterns[36063] = 25'b10001100_11011101_01101001_1;
      patterns[36064] = 25'b10001100_11011110_01101010_1;
      patterns[36065] = 25'b10001100_11011111_01101011_1;
      patterns[36066] = 25'b10001100_11100000_01101100_1;
      patterns[36067] = 25'b10001100_11100001_01101101_1;
      patterns[36068] = 25'b10001100_11100010_01101110_1;
      patterns[36069] = 25'b10001100_11100011_01101111_1;
      patterns[36070] = 25'b10001100_11100100_01110000_1;
      patterns[36071] = 25'b10001100_11100101_01110001_1;
      patterns[36072] = 25'b10001100_11100110_01110010_1;
      patterns[36073] = 25'b10001100_11100111_01110011_1;
      patterns[36074] = 25'b10001100_11101000_01110100_1;
      patterns[36075] = 25'b10001100_11101001_01110101_1;
      patterns[36076] = 25'b10001100_11101010_01110110_1;
      patterns[36077] = 25'b10001100_11101011_01110111_1;
      patterns[36078] = 25'b10001100_11101100_01111000_1;
      patterns[36079] = 25'b10001100_11101101_01111001_1;
      patterns[36080] = 25'b10001100_11101110_01111010_1;
      patterns[36081] = 25'b10001100_11101111_01111011_1;
      patterns[36082] = 25'b10001100_11110000_01111100_1;
      patterns[36083] = 25'b10001100_11110001_01111101_1;
      patterns[36084] = 25'b10001100_11110010_01111110_1;
      patterns[36085] = 25'b10001100_11110011_01111111_1;
      patterns[36086] = 25'b10001100_11110100_10000000_1;
      patterns[36087] = 25'b10001100_11110101_10000001_1;
      patterns[36088] = 25'b10001100_11110110_10000010_1;
      patterns[36089] = 25'b10001100_11110111_10000011_1;
      patterns[36090] = 25'b10001100_11111000_10000100_1;
      patterns[36091] = 25'b10001100_11111001_10000101_1;
      patterns[36092] = 25'b10001100_11111010_10000110_1;
      patterns[36093] = 25'b10001100_11111011_10000111_1;
      patterns[36094] = 25'b10001100_11111100_10001000_1;
      patterns[36095] = 25'b10001100_11111101_10001001_1;
      patterns[36096] = 25'b10001100_11111110_10001010_1;
      patterns[36097] = 25'b10001100_11111111_10001011_1;
      patterns[36098] = 25'b10001101_00000000_10001101_0;
      patterns[36099] = 25'b10001101_00000001_10001110_0;
      patterns[36100] = 25'b10001101_00000010_10001111_0;
      patterns[36101] = 25'b10001101_00000011_10010000_0;
      patterns[36102] = 25'b10001101_00000100_10010001_0;
      patterns[36103] = 25'b10001101_00000101_10010010_0;
      patterns[36104] = 25'b10001101_00000110_10010011_0;
      patterns[36105] = 25'b10001101_00000111_10010100_0;
      patterns[36106] = 25'b10001101_00001000_10010101_0;
      patterns[36107] = 25'b10001101_00001001_10010110_0;
      patterns[36108] = 25'b10001101_00001010_10010111_0;
      patterns[36109] = 25'b10001101_00001011_10011000_0;
      patterns[36110] = 25'b10001101_00001100_10011001_0;
      patterns[36111] = 25'b10001101_00001101_10011010_0;
      patterns[36112] = 25'b10001101_00001110_10011011_0;
      patterns[36113] = 25'b10001101_00001111_10011100_0;
      patterns[36114] = 25'b10001101_00010000_10011101_0;
      patterns[36115] = 25'b10001101_00010001_10011110_0;
      patterns[36116] = 25'b10001101_00010010_10011111_0;
      patterns[36117] = 25'b10001101_00010011_10100000_0;
      patterns[36118] = 25'b10001101_00010100_10100001_0;
      patterns[36119] = 25'b10001101_00010101_10100010_0;
      patterns[36120] = 25'b10001101_00010110_10100011_0;
      patterns[36121] = 25'b10001101_00010111_10100100_0;
      patterns[36122] = 25'b10001101_00011000_10100101_0;
      patterns[36123] = 25'b10001101_00011001_10100110_0;
      patterns[36124] = 25'b10001101_00011010_10100111_0;
      patterns[36125] = 25'b10001101_00011011_10101000_0;
      patterns[36126] = 25'b10001101_00011100_10101001_0;
      patterns[36127] = 25'b10001101_00011101_10101010_0;
      patterns[36128] = 25'b10001101_00011110_10101011_0;
      patterns[36129] = 25'b10001101_00011111_10101100_0;
      patterns[36130] = 25'b10001101_00100000_10101101_0;
      patterns[36131] = 25'b10001101_00100001_10101110_0;
      patterns[36132] = 25'b10001101_00100010_10101111_0;
      patterns[36133] = 25'b10001101_00100011_10110000_0;
      patterns[36134] = 25'b10001101_00100100_10110001_0;
      patterns[36135] = 25'b10001101_00100101_10110010_0;
      patterns[36136] = 25'b10001101_00100110_10110011_0;
      patterns[36137] = 25'b10001101_00100111_10110100_0;
      patterns[36138] = 25'b10001101_00101000_10110101_0;
      patterns[36139] = 25'b10001101_00101001_10110110_0;
      patterns[36140] = 25'b10001101_00101010_10110111_0;
      patterns[36141] = 25'b10001101_00101011_10111000_0;
      patterns[36142] = 25'b10001101_00101100_10111001_0;
      patterns[36143] = 25'b10001101_00101101_10111010_0;
      patterns[36144] = 25'b10001101_00101110_10111011_0;
      patterns[36145] = 25'b10001101_00101111_10111100_0;
      patterns[36146] = 25'b10001101_00110000_10111101_0;
      patterns[36147] = 25'b10001101_00110001_10111110_0;
      patterns[36148] = 25'b10001101_00110010_10111111_0;
      patterns[36149] = 25'b10001101_00110011_11000000_0;
      patterns[36150] = 25'b10001101_00110100_11000001_0;
      patterns[36151] = 25'b10001101_00110101_11000010_0;
      patterns[36152] = 25'b10001101_00110110_11000011_0;
      patterns[36153] = 25'b10001101_00110111_11000100_0;
      patterns[36154] = 25'b10001101_00111000_11000101_0;
      patterns[36155] = 25'b10001101_00111001_11000110_0;
      patterns[36156] = 25'b10001101_00111010_11000111_0;
      patterns[36157] = 25'b10001101_00111011_11001000_0;
      patterns[36158] = 25'b10001101_00111100_11001001_0;
      patterns[36159] = 25'b10001101_00111101_11001010_0;
      patterns[36160] = 25'b10001101_00111110_11001011_0;
      patterns[36161] = 25'b10001101_00111111_11001100_0;
      patterns[36162] = 25'b10001101_01000000_11001101_0;
      patterns[36163] = 25'b10001101_01000001_11001110_0;
      patterns[36164] = 25'b10001101_01000010_11001111_0;
      patterns[36165] = 25'b10001101_01000011_11010000_0;
      patterns[36166] = 25'b10001101_01000100_11010001_0;
      patterns[36167] = 25'b10001101_01000101_11010010_0;
      patterns[36168] = 25'b10001101_01000110_11010011_0;
      patterns[36169] = 25'b10001101_01000111_11010100_0;
      patterns[36170] = 25'b10001101_01001000_11010101_0;
      patterns[36171] = 25'b10001101_01001001_11010110_0;
      patterns[36172] = 25'b10001101_01001010_11010111_0;
      patterns[36173] = 25'b10001101_01001011_11011000_0;
      patterns[36174] = 25'b10001101_01001100_11011001_0;
      patterns[36175] = 25'b10001101_01001101_11011010_0;
      patterns[36176] = 25'b10001101_01001110_11011011_0;
      patterns[36177] = 25'b10001101_01001111_11011100_0;
      patterns[36178] = 25'b10001101_01010000_11011101_0;
      patterns[36179] = 25'b10001101_01010001_11011110_0;
      patterns[36180] = 25'b10001101_01010010_11011111_0;
      patterns[36181] = 25'b10001101_01010011_11100000_0;
      patterns[36182] = 25'b10001101_01010100_11100001_0;
      patterns[36183] = 25'b10001101_01010101_11100010_0;
      patterns[36184] = 25'b10001101_01010110_11100011_0;
      patterns[36185] = 25'b10001101_01010111_11100100_0;
      patterns[36186] = 25'b10001101_01011000_11100101_0;
      patterns[36187] = 25'b10001101_01011001_11100110_0;
      patterns[36188] = 25'b10001101_01011010_11100111_0;
      patterns[36189] = 25'b10001101_01011011_11101000_0;
      patterns[36190] = 25'b10001101_01011100_11101001_0;
      patterns[36191] = 25'b10001101_01011101_11101010_0;
      patterns[36192] = 25'b10001101_01011110_11101011_0;
      patterns[36193] = 25'b10001101_01011111_11101100_0;
      patterns[36194] = 25'b10001101_01100000_11101101_0;
      patterns[36195] = 25'b10001101_01100001_11101110_0;
      patterns[36196] = 25'b10001101_01100010_11101111_0;
      patterns[36197] = 25'b10001101_01100011_11110000_0;
      patterns[36198] = 25'b10001101_01100100_11110001_0;
      patterns[36199] = 25'b10001101_01100101_11110010_0;
      patterns[36200] = 25'b10001101_01100110_11110011_0;
      patterns[36201] = 25'b10001101_01100111_11110100_0;
      patterns[36202] = 25'b10001101_01101000_11110101_0;
      patterns[36203] = 25'b10001101_01101001_11110110_0;
      patterns[36204] = 25'b10001101_01101010_11110111_0;
      patterns[36205] = 25'b10001101_01101011_11111000_0;
      patterns[36206] = 25'b10001101_01101100_11111001_0;
      patterns[36207] = 25'b10001101_01101101_11111010_0;
      patterns[36208] = 25'b10001101_01101110_11111011_0;
      patterns[36209] = 25'b10001101_01101111_11111100_0;
      patterns[36210] = 25'b10001101_01110000_11111101_0;
      patterns[36211] = 25'b10001101_01110001_11111110_0;
      patterns[36212] = 25'b10001101_01110010_11111111_0;
      patterns[36213] = 25'b10001101_01110011_00000000_1;
      patterns[36214] = 25'b10001101_01110100_00000001_1;
      patterns[36215] = 25'b10001101_01110101_00000010_1;
      patterns[36216] = 25'b10001101_01110110_00000011_1;
      patterns[36217] = 25'b10001101_01110111_00000100_1;
      patterns[36218] = 25'b10001101_01111000_00000101_1;
      patterns[36219] = 25'b10001101_01111001_00000110_1;
      patterns[36220] = 25'b10001101_01111010_00000111_1;
      patterns[36221] = 25'b10001101_01111011_00001000_1;
      patterns[36222] = 25'b10001101_01111100_00001001_1;
      patterns[36223] = 25'b10001101_01111101_00001010_1;
      patterns[36224] = 25'b10001101_01111110_00001011_1;
      patterns[36225] = 25'b10001101_01111111_00001100_1;
      patterns[36226] = 25'b10001101_10000000_00001101_1;
      patterns[36227] = 25'b10001101_10000001_00001110_1;
      patterns[36228] = 25'b10001101_10000010_00001111_1;
      patterns[36229] = 25'b10001101_10000011_00010000_1;
      patterns[36230] = 25'b10001101_10000100_00010001_1;
      patterns[36231] = 25'b10001101_10000101_00010010_1;
      patterns[36232] = 25'b10001101_10000110_00010011_1;
      patterns[36233] = 25'b10001101_10000111_00010100_1;
      patterns[36234] = 25'b10001101_10001000_00010101_1;
      patterns[36235] = 25'b10001101_10001001_00010110_1;
      patterns[36236] = 25'b10001101_10001010_00010111_1;
      patterns[36237] = 25'b10001101_10001011_00011000_1;
      patterns[36238] = 25'b10001101_10001100_00011001_1;
      patterns[36239] = 25'b10001101_10001101_00011010_1;
      patterns[36240] = 25'b10001101_10001110_00011011_1;
      patterns[36241] = 25'b10001101_10001111_00011100_1;
      patterns[36242] = 25'b10001101_10010000_00011101_1;
      patterns[36243] = 25'b10001101_10010001_00011110_1;
      patterns[36244] = 25'b10001101_10010010_00011111_1;
      patterns[36245] = 25'b10001101_10010011_00100000_1;
      patterns[36246] = 25'b10001101_10010100_00100001_1;
      patterns[36247] = 25'b10001101_10010101_00100010_1;
      patterns[36248] = 25'b10001101_10010110_00100011_1;
      patterns[36249] = 25'b10001101_10010111_00100100_1;
      patterns[36250] = 25'b10001101_10011000_00100101_1;
      patterns[36251] = 25'b10001101_10011001_00100110_1;
      patterns[36252] = 25'b10001101_10011010_00100111_1;
      patterns[36253] = 25'b10001101_10011011_00101000_1;
      patterns[36254] = 25'b10001101_10011100_00101001_1;
      patterns[36255] = 25'b10001101_10011101_00101010_1;
      patterns[36256] = 25'b10001101_10011110_00101011_1;
      patterns[36257] = 25'b10001101_10011111_00101100_1;
      patterns[36258] = 25'b10001101_10100000_00101101_1;
      patterns[36259] = 25'b10001101_10100001_00101110_1;
      patterns[36260] = 25'b10001101_10100010_00101111_1;
      patterns[36261] = 25'b10001101_10100011_00110000_1;
      patterns[36262] = 25'b10001101_10100100_00110001_1;
      patterns[36263] = 25'b10001101_10100101_00110010_1;
      patterns[36264] = 25'b10001101_10100110_00110011_1;
      patterns[36265] = 25'b10001101_10100111_00110100_1;
      patterns[36266] = 25'b10001101_10101000_00110101_1;
      patterns[36267] = 25'b10001101_10101001_00110110_1;
      patterns[36268] = 25'b10001101_10101010_00110111_1;
      patterns[36269] = 25'b10001101_10101011_00111000_1;
      patterns[36270] = 25'b10001101_10101100_00111001_1;
      patterns[36271] = 25'b10001101_10101101_00111010_1;
      patterns[36272] = 25'b10001101_10101110_00111011_1;
      patterns[36273] = 25'b10001101_10101111_00111100_1;
      patterns[36274] = 25'b10001101_10110000_00111101_1;
      patterns[36275] = 25'b10001101_10110001_00111110_1;
      patterns[36276] = 25'b10001101_10110010_00111111_1;
      patterns[36277] = 25'b10001101_10110011_01000000_1;
      patterns[36278] = 25'b10001101_10110100_01000001_1;
      patterns[36279] = 25'b10001101_10110101_01000010_1;
      patterns[36280] = 25'b10001101_10110110_01000011_1;
      patterns[36281] = 25'b10001101_10110111_01000100_1;
      patterns[36282] = 25'b10001101_10111000_01000101_1;
      patterns[36283] = 25'b10001101_10111001_01000110_1;
      patterns[36284] = 25'b10001101_10111010_01000111_1;
      patterns[36285] = 25'b10001101_10111011_01001000_1;
      patterns[36286] = 25'b10001101_10111100_01001001_1;
      patterns[36287] = 25'b10001101_10111101_01001010_1;
      patterns[36288] = 25'b10001101_10111110_01001011_1;
      patterns[36289] = 25'b10001101_10111111_01001100_1;
      patterns[36290] = 25'b10001101_11000000_01001101_1;
      patterns[36291] = 25'b10001101_11000001_01001110_1;
      patterns[36292] = 25'b10001101_11000010_01001111_1;
      patterns[36293] = 25'b10001101_11000011_01010000_1;
      patterns[36294] = 25'b10001101_11000100_01010001_1;
      patterns[36295] = 25'b10001101_11000101_01010010_1;
      patterns[36296] = 25'b10001101_11000110_01010011_1;
      patterns[36297] = 25'b10001101_11000111_01010100_1;
      patterns[36298] = 25'b10001101_11001000_01010101_1;
      patterns[36299] = 25'b10001101_11001001_01010110_1;
      patterns[36300] = 25'b10001101_11001010_01010111_1;
      patterns[36301] = 25'b10001101_11001011_01011000_1;
      patterns[36302] = 25'b10001101_11001100_01011001_1;
      patterns[36303] = 25'b10001101_11001101_01011010_1;
      patterns[36304] = 25'b10001101_11001110_01011011_1;
      patterns[36305] = 25'b10001101_11001111_01011100_1;
      patterns[36306] = 25'b10001101_11010000_01011101_1;
      patterns[36307] = 25'b10001101_11010001_01011110_1;
      patterns[36308] = 25'b10001101_11010010_01011111_1;
      patterns[36309] = 25'b10001101_11010011_01100000_1;
      patterns[36310] = 25'b10001101_11010100_01100001_1;
      patterns[36311] = 25'b10001101_11010101_01100010_1;
      patterns[36312] = 25'b10001101_11010110_01100011_1;
      patterns[36313] = 25'b10001101_11010111_01100100_1;
      patterns[36314] = 25'b10001101_11011000_01100101_1;
      patterns[36315] = 25'b10001101_11011001_01100110_1;
      patterns[36316] = 25'b10001101_11011010_01100111_1;
      patterns[36317] = 25'b10001101_11011011_01101000_1;
      patterns[36318] = 25'b10001101_11011100_01101001_1;
      patterns[36319] = 25'b10001101_11011101_01101010_1;
      patterns[36320] = 25'b10001101_11011110_01101011_1;
      patterns[36321] = 25'b10001101_11011111_01101100_1;
      patterns[36322] = 25'b10001101_11100000_01101101_1;
      patterns[36323] = 25'b10001101_11100001_01101110_1;
      patterns[36324] = 25'b10001101_11100010_01101111_1;
      patterns[36325] = 25'b10001101_11100011_01110000_1;
      patterns[36326] = 25'b10001101_11100100_01110001_1;
      patterns[36327] = 25'b10001101_11100101_01110010_1;
      patterns[36328] = 25'b10001101_11100110_01110011_1;
      patterns[36329] = 25'b10001101_11100111_01110100_1;
      patterns[36330] = 25'b10001101_11101000_01110101_1;
      patterns[36331] = 25'b10001101_11101001_01110110_1;
      patterns[36332] = 25'b10001101_11101010_01110111_1;
      patterns[36333] = 25'b10001101_11101011_01111000_1;
      patterns[36334] = 25'b10001101_11101100_01111001_1;
      patterns[36335] = 25'b10001101_11101101_01111010_1;
      patterns[36336] = 25'b10001101_11101110_01111011_1;
      patterns[36337] = 25'b10001101_11101111_01111100_1;
      patterns[36338] = 25'b10001101_11110000_01111101_1;
      patterns[36339] = 25'b10001101_11110001_01111110_1;
      patterns[36340] = 25'b10001101_11110010_01111111_1;
      patterns[36341] = 25'b10001101_11110011_10000000_1;
      patterns[36342] = 25'b10001101_11110100_10000001_1;
      patterns[36343] = 25'b10001101_11110101_10000010_1;
      patterns[36344] = 25'b10001101_11110110_10000011_1;
      patterns[36345] = 25'b10001101_11110111_10000100_1;
      patterns[36346] = 25'b10001101_11111000_10000101_1;
      patterns[36347] = 25'b10001101_11111001_10000110_1;
      patterns[36348] = 25'b10001101_11111010_10000111_1;
      patterns[36349] = 25'b10001101_11111011_10001000_1;
      patterns[36350] = 25'b10001101_11111100_10001001_1;
      patterns[36351] = 25'b10001101_11111101_10001010_1;
      patterns[36352] = 25'b10001101_11111110_10001011_1;
      patterns[36353] = 25'b10001101_11111111_10001100_1;
      patterns[36354] = 25'b10001110_00000000_10001110_0;
      patterns[36355] = 25'b10001110_00000001_10001111_0;
      patterns[36356] = 25'b10001110_00000010_10010000_0;
      patterns[36357] = 25'b10001110_00000011_10010001_0;
      patterns[36358] = 25'b10001110_00000100_10010010_0;
      patterns[36359] = 25'b10001110_00000101_10010011_0;
      patterns[36360] = 25'b10001110_00000110_10010100_0;
      patterns[36361] = 25'b10001110_00000111_10010101_0;
      patterns[36362] = 25'b10001110_00001000_10010110_0;
      patterns[36363] = 25'b10001110_00001001_10010111_0;
      patterns[36364] = 25'b10001110_00001010_10011000_0;
      patterns[36365] = 25'b10001110_00001011_10011001_0;
      patterns[36366] = 25'b10001110_00001100_10011010_0;
      patterns[36367] = 25'b10001110_00001101_10011011_0;
      patterns[36368] = 25'b10001110_00001110_10011100_0;
      patterns[36369] = 25'b10001110_00001111_10011101_0;
      patterns[36370] = 25'b10001110_00010000_10011110_0;
      patterns[36371] = 25'b10001110_00010001_10011111_0;
      patterns[36372] = 25'b10001110_00010010_10100000_0;
      patterns[36373] = 25'b10001110_00010011_10100001_0;
      patterns[36374] = 25'b10001110_00010100_10100010_0;
      patterns[36375] = 25'b10001110_00010101_10100011_0;
      patterns[36376] = 25'b10001110_00010110_10100100_0;
      patterns[36377] = 25'b10001110_00010111_10100101_0;
      patterns[36378] = 25'b10001110_00011000_10100110_0;
      patterns[36379] = 25'b10001110_00011001_10100111_0;
      patterns[36380] = 25'b10001110_00011010_10101000_0;
      patterns[36381] = 25'b10001110_00011011_10101001_0;
      patterns[36382] = 25'b10001110_00011100_10101010_0;
      patterns[36383] = 25'b10001110_00011101_10101011_0;
      patterns[36384] = 25'b10001110_00011110_10101100_0;
      patterns[36385] = 25'b10001110_00011111_10101101_0;
      patterns[36386] = 25'b10001110_00100000_10101110_0;
      patterns[36387] = 25'b10001110_00100001_10101111_0;
      patterns[36388] = 25'b10001110_00100010_10110000_0;
      patterns[36389] = 25'b10001110_00100011_10110001_0;
      patterns[36390] = 25'b10001110_00100100_10110010_0;
      patterns[36391] = 25'b10001110_00100101_10110011_0;
      patterns[36392] = 25'b10001110_00100110_10110100_0;
      patterns[36393] = 25'b10001110_00100111_10110101_0;
      patterns[36394] = 25'b10001110_00101000_10110110_0;
      patterns[36395] = 25'b10001110_00101001_10110111_0;
      patterns[36396] = 25'b10001110_00101010_10111000_0;
      patterns[36397] = 25'b10001110_00101011_10111001_0;
      patterns[36398] = 25'b10001110_00101100_10111010_0;
      patterns[36399] = 25'b10001110_00101101_10111011_0;
      patterns[36400] = 25'b10001110_00101110_10111100_0;
      patterns[36401] = 25'b10001110_00101111_10111101_0;
      patterns[36402] = 25'b10001110_00110000_10111110_0;
      patterns[36403] = 25'b10001110_00110001_10111111_0;
      patterns[36404] = 25'b10001110_00110010_11000000_0;
      patterns[36405] = 25'b10001110_00110011_11000001_0;
      patterns[36406] = 25'b10001110_00110100_11000010_0;
      patterns[36407] = 25'b10001110_00110101_11000011_0;
      patterns[36408] = 25'b10001110_00110110_11000100_0;
      patterns[36409] = 25'b10001110_00110111_11000101_0;
      patterns[36410] = 25'b10001110_00111000_11000110_0;
      patterns[36411] = 25'b10001110_00111001_11000111_0;
      patterns[36412] = 25'b10001110_00111010_11001000_0;
      patterns[36413] = 25'b10001110_00111011_11001001_0;
      patterns[36414] = 25'b10001110_00111100_11001010_0;
      patterns[36415] = 25'b10001110_00111101_11001011_0;
      patterns[36416] = 25'b10001110_00111110_11001100_0;
      patterns[36417] = 25'b10001110_00111111_11001101_0;
      patterns[36418] = 25'b10001110_01000000_11001110_0;
      patterns[36419] = 25'b10001110_01000001_11001111_0;
      patterns[36420] = 25'b10001110_01000010_11010000_0;
      patterns[36421] = 25'b10001110_01000011_11010001_0;
      patterns[36422] = 25'b10001110_01000100_11010010_0;
      patterns[36423] = 25'b10001110_01000101_11010011_0;
      patterns[36424] = 25'b10001110_01000110_11010100_0;
      patterns[36425] = 25'b10001110_01000111_11010101_0;
      patterns[36426] = 25'b10001110_01001000_11010110_0;
      patterns[36427] = 25'b10001110_01001001_11010111_0;
      patterns[36428] = 25'b10001110_01001010_11011000_0;
      patterns[36429] = 25'b10001110_01001011_11011001_0;
      patterns[36430] = 25'b10001110_01001100_11011010_0;
      patterns[36431] = 25'b10001110_01001101_11011011_0;
      patterns[36432] = 25'b10001110_01001110_11011100_0;
      patterns[36433] = 25'b10001110_01001111_11011101_0;
      patterns[36434] = 25'b10001110_01010000_11011110_0;
      patterns[36435] = 25'b10001110_01010001_11011111_0;
      patterns[36436] = 25'b10001110_01010010_11100000_0;
      patterns[36437] = 25'b10001110_01010011_11100001_0;
      patterns[36438] = 25'b10001110_01010100_11100010_0;
      patterns[36439] = 25'b10001110_01010101_11100011_0;
      patterns[36440] = 25'b10001110_01010110_11100100_0;
      patterns[36441] = 25'b10001110_01010111_11100101_0;
      patterns[36442] = 25'b10001110_01011000_11100110_0;
      patterns[36443] = 25'b10001110_01011001_11100111_0;
      patterns[36444] = 25'b10001110_01011010_11101000_0;
      patterns[36445] = 25'b10001110_01011011_11101001_0;
      patterns[36446] = 25'b10001110_01011100_11101010_0;
      patterns[36447] = 25'b10001110_01011101_11101011_0;
      patterns[36448] = 25'b10001110_01011110_11101100_0;
      patterns[36449] = 25'b10001110_01011111_11101101_0;
      patterns[36450] = 25'b10001110_01100000_11101110_0;
      patterns[36451] = 25'b10001110_01100001_11101111_0;
      patterns[36452] = 25'b10001110_01100010_11110000_0;
      patterns[36453] = 25'b10001110_01100011_11110001_0;
      patterns[36454] = 25'b10001110_01100100_11110010_0;
      patterns[36455] = 25'b10001110_01100101_11110011_0;
      patterns[36456] = 25'b10001110_01100110_11110100_0;
      patterns[36457] = 25'b10001110_01100111_11110101_0;
      patterns[36458] = 25'b10001110_01101000_11110110_0;
      patterns[36459] = 25'b10001110_01101001_11110111_0;
      patterns[36460] = 25'b10001110_01101010_11111000_0;
      patterns[36461] = 25'b10001110_01101011_11111001_0;
      patterns[36462] = 25'b10001110_01101100_11111010_0;
      patterns[36463] = 25'b10001110_01101101_11111011_0;
      patterns[36464] = 25'b10001110_01101110_11111100_0;
      patterns[36465] = 25'b10001110_01101111_11111101_0;
      patterns[36466] = 25'b10001110_01110000_11111110_0;
      patterns[36467] = 25'b10001110_01110001_11111111_0;
      patterns[36468] = 25'b10001110_01110010_00000000_1;
      patterns[36469] = 25'b10001110_01110011_00000001_1;
      patterns[36470] = 25'b10001110_01110100_00000010_1;
      patterns[36471] = 25'b10001110_01110101_00000011_1;
      patterns[36472] = 25'b10001110_01110110_00000100_1;
      patterns[36473] = 25'b10001110_01110111_00000101_1;
      patterns[36474] = 25'b10001110_01111000_00000110_1;
      patterns[36475] = 25'b10001110_01111001_00000111_1;
      patterns[36476] = 25'b10001110_01111010_00001000_1;
      patterns[36477] = 25'b10001110_01111011_00001001_1;
      patterns[36478] = 25'b10001110_01111100_00001010_1;
      patterns[36479] = 25'b10001110_01111101_00001011_1;
      patterns[36480] = 25'b10001110_01111110_00001100_1;
      patterns[36481] = 25'b10001110_01111111_00001101_1;
      patterns[36482] = 25'b10001110_10000000_00001110_1;
      patterns[36483] = 25'b10001110_10000001_00001111_1;
      patterns[36484] = 25'b10001110_10000010_00010000_1;
      patterns[36485] = 25'b10001110_10000011_00010001_1;
      patterns[36486] = 25'b10001110_10000100_00010010_1;
      patterns[36487] = 25'b10001110_10000101_00010011_1;
      patterns[36488] = 25'b10001110_10000110_00010100_1;
      patterns[36489] = 25'b10001110_10000111_00010101_1;
      patterns[36490] = 25'b10001110_10001000_00010110_1;
      patterns[36491] = 25'b10001110_10001001_00010111_1;
      patterns[36492] = 25'b10001110_10001010_00011000_1;
      patterns[36493] = 25'b10001110_10001011_00011001_1;
      patterns[36494] = 25'b10001110_10001100_00011010_1;
      patterns[36495] = 25'b10001110_10001101_00011011_1;
      patterns[36496] = 25'b10001110_10001110_00011100_1;
      patterns[36497] = 25'b10001110_10001111_00011101_1;
      patterns[36498] = 25'b10001110_10010000_00011110_1;
      patterns[36499] = 25'b10001110_10010001_00011111_1;
      patterns[36500] = 25'b10001110_10010010_00100000_1;
      patterns[36501] = 25'b10001110_10010011_00100001_1;
      patterns[36502] = 25'b10001110_10010100_00100010_1;
      patterns[36503] = 25'b10001110_10010101_00100011_1;
      patterns[36504] = 25'b10001110_10010110_00100100_1;
      patterns[36505] = 25'b10001110_10010111_00100101_1;
      patterns[36506] = 25'b10001110_10011000_00100110_1;
      patterns[36507] = 25'b10001110_10011001_00100111_1;
      patterns[36508] = 25'b10001110_10011010_00101000_1;
      patterns[36509] = 25'b10001110_10011011_00101001_1;
      patterns[36510] = 25'b10001110_10011100_00101010_1;
      patterns[36511] = 25'b10001110_10011101_00101011_1;
      patterns[36512] = 25'b10001110_10011110_00101100_1;
      patterns[36513] = 25'b10001110_10011111_00101101_1;
      patterns[36514] = 25'b10001110_10100000_00101110_1;
      patterns[36515] = 25'b10001110_10100001_00101111_1;
      patterns[36516] = 25'b10001110_10100010_00110000_1;
      patterns[36517] = 25'b10001110_10100011_00110001_1;
      patterns[36518] = 25'b10001110_10100100_00110010_1;
      patterns[36519] = 25'b10001110_10100101_00110011_1;
      patterns[36520] = 25'b10001110_10100110_00110100_1;
      patterns[36521] = 25'b10001110_10100111_00110101_1;
      patterns[36522] = 25'b10001110_10101000_00110110_1;
      patterns[36523] = 25'b10001110_10101001_00110111_1;
      patterns[36524] = 25'b10001110_10101010_00111000_1;
      patterns[36525] = 25'b10001110_10101011_00111001_1;
      patterns[36526] = 25'b10001110_10101100_00111010_1;
      patterns[36527] = 25'b10001110_10101101_00111011_1;
      patterns[36528] = 25'b10001110_10101110_00111100_1;
      patterns[36529] = 25'b10001110_10101111_00111101_1;
      patterns[36530] = 25'b10001110_10110000_00111110_1;
      patterns[36531] = 25'b10001110_10110001_00111111_1;
      patterns[36532] = 25'b10001110_10110010_01000000_1;
      patterns[36533] = 25'b10001110_10110011_01000001_1;
      patterns[36534] = 25'b10001110_10110100_01000010_1;
      patterns[36535] = 25'b10001110_10110101_01000011_1;
      patterns[36536] = 25'b10001110_10110110_01000100_1;
      patterns[36537] = 25'b10001110_10110111_01000101_1;
      patterns[36538] = 25'b10001110_10111000_01000110_1;
      patterns[36539] = 25'b10001110_10111001_01000111_1;
      patterns[36540] = 25'b10001110_10111010_01001000_1;
      patterns[36541] = 25'b10001110_10111011_01001001_1;
      patterns[36542] = 25'b10001110_10111100_01001010_1;
      patterns[36543] = 25'b10001110_10111101_01001011_1;
      patterns[36544] = 25'b10001110_10111110_01001100_1;
      patterns[36545] = 25'b10001110_10111111_01001101_1;
      patterns[36546] = 25'b10001110_11000000_01001110_1;
      patterns[36547] = 25'b10001110_11000001_01001111_1;
      patterns[36548] = 25'b10001110_11000010_01010000_1;
      patterns[36549] = 25'b10001110_11000011_01010001_1;
      patterns[36550] = 25'b10001110_11000100_01010010_1;
      patterns[36551] = 25'b10001110_11000101_01010011_1;
      patterns[36552] = 25'b10001110_11000110_01010100_1;
      patterns[36553] = 25'b10001110_11000111_01010101_1;
      patterns[36554] = 25'b10001110_11001000_01010110_1;
      patterns[36555] = 25'b10001110_11001001_01010111_1;
      patterns[36556] = 25'b10001110_11001010_01011000_1;
      patterns[36557] = 25'b10001110_11001011_01011001_1;
      patterns[36558] = 25'b10001110_11001100_01011010_1;
      patterns[36559] = 25'b10001110_11001101_01011011_1;
      patterns[36560] = 25'b10001110_11001110_01011100_1;
      patterns[36561] = 25'b10001110_11001111_01011101_1;
      patterns[36562] = 25'b10001110_11010000_01011110_1;
      patterns[36563] = 25'b10001110_11010001_01011111_1;
      patterns[36564] = 25'b10001110_11010010_01100000_1;
      patterns[36565] = 25'b10001110_11010011_01100001_1;
      patterns[36566] = 25'b10001110_11010100_01100010_1;
      patterns[36567] = 25'b10001110_11010101_01100011_1;
      patterns[36568] = 25'b10001110_11010110_01100100_1;
      patterns[36569] = 25'b10001110_11010111_01100101_1;
      patterns[36570] = 25'b10001110_11011000_01100110_1;
      patterns[36571] = 25'b10001110_11011001_01100111_1;
      patterns[36572] = 25'b10001110_11011010_01101000_1;
      patterns[36573] = 25'b10001110_11011011_01101001_1;
      patterns[36574] = 25'b10001110_11011100_01101010_1;
      patterns[36575] = 25'b10001110_11011101_01101011_1;
      patterns[36576] = 25'b10001110_11011110_01101100_1;
      patterns[36577] = 25'b10001110_11011111_01101101_1;
      patterns[36578] = 25'b10001110_11100000_01101110_1;
      patterns[36579] = 25'b10001110_11100001_01101111_1;
      patterns[36580] = 25'b10001110_11100010_01110000_1;
      patterns[36581] = 25'b10001110_11100011_01110001_1;
      patterns[36582] = 25'b10001110_11100100_01110010_1;
      patterns[36583] = 25'b10001110_11100101_01110011_1;
      patterns[36584] = 25'b10001110_11100110_01110100_1;
      patterns[36585] = 25'b10001110_11100111_01110101_1;
      patterns[36586] = 25'b10001110_11101000_01110110_1;
      patterns[36587] = 25'b10001110_11101001_01110111_1;
      patterns[36588] = 25'b10001110_11101010_01111000_1;
      patterns[36589] = 25'b10001110_11101011_01111001_1;
      patterns[36590] = 25'b10001110_11101100_01111010_1;
      patterns[36591] = 25'b10001110_11101101_01111011_1;
      patterns[36592] = 25'b10001110_11101110_01111100_1;
      patterns[36593] = 25'b10001110_11101111_01111101_1;
      patterns[36594] = 25'b10001110_11110000_01111110_1;
      patterns[36595] = 25'b10001110_11110001_01111111_1;
      patterns[36596] = 25'b10001110_11110010_10000000_1;
      patterns[36597] = 25'b10001110_11110011_10000001_1;
      patterns[36598] = 25'b10001110_11110100_10000010_1;
      patterns[36599] = 25'b10001110_11110101_10000011_1;
      patterns[36600] = 25'b10001110_11110110_10000100_1;
      patterns[36601] = 25'b10001110_11110111_10000101_1;
      patterns[36602] = 25'b10001110_11111000_10000110_1;
      patterns[36603] = 25'b10001110_11111001_10000111_1;
      patterns[36604] = 25'b10001110_11111010_10001000_1;
      patterns[36605] = 25'b10001110_11111011_10001001_1;
      patterns[36606] = 25'b10001110_11111100_10001010_1;
      patterns[36607] = 25'b10001110_11111101_10001011_1;
      patterns[36608] = 25'b10001110_11111110_10001100_1;
      patterns[36609] = 25'b10001110_11111111_10001101_1;
      patterns[36610] = 25'b10001111_00000000_10001111_0;
      patterns[36611] = 25'b10001111_00000001_10010000_0;
      patterns[36612] = 25'b10001111_00000010_10010001_0;
      patterns[36613] = 25'b10001111_00000011_10010010_0;
      patterns[36614] = 25'b10001111_00000100_10010011_0;
      patterns[36615] = 25'b10001111_00000101_10010100_0;
      patterns[36616] = 25'b10001111_00000110_10010101_0;
      patterns[36617] = 25'b10001111_00000111_10010110_0;
      patterns[36618] = 25'b10001111_00001000_10010111_0;
      patterns[36619] = 25'b10001111_00001001_10011000_0;
      patterns[36620] = 25'b10001111_00001010_10011001_0;
      patterns[36621] = 25'b10001111_00001011_10011010_0;
      patterns[36622] = 25'b10001111_00001100_10011011_0;
      patterns[36623] = 25'b10001111_00001101_10011100_0;
      patterns[36624] = 25'b10001111_00001110_10011101_0;
      patterns[36625] = 25'b10001111_00001111_10011110_0;
      patterns[36626] = 25'b10001111_00010000_10011111_0;
      patterns[36627] = 25'b10001111_00010001_10100000_0;
      patterns[36628] = 25'b10001111_00010010_10100001_0;
      patterns[36629] = 25'b10001111_00010011_10100010_0;
      patterns[36630] = 25'b10001111_00010100_10100011_0;
      patterns[36631] = 25'b10001111_00010101_10100100_0;
      patterns[36632] = 25'b10001111_00010110_10100101_0;
      patterns[36633] = 25'b10001111_00010111_10100110_0;
      patterns[36634] = 25'b10001111_00011000_10100111_0;
      patterns[36635] = 25'b10001111_00011001_10101000_0;
      patterns[36636] = 25'b10001111_00011010_10101001_0;
      patterns[36637] = 25'b10001111_00011011_10101010_0;
      patterns[36638] = 25'b10001111_00011100_10101011_0;
      patterns[36639] = 25'b10001111_00011101_10101100_0;
      patterns[36640] = 25'b10001111_00011110_10101101_0;
      patterns[36641] = 25'b10001111_00011111_10101110_0;
      patterns[36642] = 25'b10001111_00100000_10101111_0;
      patterns[36643] = 25'b10001111_00100001_10110000_0;
      patterns[36644] = 25'b10001111_00100010_10110001_0;
      patterns[36645] = 25'b10001111_00100011_10110010_0;
      patterns[36646] = 25'b10001111_00100100_10110011_0;
      patterns[36647] = 25'b10001111_00100101_10110100_0;
      patterns[36648] = 25'b10001111_00100110_10110101_0;
      patterns[36649] = 25'b10001111_00100111_10110110_0;
      patterns[36650] = 25'b10001111_00101000_10110111_0;
      patterns[36651] = 25'b10001111_00101001_10111000_0;
      patterns[36652] = 25'b10001111_00101010_10111001_0;
      patterns[36653] = 25'b10001111_00101011_10111010_0;
      patterns[36654] = 25'b10001111_00101100_10111011_0;
      patterns[36655] = 25'b10001111_00101101_10111100_0;
      patterns[36656] = 25'b10001111_00101110_10111101_0;
      patterns[36657] = 25'b10001111_00101111_10111110_0;
      patterns[36658] = 25'b10001111_00110000_10111111_0;
      patterns[36659] = 25'b10001111_00110001_11000000_0;
      patterns[36660] = 25'b10001111_00110010_11000001_0;
      patterns[36661] = 25'b10001111_00110011_11000010_0;
      patterns[36662] = 25'b10001111_00110100_11000011_0;
      patterns[36663] = 25'b10001111_00110101_11000100_0;
      patterns[36664] = 25'b10001111_00110110_11000101_0;
      patterns[36665] = 25'b10001111_00110111_11000110_0;
      patterns[36666] = 25'b10001111_00111000_11000111_0;
      patterns[36667] = 25'b10001111_00111001_11001000_0;
      patterns[36668] = 25'b10001111_00111010_11001001_0;
      patterns[36669] = 25'b10001111_00111011_11001010_0;
      patterns[36670] = 25'b10001111_00111100_11001011_0;
      patterns[36671] = 25'b10001111_00111101_11001100_0;
      patterns[36672] = 25'b10001111_00111110_11001101_0;
      patterns[36673] = 25'b10001111_00111111_11001110_0;
      patterns[36674] = 25'b10001111_01000000_11001111_0;
      patterns[36675] = 25'b10001111_01000001_11010000_0;
      patterns[36676] = 25'b10001111_01000010_11010001_0;
      patterns[36677] = 25'b10001111_01000011_11010010_0;
      patterns[36678] = 25'b10001111_01000100_11010011_0;
      patterns[36679] = 25'b10001111_01000101_11010100_0;
      patterns[36680] = 25'b10001111_01000110_11010101_0;
      patterns[36681] = 25'b10001111_01000111_11010110_0;
      patterns[36682] = 25'b10001111_01001000_11010111_0;
      patterns[36683] = 25'b10001111_01001001_11011000_0;
      patterns[36684] = 25'b10001111_01001010_11011001_0;
      patterns[36685] = 25'b10001111_01001011_11011010_0;
      patterns[36686] = 25'b10001111_01001100_11011011_0;
      patterns[36687] = 25'b10001111_01001101_11011100_0;
      patterns[36688] = 25'b10001111_01001110_11011101_0;
      patterns[36689] = 25'b10001111_01001111_11011110_0;
      patterns[36690] = 25'b10001111_01010000_11011111_0;
      patterns[36691] = 25'b10001111_01010001_11100000_0;
      patterns[36692] = 25'b10001111_01010010_11100001_0;
      patterns[36693] = 25'b10001111_01010011_11100010_0;
      patterns[36694] = 25'b10001111_01010100_11100011_0;
      patterns[36695] = 25'b10001111_01010101_11100100_0;
      patterns[36696] = 25'b10001111_01010110_11100101_0;
      patterns[36697] = 25'b10001111_01010111_11100110_0;
      patterns[36698] = 25'b10001111_01011000_11100111_0;
      patterns[36699] = 25'b10001111_01011001_11101000_0;
      patterns[36700] = 25'b10001111_01011010_11101001_0;
      patterns[36701] = 25'b10001111_01011011_11101010_0;
      patterns[36702] = 25'b10001111_01011100_11101011_0;
      patterns[36703] = 25'b10001111_01011101_11101100_0;
      patterns[36704] = 25'b10001111_01011110_11101101_0;
      patterns[36705] = 25'b10001111_01011111_11101110_0;
      patterns[36706] = 25'b10001111_01100000_11101111_0;
      patterns[36707] = 25'b10001111_01100001_11110000_0;
      patterns[36708] = 25'b10001111_01100010_11110001_0;
      patterns[36709] = 25'b10001111_01100011_11110010_0;
      patterns[36710] = 25'b10001111_01100100_11110011_0;
      patterns[36711] = 25'b10001111_01100101_11110100_0;
      patterns[36712] = 25'b10001111_01100110_11110101_0;
      patterns[36713] = 25'b10001111_01100111_11110110_0;
      patterns[36714] = 25'b10001111_01101000_11110111_0;
      patterns[36715] = 25'b10001111_01101001_11111000_0;
      patterns[36716] = 25'b10001111_01101010_11111001_0;
      patterns[36717] = 25'b10001111_01101011_11111010_0;
      patterns[36718] = 25'b10001111_01101100_11111011_0;
      patterns[36719] = 25'b10001111_01101101_11111100_0;
      patterns[36720] = 25'b10001111_01101110_11111101_0;
      patterns[36721] = 25'b10001111_01101111_11111110_0;
      patterns[36722] = 25'b10001111_01110000_11111111_0;
      patterns[36723] = 25'b10001111_01110001_00000000_1;
      patterns[36724] = 25'b10001111_01110010_00000001_1;
      patterns[36725] = 25'b10001111_01110011_00000010_1;
      patterns[36726] = 25'b10001111_01110100_00000011_1;
      patterns[36727] = 25'b10001111_01110101_00000100_1;
      patterns[36728] = 25'b10001111_01110110_00000101_1;
      patterns[36729] = 25'b10001111_01110111_00000110_1;
      patterns[36730] = 25'b10001111_01111000_00000111_1;
      patterns[36731] = 25'b10001111_01111001_00001000_1;
      patterns[36732] = 25'b10001111_01111010_00001001_1;
      patterns[36733] = 25'b10001111_01111011_00001010_1;
      patterns[36734] = 25'b10001111_01111100_00001011_1;
      patterns[36735] = 25'b10001111_01111101_00001100_1;
      patterns[36736] = 25'b10001111_01111110_00001101_1;
      patterns[36737] = 25'b10001111_01111111_00001110_1;
      patterns[36738] = 25'b10001111_10000000_00001111_1;
      patterns[36739] = 25'b10001111_10000001_00010000_1;
      patterns[36740] = 25'b10001111_10000010_00010001_1;
      patterns[36741] = 25'b10001111_10000011_00010010_1;
      patterns[36742] = 25'b10001111_10000100_00010011_1;
      patterns[36743] = 25'b10001111_10000101_00010100_1;
      patterns[36744] = 25'b10001111_10000110_00010101_1;
      patterns[36745] = 25'b10001111_10000111_00010110_1;
      patterns[36746] = 25'b10001111_10001000_00010111_1;
      patterns[36747] = 25'b10001111_10001001_00011000_1;
      patterns[36748] = 25'b10001111_10001010_00011001_1;
      patterns[36749] = 25'b10001111_10001011_00011010_1;
      patterns[36750] = 25'b10001111_10001100_00011011_1;
      patterns[36751] = 25'b10001111_10001101_00011100_1;
      patterns[36752] = 25'b10001111_10001110_00011101_1;
      patterns[36753] = 25'b10001111_10001111_00011110_1;
      patterns[36754] = 25'b10001111_10010000_00011111_1;
      patterns[36755] = 25'b10001111_10010001_00100000_1;
      patterns[36756] = 25'b10001111_10010010_00100001_1;
      patterns[36757] = 25'b10001111_10010011_00100010_1;
      patterns[36758] = 25'b10001111_10010100_00100011_1;
      patterns[36759] = 25'b10001111_10010101_00100100_1;
      patterns[36760] = 25'b10001111_10010110_00100101_1;
      patterns[36761] = 25'b10001111_10010111_00100110_1;
      patterns[36762] = 25'b10001111_10011000_00100111_1;
      patterns[36763] = 25'b10001111_10011001_00101000_1;
      patterns[36764] = 25'b10001111_10011010_00101001_1;
      patterns[36765] = 25'b10001111_10011011_00101010_1;
      patterns[36766] = 25'b10001111_10011100_00101011_1;
      patterns[36767] = 25'b10001111_10011101_00101100_1;
      patterns[36768] = 25'b10001111_10011110_00101101_1;
      patterns[36769] = 25'b10001111_10011111_00101110_1;
      patterns[36770] = 25'b10001111_10100000_00101111_1;
      patterns[36771] = 25'b10001111_10100001_00110000_1;
      patterns[36772] = 25'b10001111_10100010_00110001_1;
      patterns[36773] = 25'b10001111_10100011_00110010_1;
      patterns[36774] = 25'b10001111_10100100_00110011_1;
      patterns[36775] = 25'b10001111_10100101_00110100_1;
      patterns[36776] = 25'b10001111_10100110_00110101_1;
      patterns[36777] = 25'b10001111_10100111_00110110_1;
      patterns[36778] = 25'b10001111_10101000_00110111_1;
      patterns[36779] = 25'b10001111_10101001_00111000_1;
      patterns[36780] = 25'b10001111_10101010_00111001_1;
      patterns[36781] = 25'b10001111_10101011_00111010_1;
      patterns[36782] = 25'b10001111_10101100_00111011_1;
      patterns[36783] = 25'b10001111_10101101_00111100_1;
      patterns[36784] = 25'b10001111_10101110_00111101_1;
      patterns[36785] = 25'b10001111_10101111_00111110_1;
      patterns[36786] = 25'b10001111_10110000_00111111_1;
      patterns[36787] = 25'b10001111_10110001_01000000_1;
      patterns[36788] = 25'b10001111_10110010_01000001_1;
      patterns[36789] = 25'b10001111_10110011_01000010_1;
      patterns[36790] = 25'b10001111_10110100_01000011_1;
      patterns[36791] = 25'b10001111_10110101_01000100_1;
      patterns[36792] = 25'b10001111_10110110_01000101_1;
      patterns[36793] = 25'b10001111_10110111_01000110_1;
      patterns[36794] = 25'b10001111_10111000_01000111_1;
      patterns[36795] = 25'b10001111_10111001_01001000_1;
      patterns[36796] = 25'b10001111_10111010_01001001_1;
      patterns[36797] = 25'b10001111_10111011_01001010_1;
      patterns[36798] = 25'b10001111_10111100_01001011_1;
      patterns[36799] = 25'b10001111_10111101_01001100_1;
      patterns[36800] = 25'b10001111_10111110_01001101_1;
      patterns[36801] = 25'b10001111_10111111_01001110_1;
      patterns[36802] = 25'b10001111_11000000_01001111_1;
      patterns[36803] = 25'b10001111_11000001_01010000_1;
      patterns[36804] = 25'b10001111_11000010_01010001_1;
      patterns[36805] = 25'b10001111_11000011_01010010_1;
      patterns[36806] = 25'b10001111_11000100_01010011_1;
      patterns[36807] = 25'b10001111_11000101_01010100_1;
      patterns[36808] = 25'b10001111_11000110_01010101_1;
      patterns[36809] = 25'b10001111_11000111_01010110_1;
      patterns[36810] = 25'b10001111_11001000_01010111_1;
      patterns[36811] = 25'b10001111_11001001_01011000_1;
      patterns[36812] = 25'b10001111_11001010_01011001_1;
      patterns[36813] = 25'b10001111_11001011_01011010_1;
      patterns[36814] = 25'b10001111_11001100_01011011_1;
      patterns[36815] = 25'b10001111_11001101_01011100_1;
      patterns[36816] = 25'b10001111_11001110_01011101_1;
      patterns[36817] = 25'b10001111_11001111_01011110_1;
      patterns[36818] = 25'b10001111_11010000_01011111_1;
      patterns[36819] = 25'b10001111_11010001_01100000_1;
      patterns[36820] = 25'b10001111_11010010_01100001_1;
      patterns[36821] = 25'b10001111_11010011_01100010_1;
      patterns[36822] = 25'b10001111_11010100_01100011_1;
      patterns[36823] = 25'b10001111_11010101_01100100_1;
      patterns[36824] = 25'b10001111_11010110_01100101_1;
      patterns[36825] = 25'b10001111_11010111_01100110_1;
      patterns[36826] = 25'b10001111_11011000_01100111_1;
      patterns[36827] = 25'b10001111_11011001_01101000_1;
      patterns[36828] = 25'b10001111_11011010_01101001_1;
      patterns[36829] = 25'b10001111_11011011_01101010_1;
      patterns[36830] = 25'b10001111_11011100_01101011_1;
      patterns[36831] = 25'b10001111_11011101_01101100_1;
      patterns[36832] = 25'b10001111_11011110_01101101_1;
      patterns[36833] = 25'b10001111_11011111_01101110_1;
      patterns[36834] = 25'b10001111_11100000_01101111_1;
      patterns[36835] = 25'b10001111_11100001_01110000_1;
      patterns[36836] = 25'b10001111_11100010_01110001_1;
      patterns[36837] = 25'b10001111_11100011_01110010_1;
      patterns[36838] = 25'b10001111_11100100_01110011_1;
      patterns[36839] = 25'b10001111_11100101_01110100_1;
      patterns[36840] = 25'b10001111_11100110_01110101_1;
      patterns[36841] = 25'b10001111_11100111_01110110_1;
      patterns[36842] = 25'b10001111_11101000_01110111_1;
      patterns[36843] = 25'b10001111_11101001_01111000_1;
      patterns[36844] = 25'b10001111_11101010_01111001_1;
      patterns[36845] = 25'b10001111_11101011_01111010_1;
      patterns[36846] = 25'b10001111_11101100_01111011_1;
      patterns[36847] = 25'b10001111_11101101_01111100_1;
      patterns[36848] = 25'b10001111_11101110_01111101_1;
      patterns[36849] = 25'b10001111_11101111_01111110_1;
      patterns[36850] = 25'b10001111_11110000_01111111_1;
      patterns[36851] = 25'b10001111_11110001_10000000_1;
      patterns[36852] = 25'b10001111_11110010_10000001_1;
      patterns[36853] = 25'b10001111_11110011_10000010_1;
      patterns[36854] = 25'b10001111_11110100_10000011_1;
      patterns[36855] = 25'b10001111_11110101_10000100_1;
      patterns[36856] = 25'b10001111_11110110_10000101_1;
      patterns[36857] = 25'b10001111_11110111_10000110_1;
      patterns[36858] = 25'b10001111_11111000_10000111_1;
      patterns[36859] = 25'b10001111_11111001_10001000_1;
      patterns[36860] = 25'b10001111_11111010_10001001_1;
      patterns[36861] = 25'b10001111_11111011_10001010_1;
      patterns[36862] = 25'b10001111_11111100_10001011_1;
      patterns[36863] = 25'b10001111_11111101_10001100_1;
      patterns[36864] = 25'b10001111_11111110_10001101_1;
      patterns[36865] = 25'b10001111_11111111_10001110_1;
      patterns[36866] = 25'b10010000_00000000_10010000_0;
      patterns[36867] = 25'b10010000_00000001_10010001_0;
      patterns[36868] = 25'b10010000_00000010_10010010_0;
      patterns[36869] = 25'b10010000_00000011_10010011_0;
      patterns[36870] = 25'b10010000_00000100_10010100_0;
      patterns[36871] = 25'b10010000_00000101_10010101_0;
      patterns[36872] = 25'b10010000_00000110_10010110_0;
      patterns[36873] = 25'b10010000_00000111_10010111_0;
      patterns[36874] = 25'b10010000_00001000_10011000_0;
      patterns[36875] = 25'b10010000_00001001_10011001_0;
      patterns[36876] = 25'b10010000_00001010_10011010_0;
      patterns[36877] = 25'b10010000_00001011_10011011_0;
      patterns[36878] = 25'b10010000_00001100_10011100_0;
      patterns[36879] = 25'b10010000_00001101_10011101_0;
      patterns[36880] = 25'b10010000_00001110_10011110_0;
      patterns[36881] = 25'b10010000_00001111_10011111_0;
      patterns[36882] = 25'b10010000_00010000_10100000_0;
      patterns[36883] = 25'b10010000_00010001_10100001_0;
      patterns[36884] = 25'b10010000_00010010_10100010_0;
      patterns[36885] = 25'b10010000_00010011_10100011_0;
      patterns[36886] = 25'b10010000_00010100_10100100_0;
      patterns[36887] = 25'b10010000_00010101_10100101_0;
      patterns[36888] = 25'b10010000_00010110_10100110_0;
      patterns[36889] = 25'b10010000_00010111_10100111_0;
      patterns[36890] = 25'b10010000_00011000_10101000_0;
      patterns[36891] = 25'b10010000_00011001_10101001_0;
      patterns[36892] = 25'b10010000_00011010_10101010_0;
      patterns[36893] = 25'b10010000_00011011_10101011_0;
      patterns[36894] = 25'b10010000_00011100_10101100_0;
      patterns[36895] = 25'b10010000_00011101_10101101_0;
      patterns[36896] = 25'b10010000_00011110_10101110_0;
      patterns[36897] = 25'b10010000_00011111_10101111_0;
      patterns[36898] = 25'b10010000_00100000_10110000_0;
      patterns[36899] = 25'b10010000_00100001_10110001_0;
      patterns[36900] = 25'b10010000_00100010_10110010_0;
      patterns[36901] = 25'b10010000_00100011_10110011_0;
      patterns[36902] = 25'b10010000_00100100_10110100_0;
      patterns[36903] = 25'b10010000_00100101_10110101_0;
      patterns[36904] = 25'b10010000_00100110_10110110_0;
      patterns[36905] = 25'b10010000_00100111_10110111_0;
      patterns[36906] = 25'b10010000_00101000_10111000_0;
      patterns[36907] = 25'b10010000_00101001_10111001_0;
      patterns[36908] = 25'b10010000_00101010_10111010_0;
      patterns[36909] = 25'b10010000_00101011_10111011_0;
      patterns[36910] = 25'b10010000_00101100_10111100_0;
      patterns[36911] = 25'b10010000_00101101_10111101_0;
      patterns[36912] = 25'b10010000_00101110_10111110_0;
      patterns[36913] = 25'b10010000_00101111_10111111_0;
      patterns[36914] = 25'b10010000_00110000_11000000_0;
      patterns[36915] = 25'b10010000_00110001_11000001_0;
      patterns[36916] = 25'b10010000_00110010_11000010_0;
      patterns[36917] = 25'b10010000_00110011_11000011_0;
      patterns[36918] = 25'b10010000_00110100_11000100_0;
      patterns[36919] = 25'b10010000_00110101_11000101_0;
      patterns[36920] = 25'b10010000_00110110_11000110_0;
      patterns[36921] = 25'b10010000_00110111_11000111_0;
      patterns[36922] = 25'b10010000_00111000_11001000_0;
      patterns[36923] = 25'b10010000_00111001_11001001_0;
      patterns[36924] = 25'b10010000_00111010_11001010_0;
      patterns[36925] = 25'b10010000_00111011_11001011_0;
      patterns[36926] = 25'b10010000_00111100_11001100_0;
      patterns[36927] = 25'b10010000_00111101_11001101_0;
      patterns[36928] = 25'b10010000_00111110_11001110_0;
      patterns[36929] = 25'b10010000_00111111_11001111_0;
      patterns[36930] = 25'b10010000_01000000_11010000_0;
      patterns[36931] = 25'b10010000_01000001_11010001_0;
      patterns[36932] = 25'b10010000_01000010_11010010_0;
      patterns[36933] = 25'b10010000_01000011_11010011_0;
      patterns[36934] = 25'b10010000_01000100_11010100_0;
      patterns[36935] = 25'b10010000_01000101_11010101_0;
      patterns[36936] = 25'b10010000_01000110_11010110_0;
      patterns[36937] = 25'b10010000_01000111_11010111_0;
      patterns[36938] = 25'b10010000_01001000_11011000_0;
      patterns[36939] = 25'b10010000_01001001_11011001_0;
      patterns[36940] = 25'b10010000_01001010_11011010_0;
      patterns[36941] = 25'b10010000_01001011_11011011_0;
      patterns[36942] = 25'b10010000_01001100_11011100_0;
      patterns[36943] = 25'b10010000_01001101_11011101_0;
      patterns[36944] = 25'b10010000_01001110_11011110_0;
      patterns[36945] = 25'b10010000_01001111_11011111_0;
      patterns[36946] = 25'b10010000_01010000_11100000_0;
      patterns[36947] = 25'b10010000_01010001_11100001_0;
      patterns[36948] = 25'b10010000_01010010_11100010_0;
      patterns[36949] = 25'b10010000_01010011_11100011_0;
      patterns[36950] = 25'b10010000_01010100_11100100_0;
      patterns[36951] = 25'b10010000_01010101_11100101_0;
      patterns[36952] = 25'b10010000_01010110_11100110_0;
      patterns[36953] = 25'b10010000_01010111_11100111_0;
      patterns[36954] = 25'b10010000_01011000_11101000_0;
      patterns[36955] = 25'b10010000_01011001_11101001_0;
      patterns[36956] = 25'b10010000_01011010_11101010_0;
      patterns[36957] = 25'b10010000_01011011_11101011_0;
      patterns[36958] = 25'b10010000_01011100_11101100_0;
      patterns[36959] = 25'b10010000_01011101_11101101_0;
      patterns[36960] = 25'b10010000_01011110_11101110_0;
      patterns[36961] = 25'b10010000_01011111_11101111_0;
      patterns[36962] = 25'b10010000_01100000_11110000_0;
      patterns[36963] = 25'b10010000_01100001_11110001_0;
      patterns[36964] = 25'b10010000_01100010_11110010_0;
      patterns[36965] = 25'b10010000_01100011_11110011_0;
      patterns[36966] = 25'b10010000_01100100_11110100_0;
      patterns[36967] = 25'b10010000_01100101_11110101_0;
      patterns[36968] = 25'b10010000_01100110_11110110_0;
      patterns[36969] = 25'b10010000_01100111_11110111_0;
      patterns[36970] = 25'b10010000_01101000_11111000_0;
      patterns[36971] = 25'b10010000_01101001_11111001_0;
      patterns[36972] = 25'b10010000_01101010_11111010_0;
      patterns[36973] = 25'b10010000_01101011_11111011_0;
      patterns[36974] = 25'b10010000_01101100_11111100_0;
      patterns[36975] = 25'b10010000_01101101_11111101_0;
      patterns[36976] = 25'b10010000_01101110_11111110_0;
      patterns[36977] = 25'b10010000_01101111_11111111_0;
      patterns[36978] = 25'b10010000_01110000_00000000_1;
      patterns[36979] = 25'b10010000_01110001_00000001_1;
      patterns[36980] = 25'b10010000_01110010_00000010_1;
      patterns[36981] = 25'b10010000_01110011_00000011_1;
      patterns[36982] = 25'b10010000_01110100_00000100_1;
      patterns[36983] = 25'b10010000_01110101_00000101_1;
      patterns[36984] = 25'b10010000_01110110_00000110_1;
      patterns[36985] = 25'b10010000_01110111_00000111_1;
      patterns[36986] = 25'b10010000_01111000_00001000_1;
      patterns[36987] = 25'b10010000_01111001_00001001_1;
      patterns[36988] = 25'b10010000_01111010_00001010_1;
      patterns[36989] = 25'b10010000_01111011_00001011_1;
      patterns[36990] = 25'b10010000_01111100_00001100_1;
      patterns[36991] = 25'b10010000_01111101_00001101_1;
      patterns[36992] = 25'b10010000_01111110_00001110_1;
      patterns[36993] = 25'b10010000_01111111_00001111_1;
      patterns[36994] = 25'b10010000_10000000_00010000_1;
      patterns[36995] = 25'b10010000_10000001_00010001_1;
      patterns[36996] = 25'b10010000_10000010_00010010_1;
      patterns[36997] = 25'b10010000_10000011_00010011_1;
      patterns[36998] = 25'b10010000_10000100_00010100_1;
      patterns[36999] = 25'b10010000_10000101_00010101_1;
      patterns[37000] = 25'b10010000_10000110_00010110_1;
      patterns[37001] = 25'b10010000_10000111_00010111_1;
      patterns[37002] = 25'b10010000_10001000_00011000_1;
      patterns[37003] = 25'b10010000_10001001_00011001_1;
      patterns[37004] = 25'b10010000_10001010_00011010_1;
      patterns[37005] = 25'b10010000_10001011_00011011_1;
      patterns[37006] = 25'b10010000_10001100_00011100_1;
      patterns[37007] = 25'b10010000_10001101_00011101_1;
      patterns[37008] = 25'b10010000_10001110_00011110_1;
      patterns[37009] = 25'b10010000_10001111_00011111_1;
      patterns[37010] = 25'b10010000_10010000_00100000_1;
      patterns[37011] = 25'b10010000_10010001_00100001_1;
      patterns[37012] = 25'b10010000_10010010_00100010_1;
      patterns[37013] = 25'b10010000_10010011_00100011_1;
      patterns[37014] = 25'b10010000_10010100_00100100_1;
      patterns[37015] = 25'b10010000_10010101_00100101_1;
      patterns[37016] = 25'b10010000_10010110_00100110_1;
      patterns[37017] = 25'b10010000_10010111_00100111_1;
      patterns[37018] = 25'b10010000_10011000_00101000_1;
      patterns[37019] = 25'b10010000_10011001_00101001_1;
      patterns[37020] = 25'b10010000_10011010_00101010_1;
      patterns[37021] = 25'b10010000_10011011_00101011_1;
      patterns[37022] = 25'b10010000_10011100_00101100_1;
      patterns[37023] = 25'b10010000_10011101_00101101_1;
      patterns[37024] = 25'b10010000_10011110_00101110_1;
      patterns[37025] = 25'b10010000_10011111_00101111_1;
      patterns[37026] = 25'b10010000_10100000_00110000_1;
      patterns[37027] = 25'b10010000_10100001_00110001_1;
      patterns[37028] = 25'b10010000_10100010_00110010_1;
      patterns[37029] = 25'b10010000_10100011_00110011_1;
      patterns[37030] = 25'b10010000_10100100_00110100_1;
      patterns[37031] = 25'b10010000_10100101_00110101_1;
      patterns[37032] = 25'b10010000_10100110_00110110_1;
      patterns[37033] = 25'b10010000_10100111_00110111_1;
      patterns[37034] = 25'b10010000_10101000_00111000_1;
      patterns[37035] = 25'b10010000_10101001_00111001_1;
      patterns[37036] = 25'b10010000_10101010_00111010_1;
      patterns[37037] = 25'b10010000_10101011_00111011_1;
      patterns[37038] = 25'b10010000_10101100_00111100_1;
      patterns[37039] = 25'b10010000_10101101_00111101_1;
      patterns[37040] = 25'b10010000_10101110_00111110_1;
      patterns[37041] = 25'b10010000_10101111_00111111_1;
      patterns[37042] = 25'b10010000_10110000_01000000_1;
      patterns[37043] = 25'b10010000_10110001_01000001_1;
      patterns[37044] = 25'b10010000_10110010_01000010_1;
      patterns[37045] = 25'b10010000_10110011_01000011_1;
      patterns[37046] = 25'b10010000_10110100_01000100_1;
      patterns[37047] = 25'b10010000_10110101_01000101_1;
      patterns[37048] = 25'b10010000_10110110_01000110_1;
      patterns[37049] = 25'b10010000_10110111_01000111_1;
      patterns[37050] = 25'b10010000_10111000_01001000_1;
      patterns[37051] = 25'b10010000_10111001_01001001_1;
      patterns[37052] = 25'b10010000_10111010_01001010_1;
      patterns[37053] = 25'b10010000_10111011_01001011_1;
      patterns[37054] = 25'b10010000_10111100_01001100_1;
      patterns[37055] = 25'b10010000_10111101_01001101_1;
      patterns[37056] = 25'b10010000_10111110_01001110_1;
      patterns[37057] = 25'b10010000_10111111_01001111_1;
      patterns[37058] = 25'b10010000_11000000_01010000_1;
      patterns[37059] = 25'b10010000_11000001_01010001_1;
      patterns[37060] = 25'b10010000_11000010_01010010_1;
      patterns[37061] = 25'b10010000_11000011_01010011_1;
      patterns[37062] = 25'b10010000_11000100_01010100_1;
      patterns[37063] = 25'b10010000_11000101_01010101_1;
      patterns[37064] = 25'b10010000_11000110_01010110_1;
      patterns[37065] = 25'b10010000_11000111_01010111_1;
      patterns[37066] = 25'b10010000_11001000_01011000_1;
      patterns[37067] = 25'b10010000_11001001_01011001_1;
      patterns[37068] = 25'b10010000_11001010_01011010_1;
      patterns[37069] = 25'b10010000_11001011_01011011_1;
      patterns[37070] = 25'b10010000_11001100_01011100_1;
      patterns[37071] = 25'b10010000_11001101_01011101_1;
      patterns[37072] = 25'b10010000_11001110_01011110_1;
      patterns[37073] = 25'b10010000_11001111_01011111_1;
      patterns[37074] = 25'b10010000_11010000_01100000_1;
      patterns[37075] = 25'b10010000_11010001_01100001_1;
      patterns[37076] = 25'b10010000_11010010_01100010_1;
      patterns[37077] = 25'b10010000_11010011_01100011_1;
      patterns[37078] = 25'b10010000_11010100_01100100_1;
      patterns[37079] = 25'b10010000_11010101_01100101_1;
      patterns[37080] = 25'b10010000_11010110_01100110_1;
      patterns[37081] = 25'b10010000_11010111_01100111_1;
      patterns[37082] = 25'b10010000_11011000_01101000_1;
      patterns[37083] = 25'b10010000_11011001_01101001_1;
      patterns[37084] = 25'b10010000_11011010_01101010_1;
      patterns[37085] = 25'b10010000_11011011_01101011_1;
      patterns[37086] = 25'b10010000_11011100_01101100_1;
      patterns[37087] = 25'b10010000_11011101_01101101_1;
      patterns[37088] = 25'b10010000_11011110_01101110_1;
      patterns[37089] = 25'b10010000_11011111_01101111_1;
      patterns[37090] = 25'b10010000_11100000_01110000_1;
      patterns[37091] = 25'b10010000_11100001_01110001_1;
      patterns[37092] = 25'b10010000_11100010_01110010_1;
      patterns[37093] = 25'b10010000_11100011_01110011_1;
      patterns[37094] = 25'b10010000_11100100_01110100_1;
      patterns[37095] = 25'b10010000_11100101_01110101_1;
      patterns[37096] = 25'b10010000_11100110_01110110_1;
      patterns[37097] = 25'b10010000_11100111_01110111_1;
      patterns[37098] = 25'b10010000_11101000_01111000_1;
      patterns[37099] = 25'b10010000_11101001_01111001_1;
      patterns[37100] = 25'b10010000_11101010_01111010_1;
      patterns[37101] = 25'b10010000_11101011_01111011_1;
      patterns[37102] = 25'b10010000_11101100_01111100_1;
      patterns[37103] = 25'b10010000_11101101_01111101_1;
      patterns[37104] = 25'b10010000_11101110_01111110_1;
      patterns[37105] = 25'b10010000_11101111_01111111_1;
      patterns[37106] = 25'b10010000_11110000_10000000_1;
      patterns[37107] = 25'b10010000_11110001_10000001_1;
      patterns[37108] = 25'b10010000_11110010_10000010_1;
      patterns[37109] = 25'b10010000_11110011_10000011_1;
      patterns[37110] = 25'b10010000_11110100_10000100_1;
      patterns[37111] = 25'b10010000_11110101_10000101_1;
      patterns[37112] = 25'b10010000_11110110_10000110_1;
      patterns[37113] = 25'b10010000_11110111_10000111_1;
      patterns[37114] = 25'b10010000_11111000_10001000_1;
      patterns[37115] = 25'b10010000_11111001_10001001_1;
      patterns[37116] = 25'b10010000_11111010_10001010_1;
      patterns[37117] = 25'b10010000_11111011_10001011_1;
      patterns[37118] = 25'b10010000_11111100_10001100_1;
      patterns[37119] = 25'b10010000_11111101_10001101_1;
      patterns[37120] = 25'b10010000_11111110_10001110_1;
      patterns[37121] = 25'b10010000_11111111_10001111_1;
      patterns[37122] = 25'b10010001_00000000_10010001_0;
      patterns[37123] = 25'b10010001_00000001_10010010_0;
      patterns[37124] = 25'b10010001_00000010_10010011_0;
      patterns[37125] = 25'b10010001_00000011_10010100_0;
      patterns[37126] = 25'b10010001_00000100_10010101_0;
      patterns[37127] = 25'b10010001_00000101_10010110_0;
      patterns[37128] = 25'b10010001_00000110_10010111_0;
      patterns[37129] = 25'b10010001_00000111_10011000_0;
      patterns[37130] = 25'b10010001_00001000_10011001_0;
      patterns[37131] = 25'b10010001_00001001_10011010_0;
      patterns[37132] = 25'b10010001_00001010_10011011_0;
      patterns[37133] = 25'b10010001_00001011_10011100_0;
      patterns[37134] = 25'b10010001_00001100_10011101_0;
      patterns[37135] = 25'b10010001_00001101_10011110_0;
      patterns[37136] = 25'b10010001_00001110_10011111_0;
      patterns[37137] = 25'b10010001_00001111_10100000_0;
      patterns[37138] = 25'b10010001_00010000_10100001_0;
      patterns[37139] = 25'b10010001_00010001_10100010_0;
      patterns[37140] = 25'b10010001_00010010_10100011_0;
      patterns[37141] = 25'b10010001_00010011_10100100_0;
      patterns[37142] = 25'b10010001_00010100_10100101_0;
      patterns[37143] = 25'b10010001_00010101_10100110_0;
      patterns[37144] = 25'b10010001_00010110_10100111_0;
      patterns[37145] = 25'b10010001_00010111_10101000_0;
      patterns[37146] = 25'b10010001_00011000_10101001_0;
      patterns[37147] = 25'b10010001_00011001_10101010_0;
      patterns[37148] = 25'b10010001_00011010_10101011_0;
      patterns[37149] = 25'b10010001_00011011_10101100_0;
      patterns[37150] = 25'b10010001_00011100_10101101_0;
      patterns[37151] = 25'b10010001_00011101_10101110_0;
      patterns[37152] = 25'b10010001_00011110_10101111_0;
      patterns[37153] = 25'b10010001_00011111_10110000_0;
      patterns[37154] = 25'b10010001_00100000_10110001_0;
      patterns[37155] = 25'b10010001_00100001_10110010_0;
      patterns[37156] = 25'b10010001_00100010_10110011_0;
      patterns[37157] = 25'b10010001_00100011_10110100_0;
      patterns[37158] = 25'b10010001_00100100_10110101_0;
      patterns[37159] = 25'b10010001_00100101_10110110_0;
      patterns[37160] = 25'b10010001_00100110_10110111_0;
      patterns[37161] = 25'b10010001_00100111_10111000_0;
      patterns[37162] = 25'b10010001_00101000_10111001_0;
      patterns[37163] = 25'b10010001_00101001_10111010_0;
      patterns[37164] = 25'b10010001_00101010_10111011_0;
      patterns[37165] = 25'b10010001_00101011_10111100_0;
      patterns[37166] = 25'b10010001_00101100_10111101_0;
      patterns[37167] = 25'b10010001_00101101_10111110_0;
      patterns[37168] = 25'b10010001_00101110_10111111_0;
      patterns[37169] = 25'b10010001_00101111_11000000_0;
      patterns[37170] = 25'b10010001_00110000_11000001_0;
      patterns[37171] = 25'b10010001_00110001_11000010_0;
      patterns[37172] = 25'b10010001_00110010_11000011_0;
      patterns[37173] = 25'b10010001_00110011_11000100_0;
      patterns[37174] = 25'b10010001_00110100_11000101_0;
      patterns[37175] = 25'b10010001_00110101_11000110_0;
      patterns[37176] = 25'b10010001_00110110_11000111_0;
      patterns[37177] = 25'b10010001_00110111_11001000_0;
      patterns[37178] = 25'b10010001_00111000_11001001_0;
      patterns[37179] = 25'b10010001_00111001_11001010_0;
      patterns[37180] = 25'b10010001_00111010_11001011_0;
      patterns[37181] = 25'b10010001_00111011_11001100_0;
      patterns[37182] = 25'b10010001_00111100_11001101_0;
      patterns[37183] = 25'b10010001_00111101_11001110_0;
      patterns[37184] = 25'b10010001_00111110_11001111_0;
      patterns[37185] = 25'b10010001_00111111_11010000_0;
      patterns[37186] = 25'b10010001_01000000_11010001_0;
      patterns[37187] = 25'b10010001_01000001_11010010_0;
      patterns[37188] = 25'b10010001_01000010_11010011_0;
      patterns[37189] = 25'b10010001_01000011_11010100_0;
      patterns[37190] = 25'b10010001_01000100_11010101_0;
      patterns[37191] = 25'b10010001_01000101_11010110_0;
      patterns[37192] = 25'b10010001_01000110_11010111_0;
      patterns[37193] = 25'b10010001_01000111_11011000_0;
      patterns[37194] = 25'b10010001_01001000_11011001_0;
      patterns[37195] = 25'b10010001_01001001_11011010_0;
      patterns[37196] = 25'b10010001_01001010_11011011_0;
      patterns[37197] = 25'b10010001_01001011_11011100_0;
      patterns[37198] = 25'b10010001_01001100_11011101_0;
      patterns[37199] = 25'b10010001_01001101_11011110_0;
      patterns[37200] = 25'b10010001_01001110_11011111_0;
      patterns[37201] = 25'b10010001_01001111_11100000_0;
      patterns[37202] = 25'b10010001_01010000_11100001_0;
      patterns[37203] = 25'b10010001_01010001_11100010_0;
      patterns[37204] = 25'b10010001_01010010_11100011_0;
      patterns[37205] = 25'b10010001_01010011_11100100_0;
      patterns[37206] = 25'b10010001_01010100_11100101_0;
      patterns[37207] = 25'b10010001_01010101_11100110_0;
      patterns[37208] = 25'b10010001_01010110_11100111_0;
      patterns[37209] = 25'b10010001_01010111_11101000_0;
      patterns[37210] = 25'b10010001_01011000_11101001_0;
      patterns[37211] = 25'b10010001_01011001_11101010_0;
      patterns[37212] = 25'b10010001_01011010_11101011_0;
      patterns[37213] = 25'b10010001_01011011_11101100_0;
      patterns[37214] = 25'b10010001_01011100_11101101_0;
      patterns[37215] = 25'b10010001_01011101_11101110_0;
      patterns[37216] = 25'b10010001_01011110_11101111_0;
      patterns[37217] = 25'b10010001_01011111_11110000_0;
      patterns[37218] = 25'b10010001_01100000_11110001_0;
      patterns[37219] = 25'b10010001_01100001_11110010_0;
      patterns[37220] = 25'b10010001_01100010_11110011_0;
      patterns[37221] = 25'b10010001_01100011_11110100_0;
      patterns[37222] = 25'b10010001_01100100_11110101_0;
      patterns[37223] = 25'b10010001_01100101_11110110_0;
      patterns[37224] = 25'b10010001_01100110_11110111_0;
      patterns[37225] = 25'b10010001_01100111_11111000_0;
      patterns[37226] = 25'b10010001_01101000_11111001_0;
      patterns[37227] = 25'b10010001_01101001_11111010_0;
      patterns[37228] = 25'b10010001_01101010_11111011_0;
      patterns[37229] = 25'b10010001_01101011_11111100_0;
      patterns[37230] = 25'b10010001_01101100_11111101_0;
      patterns[37231] = 25'b10010001_01101101_11111110_0;
      patterns[37232] = 25'b10010001_01101110_11111111_0;
      patterns[37233] = 25'b10010001_01101111_00000000_1;
      patterns[37234] = 25'b10010001_01110000_00000001_1;
      patterns[37235] = 25'b10010001_01110001_00000010_1;
      patterns[37236] = 25'b10010001_01110010_00000011_1;
      patterns[37237] = 25'b10010001_01110011_00000100_1;
      patterns[37238] = 25'b10010001_01110100_00000101_1;
      patterns[37239] = 25'b10010001_01110101_00000110_1;
      patterns[37240] = 25'b10010001_01110110_00000111_1;
      patterns[37241] = 25'b10010001_01110111_00001000_1;
      patterns[37242] = 25'b10010001_01111000_00001001_1;
      patterns[37243] = 25'b10010001_01111001_00001010_1;
      patterns[37244] = 25'b10010001_01111010_00001011_1;
      patterns[37245] = 25'b10010001_01111011_00001100_1;
      patterns[37246] = 25'b10010001_01111100_00001101_1;
      patterns[37247] = 25'b10010001_01111101_00001110_1;
      patterns[37248] = 25'b10010001_01111110_00001111_1;
      patterns[37249] = 25'b10010001_01111111_00010000_1;
      patterns[37250] = 25'b10010001_10000000_00010001_1;
      patterns[37251] = 25'b10010001_10000001_00010010_1;
      patterns[37252] = 25'b10010001_10000010_00010011_1;
      patterns[37253] = 25'b10010001_10000011_00010100_1;
      patterns[37254] = 25'b10010001_10000100_00010101_1;
      patterns[37255] = 25'b10010001_10000101_00010110_1;
      patterns[37256] = 25'b10010001_10000110_00010111_1;
      patterns[37257] = 25'b10010001_10000111_00011000_1;
      patterns[37258] = 25'b10010001_10001000_00011001_1;
      patterns[37259] = 25'b10010001_10001001_00011010_1;
      patterns[37260] = 25'b10010001_10001010_00011011_1;
      patterns[37261] = 25'b10010001_10001011_00011100_1;
      patterns[37262] = 25'b10010001_10001100_00011101_1;
      patterns[37263] = 25'b10010001_10001101_00011110_1;
      patterns[37264] = 25'b10010001_10001110_00011111_1;
      patterns[37265] = 25'b10010001_10001111_00100000_1;
      patterns[37266] = 25'b10010001_10010000_00100001_1;
      patterns[37267] = 25'b10010001_10010001_00100010_1;
      patterns[37268] = 25'b10010001_10010010_00100011_1;
      patterns[37269] = 25'b10010001_10010011_00100100_1;
      patterns[37270] = 25'b10010001_10010100_00100101_1;
      patterns[37271] = 25'b10010001_10010101_00100110_1;
      patterns[37272] = 25'b10010001_10010110_00100111_1;
      patterns[37273] = 25'b10010001_10010111_00101000_1;
      patterns[37274] = 25'b10010001_10011000_00101001_1;
      patterns[37275] = 25'b10010001_10011001_00101010_1;
      patterns[37276] = 25'b10010001_10011010_00101011_1;
      patterns[37277] = 25'b10010001_10011011_00101100_1;
      patterns[37278] = 25'b10010001_10011100_00101101_1;
      patterns[37279] = 25'b10010001_10011101_00101110_1;
      patterns[37280] = 25'b10010001_10011110_00101111_1;
      patterns[37281] = 25'b10010001_10011111_00110000_1;
      patterns[37282] = 25'b10010001_10100000_00110001_1;
      patterns[37283] = 25'b10010001_10100001_00110010_1;
      patterns[37284] = 25'b10010001_10100010_00110011_1;
      patterns[37285] = 25'b10010001_10100011_00110100_1;
      patterns[37286] = 25'b10010001_10100100_00110101_1;
      patterns[37287] = 25'b10010001_10100101_00110110_1;
      patterns[37288] = 25'b10010001_10100110_00110111_1;
      patterns[37289] = 25'b10010001_10100111_00111000_1;
      patterns[37290] = 25'b10010001_10101000_00111001_1;
      patterns[37291] = 25'b10010001_10101001_00111010_1;
      patterns[37292] = 25'b10010001_10101010_00111011_1;
      patterns[37293] = 25'b10010001_10101011_00111100_1;
      patterns[37294] = 25'b10010001_10101100_00111101_1;
      patterns[37295] = 25'b10010001_10101101_00111110_1;
      patterns[37296] = 25'b10010001_10101110_00111111_1;
      patterns[37297] = 25'b10010001_10101111_01000000_1;
      patterns[37298] = 25'b10010001_10110000_01000001_1;
      patterns[37299] = 25'b10010001_10110001_01000010_1;
      patterns[37300] = 25'b10010001_10110010_01000011_1;
      patterns[37301] = 25'b10010001_10110011_01000100_1;
      patterns[37302] = 25'b10010001_10110100_01000101_1;
      patterns[37303] = 25'b10010001_10110101_01000110_1;
      patterns[37304] = 25'b10010001_10110110_01000111_1;
      patterns[37305] = 25'b10010001_10110111_01001000_1;
      patterns[37306] = 25'b10010001_10111000_01001001_1;
      patterns[37307] = 25'b10010001_10111001_01001010_1;
      patterns[37308] = 25'b10010001_10111010_01001011_1;
      patterns[37309] = 25'b10010001_10111011_01001100_1;
      patterns[37310] = 25'b10010001_10111100_01001101_1;
      patterns[37311] = 25'b10010001_10111101_01001110_1;
      patterns[37312] = 25'b10010001_10111110_01001111_1;
      patterns[37313] = 25'b10010001_10111111_01010000_1;
      patterns[37314] = 25'b10010001_11000000_01010001_1;
      patterns[37315] = 25'b10010001_11000001_01010010_1;
      patterns[37316] = 25'b10010001_11000010_01010011_1;
      patterns[37317] = 25'b10010001_11000011_01010100_1;
      patterns[37318] = 25'b10010001_11000100_01010101_1;
      patterns[37319] = 25'b10010001_11000101_01010110_1;
      patterns[37320] = 25'b10010001_11000110_01010111_1;
      patterns[37321] = 25'b10010001_11000111_01011000_1;
      patterns[37322] = 25'b10010001_11001000_01011001_1;
      patterns[37323] = 25'b10010001_11001001_01011010_1;
      patterns[37324] = 25'b10010001_11001010_01011011_1;
      patterns[37325] = 25'b10010001_11001011_01011100_1;
      patterns[37326] = 25'b10010001_11001100_01011101_1;
      patterns[37327] = 25'b10010001_11001101_01011110_1;
      patterns[37328] = 25'b10010001_11001110_01011111_1;
      patterns[37329] = 25'b10010001_11001111_01100000_1;
      patterns[37330] = 25'b10010001_11010000_01100001_1;
      patterns[37331] = 25'b10010001_11010001_01100010_1;
      patterns[37332] = 25'b10010001_11010010_01100011_1;
      patterns[37333] = 25'b10010001_11010011_01100100_1;
      patterns[37334] = 25'b10010001_11010100_01100101_1;
      patterns[37335] = 25'b10010001_11010101_01100110_1;
      patterns[37336] = 25'b10010001_11010110_01100111_1;
      patterns[37337] = 25'b10010001_11010111_01101000_1;
      patterns[37338] = 25'b10010001_11011000_01101001_1;
      patterns[37339] = 25'b10010001_11011001_01101010_1;
      patterns[37340] = 25'b10010001_11011010_01101011_1;
      patterns[37341] = 25'b10010001_11011011_01101100_1;
      patterns[37342] = 25'b10010001_11011100_01101101_1;
      patterns[37343] = 25'b10010001_11011101_01101110_1;
      patterns[37344] = 25'b10010001_11011110_01101111_1;
      patterns[37345] = 25'b10010001_11011111_01110000_1;
      patterns[37346] = 25'b10010001_11100000_01110001_1;
      patterns[37347] = 25'b10010001_11100001_01110010_1;
      patterns[37348] = 25'b10010001_11100010_01110011_1;
      patterns[37349] = 25'b10010001_11100011_01110100_1;
      patterns[37350] = 25'b10010001_11100100_01110101_1;
      patterns[37351] = 25'b10010001_11100101_01110110_1;
      patterns[37352] = 25'b10010001_11100110_01110111_1;
      patterns[37353] = 25'b10010001_11100111_01111000_1;
      patterns[37354] = 25'b10010001_11101000_01111001_1;
      patterns[37355] = 25'b10010001_11101001_01111010_1;
      patterns[37356] = 25'b10010001_11101010_01111011_1;
      patterns[37357] = 25'b10010001_11101011_01111100_1;
      patterns[37358] = 25'b10010001_11101100_01111101_1;
      patterns[37359] = 25'b10010001_11101101_01111110_1;
      patterns[37360] = 25'b10010001_11101110_01111111_1;
      patterns[37361] = 25'b10010001_11101111_10000000_1;
      patterns[37362] = 25'b10010001_11110000_10000001_1;
      patterns[37363] = 25'b10010001_11110001_10000010_1;
      patterns[37364] = 25'b10010001_11110010_10000011_1;
      patterns[37365] = 25'b10010001_11110011_10000100_1;
      patterns[37366] = 25'b10010001_11110100_10000101_1;
      patterns[37367] = 25'b10010001_11110101_10000110_1;
      patterns[37368] = 25'b10010001_11110110_10000111_1;
      patterns[37369] = 25'b10010001_11110111_10001000_1;
      patterns[37370] = 25'b10010001_11111000_10001001_1;
      patterns[37371] = 25'b10010001_11111001_10001010_1;
      patterns[37372] = 25'b10010001_11111010_10001011_1;
      patterns[37373] = 25'b10010001_11111011_10001100_1;
      patterns[37374] = 25'b10010001_11111100_10001101_1;
      patterns[37375] = 25'b10010001_11111101_10001110_1;
      patterns[37376] = 25'b10010001_11111110_10001111_1;
      patterns[37377] = 25'b10010001_11111111_10010000_1;
      patterns[37378] = 25'b10010010_00000000_10010010_0;
      patterns[37379] = 25'b10010010_00000001_10010011_0;
      patterns[37380] = 25'b10010010_00000010_10010100_0;
      patterns[37381] = 25'b10010010_00000011_10010101_0;
      patterns[37382] = 25'b10010010_00000100_10010110_0;
      patterns[37383] = 25'b10010010_00000101_10010111_0;
      patterns[37384] = 25'b10010010_00000110_10011000_0;
      patterns[37385] = 25'b10010010_00000111_10011001_0;
      patterns[37386] = 25'b10010010_00001000_10011010_0;
      patterns[37387] = 25'b10010010_00001001_10011011_0;
      patterns[37388] = 25'b10010010_00001010_10011100_0;
      patterns[37389] = 25'b10010010_00001011_10011101_0;
      patterns[37390] = 25'b10010010_00001100_10011110_0;
      patterns[37391] = 25'b10010010_00001101_10011111_0;
      patterns[37392] = 25'b10010010_00001110_10100000_0;
      patterns[37393] = 25'b10010010_00001111_10100001_0;
      patterns[37394] = 25'b10010010_00010000_10100010_0;
      patterns[37395] = 25'b10010010_00010001_10100011_0;
      patterns[37396] = 25'b10010010_00010010_10100100_0;
      patterns[37397] = 25'b10010010_00010011_10100101_0;
      patterns[37398] = 25'b10010010_00010100_10100110_0;
      patterns[37399] = 25'b10010010_00010101_10100111_0;
      patterns[37400] = 25'b10010010_00010110_10101000_0;
      patterns[37401] = 25'b10010010_00010111_10101001_0;
      patterns[37402] = 25'b10010010_00011000_10101010_0;
      patterns[37403] = 25'b10010010_00011001_10101011_0;
      patterns[37404] = 25'b10010010_00011010_10101100_0;
      patterns[37405] = 25'b10010010_00011011_10101101_0;
      patterns[37406] = 25'b10010010_00011100_10101110_0;
      patterns[37407] = 25'b10010010_00011101_10101111_0;
      patterns[37408] = 25'b10010010_00011110_10110000_0;
      patterns[37409] = 25'b10010010_00011111_10110001_0;
      patterns[37410] = 25'b10010010_00100000_10110010_0;
      patterns[37411] = 25'b10010010_00100001_10110011_0;
      patterns[37412] = 25'b10010010_00100010_10110100_0;
      patterns[37413] = 25'b10010010_00100011_10110101_0;
      patterns[37414] = 25'b10010010_00100100_10110110_0;
      patterns[37415] = 25'b10010010_00100101_10110111_0;
      patterns[37416] = 25'b10010010_00100110_10111000_0;
      patterns[37417] = 25'b10010010_00100111_10111001_0;
      patterns[37418] = 25'b10010010_00101000_10111010_0;
      patterns[37419] = 25'b10010010_00101001_10111011_0;
      patterns[37420] = 25'b10010010_00101010_10111100_0;
      patterns[37421] = 25'b10010010_00101011_10111101_0;
      patterns[37422] = 25'b10010010_00101100_10111110_0;
      patterns[37423] = 25'b10010010_00101101_10111111_0;
      patterns[37424] = 25'b10010010_00101110_11000000_0;
      patterns[37425] = 25'b10010010_00101111_11000001_0;
      patterns[37426] = 25'b10010010_00110000_11000010_0;
      patterns[37427] = 25'b10010010_00110001_11000011_0;
      patterns[37428] = 25'b10010010_00110010_11000100_0;
      patterns[37429] = 25'b10010010_00110011_11000101_0;
      patterns[37430] = 25'b10010010_00110100_11000110_0;
      patterns[37431] = 25'b10010010_00110101_11000111_0;
      patterns[37432] = 25'b10010010_00110110_11001000_0;
      patterns[37433] = 25'b10010010_00110111_11001001_0;
      patterns[37434] = 25'b10010010_00111000_11001010_0;
      patterns[37435] = 25'b10010010_00111001_11001011_0;
      patterns[37436] = 25'b10010010_00111010_11001100_0;
      patterns[37437] = 25'b10010010_00111011_11001101_0;
      patterns[37438] = 25'b10010010_00111100_11001110_0;
      patterns[37439] = 25'b10010010_00111101_11001111_0;
      patterns[37440] = 25'b10010010_00111110_11010000_0;
      patterns[37441] = 25'b10010010_00111111_11010001_0;
      patterns[37442] = 25'b10010010_01000000_11010010_0;
      patterns[37443] = 25'b10010010_01000001_11010011_0;
      patterns[37444] = 25'b10010010_01000010_11010100_0;
      patterns[37445] = 25'b10010010_01000011_11010101_0;
      patterns[37446] = 25'b10010010_01000100_11010110_0;
      patterns[37447] = 25'b10010010_01000101_11010111_0;
      patterns[37448] = 25'b10010010_01000110_11011000_0;
      patterns[37449] = 25'b10010010_01000111_11011001_0;
      patterns[37450] = 25'b10010010_01001000_11011010_0;
      patterns[37451] = 25'b10010010_01001001_11011011_0;
      patterns[37452] = 25'b10010010_01001010_11011100_0;
      patterns[37453] = 25'b10010010_01001011_11011101_0;
      patterns[37454] = 25'b10010010_01001100_11011110_0;
      patterns[37455] = 25'b10010010_01001101_11011111_0;
      patterns[37456] = 25'b10010010_01001110_11100000_0;
      patterns[37457] = 25'b10010010_01001111_11100001_0;
      patterns[37458] = 25'b10010010_01010000_11100010_0;
      patterns[37459] = 25'b10010010_01010001_11100011_0;
      patterns[37460] = 25'b10010010_01010010_11100100_0;
      patterns[37461] = 25'b10010010_01010011_11100101_0;
      patterns[37462] = 25'b10010010_01010100_11100110_0;
      patterns[37463] = 25'b10010010_01010101_11100111_0;
      patterns[37464] = 25'b10010010_01010110_11101000_0;
      patterns[37465] = 25'b10010010_01010111_11101001_0;
      patterns[37466] = 25'b10010010_01011000_11101010_0;
      patterns[37467] = 25'b10010010_01011001_11101011_0;
      patterns[37468] = 25'b10010010_01011010_11101100_0;
      patterns[37469] = 25'b10010010_01011011_11101101_0;
      patterns[37470] = 25'b10010010_01011100_11101110_0;
      patterns[37471] = 25'b10010010_01011101_11101111_0;
      patterns[37472] = 25'b10010010_01011110_11110000_0;
      patterns[37473] = 25'b10010010_01011111_11110001_0;
      patterns[37474] = 25'b10010010_01100000_11110010_0;
      patterns[37475] = 25'b10010010_01100001_11110011_0;
      patterns[37476] = 25'b10010010_01100010_11110100_0;
      patterns[37477] = 25'b10010010_01100011_11110101_0;
      patterns[37478] = 25'b10010010_01100100_11110110_0;
      patterns[37479] = 25'b10010010_01100101_11110111_0;
      patterns[37480] = 25'b10010010_01100110_11111000_0;
      patterns[37481] = 25'b10010010_01100111_11111001_0;
      patterns[37482] = 25'b10010010_01101000_11111010_0;
      patterns[37483] = 25'b10010010_01101001_11111011_0;
      patterns[37484] = 25'b10010010_01101010_11111100_0;
      patterns[37485] = 25'b10010010_01101011_11111101_0;
      patterns[37486] = 25'b10010010_01101100_11111110_0;
      patterns[37487] = 25'b10010010_01101101_11111111_0;
      patterns[37488] = 25'b10010010_01101110_00000000_1;
      patterns[37489] = 25'b10010010_01101111_00000001_1;
      patterns[37490] = 25'b10010010_01110000_00000010_1;
      patterns[37491] = 25'b10010010_01110001_00000011_1;
      patterns[37492] = 25'b10010010_01110010_00000100_1;
      patterns[37493] = 25'b10010010_01110011_00000101_1;
      patterns[37494] = 25'b10010010_01110100_00000110_1;
      patterns[37495] = 25'b10010010_01110101_00000111_1;
      patterns[37496] = 25'b10010010_01110110_00001000_1;
      patterns[37497] = 25'b10010010_01110111_00001001_1;
      patterns[37498] = 25'b10010010_01111000_00001010_1;
      patterns[37499] = 25'b10010010_01111001_00001011_1;
      patterns[37500] = 25'b10010010_01111010_00001100_1;
      patterns[37501] = 25'b10010010_01111011_00001101_1;
      patterns[37502] = 25'b10010010_01111100_00001110_1;
      patterns[37503] = 25'b10010010_01111101_00001111_1;
      patterns[37504] = 25'b10010010_01111110_00010000_1;
      patterns[37505] = 25'b10010010_01111111_00010001_1;
      patterns[37506] = 25'b10010010_10000000_00010010_1;
      patterns[37507] = 25'b10010010_10000001_00010011_1;
      patterns[37508] = 25'b10010010_10000010_00010100_1;
      patterns[37509] = 25'b10010010_10000011_00010101_1;
      patterns[37510] = 25'b10010010_10000100_00010110_1;
      patterns[37511] = 25'b10010010_10000101_00010111_1;
      patterns[37512] = 25'b10010010_10000110_00011000_1;
      patterns[37513] = 25'b10010010_10000111_00011001_1;
      patterns[37514] = 25'b10010010_10001000_00011010_1;
      patterns[37515] = 25'b10010010_10001001_00011011_1;
      patterns[37516] = 25'b10010010_10001010_00011100_1;
      patterns[37517] = 25'b10010010_10001011_00011101_1;
      patterns[37518] = 25'b10010010_10001100_00011110_1;
      patterns[37519] = 25'b10010010_10001101_00011111_1;
      patterns[37520] = 25'b10010010_10001110_00100000_1;
      patterns[37521] = 25'b10010010_10001111_00100001_1;
      patterns[37522] = 25'b10010010_10010000_00100010_1;
      patterns[37523] = 25'b10010010_10010001_00100011_1;
      patterns[37524] = 25'b10010010_10010010_00100100_1;
      patterns[37525] = 25'b10010010_10010011_00100101_1;
      patterns[37526] = 25'b10010010_10010100_00100110_1;
      patterns[37527] = 25'b10010010_10010101_00100111_1;
      patterns[37528] = 25'b10010010_10010110_00101000_1;
      patterns[37529] = 25'b10010010_10010111_00101001_1;
      patterns[37530] = 25'b10010010_10011000_00101010_1;
      patterns[37531] = 25'b10010010_10011001_00101011_1;
      patterns[37532] = 25'b10010010_10011010_00101100_1;
      patterns[37533] = 25'b10010010_10011011_00101101_1;
      patterns[37534] = 25'b10010010_10011100_00101110_1;
      patterns[37535] = 25'b10010010_10011101_00101111_1;
      patterns[37536] = 25'b10010010_10011110_00110000_1;
      patterns[37537] = 25'b10010010_10011111_00110001_1;
      patterns[37538] = 25'b10010010_10100000_00110010_1;
      patterns[37539] = 25'b10010010_10100001_00110011_1;
      patterns[37540] = 25'b10010010_10100010_00110100_1;
      patterns[37541] = 25'b10010010_10100011_00110101_1;
      patterns[37542] = 25'b10010010_10100100_00110110_1;
      patterns[37543] = 25'b10010010_10100101_00110111_1;
      patterns[37544] = 25'b10010010_10100110_00111000_1;
      patterns[37545] = 25'b10010010_10100111_00111001_1;
      patterns[37546] = 25'b10010010_10101000_00111010_1;
      patterns[37547] = 25'b10010010_10101001_00111011_1;
      patterns[37548] = 25'b10010010_10101010_00111100_1;
      patterns[37549] = 25'b10010010_10101011_00111101_1;
      patterns[37550] = 25'b10010010_10101100_00111110_1;
      patterns[37551] = 25'b10010010_10101101_00111111_1;
      patterns[37552] = 25'b10010010_10101110_01000000_1;
      patterns[37553] = 25'b10010010_10101111_01000001_1;
      patterns[37554] = 25'b10010010_10110000_01000010_1;
      patterns[37555] = 25'b10010010_10110001_01000011_1;
      patterns[37556] = 25'b10010010_10110010_01000100_1;
      patterns[37557] = 25'b10010010_10110011_01000101_1;
      patterns[37558] = 25'b10010010_10110100_01000110_1;
      patterns[37559] = 25'b10010010_10110101_01000111_1;
      patterns[37560] = 25'b10010010_10110110_01001000_1;
      patterns[37561] = 25'b10010010_10110111_01001001_1;
      patterns[37562] = 25'b10010010_10111000_01001010_1;
      patterns[37563] = 25'b10010010_10111001_01001011_1;
      patterns[37564] = 25'b10010010_10111010_01001100_1;
      patterns[37565] = 25'b10010010_10111011_01001101_1;
      patterns[37566] = 25'b10010010_10111100_01001110_1;
      patterns[37567] = 25'b10010010_10111101_01001111_1;
      patterns[37568] = 25'b10010010_10111110_01010000_1;
      patterns[37569] = 25'b10010010_10111111_01010001_1;
      patterns[37570] = 25'b10010010_11000000_01010010_1;
      patterns[37571] = 25'b10010010_11000001_01010011_1;
      patterns[37572] = 25'b10010010_11000010_01010100_1;
      patterns[37573] = 25'b10010010_11000011_01010101_1;
      patterns[37574] = 25'b10010010_11000100_01010110_1;
      patterns[37575] = 25'b10010010_11000101_01010111_1;
      patterns[37576] = 25'b10010010_11000110_01011000_1;
      patterns[37577] = 25'b10010010_11000111_01011001_1;
      patterns[37578] = 25'b10010010_11001000_01011010_1;
      patterns[37579] = 25'b10010010_11001001_01011011_1;
      patterns[37580] = 25'b10010010_11001010_01011100_1;
      patterns[37581] = 25'b10010010_11001011_01011101_1;
      patterns[37582] = 25'b10010010_11001100_01011110_1;
      patterns[37583] = 25'b10010010_11001101_01011111_1;
      patterns[37584] = 25'b10010010_11001110_01100000_1;
      patterns[37585] = 25'b10010010_11001111_01100001_1;
      patterns[37586] = 25'b10010010_11010000_01100010_1;
      patterns[37587] = 25'b10010010_11010001_01100011_1;
      patterns[37588] = 25'b10010010_11010010_01100100_1;
      patterns[37589] = 25'b10010010_11010011_01100101_1;
      patterns[37590] = 25'b10010010_11010100_01100110_1;
      patterns[37591] = 25'b10010010_11010101_01100111_1;
      patterns[37592] = 25'b10010010_11010110_01101000_1;
      patterns[37593] = 25'b10010010_11010111_01101001_1;
      patterns[37594] = 25'b10010010_11011000_01101010_1;
      patterns[37595] = 25'b10010010_11011001_01101011_1;
      patterns[37596] = 25'b10010010_11011010_01101100_1;
      patterns[37597] = 25'b10010010_11011011_01101101_1;
      patterns[37598] = 25'b10010010_11011100_01101110_1;
      patterns[37599] = 25'b10010010_11011101_01101111_1;
      patterns[37600] = 25'b10010010_11011110_01110000_1;
      patterns[37601] = 25'b10010010_11011111_01110001_1;
      patterns[37602] = 25'b10010010_11100000_01110010_1;
      patterns[37603] = 25'b10010010_11100001_01110011_1;
      patterns[37604] = 25'b10010010_11100010_01110100_1;
      patterns[37605] = 25'b10010010_11100011_01110101_1;
      patterns[37606] = 25'b10010010_11100100_01110110_1;
      patterns[37607] = 25'b10010010_11100101_01110111_1;
      patterns[37608] = 25'b10010010_11100110_01111000_1;
      patterns[37609] = 25'b10010010_11100111_01111001_1;
      patterns[37610] = 25'b10010010_11101000_01111010_1;
      patterns[37611] = 25'b10010010_11101001_01111011_1;
      patterns[37612] = 25'b10010010_11101010_01111100_1;
      patterns[37613] = 25'b10010010_11101011_01111101_1;
      patterns[37614] = 25'b10010010_11101100_01111110_1;
      patterns[37615] = 25'b10010010_11101101_01111111_1;
      patterns[37616] = 25'b10010010_11101110_10000000_1;
      patterns[37617] = 25'b10010010_11101111_10000001_1;
      patterns[37618] = 25'b10010010_11110000_10000010_1;
      patterns[37619] = 25'b10010010_11110001_10000011_1;
      patterns[37620] = 25'b10010010_11110010_10000100_1;
      patterns[37621] = 25'b10010010_11110011_10000101_1;
      patterns[37622] = 25'b10010010_11110100_10000110_1;
      patterns[37623] = 25'b10010010_11110101_10000111_1;
      patterns[37624] = 25'b10010010_11110110_10001000_1;
      patterns[37625] = 25'b10010010_11110111_10001001_1;
      patterns[37626] = 25'b10010010_11111000_10001010_1;
      patterns[37627] = 25'b10010010_11111001_10001011_1;
      patterns[37628] = 25'b10010010_11111010_10001100_1;
      patterns[37629] = 25'b10010010_11111011_10001101_1;
      patterns[37630] = 25'b10010010_11111100_10001110_1;
      patterns[37631] = 25'b10010010_11111101_10001111_1;
      patterns[37632] = 25'b10010010_11111110_10010000_1;
      patterns[37633] = 25'b10010010_11111111_10010001_1;
      patterns[37634] = 25'b10010011_00000000_10010011_0;
      patterns[37635] = 25'b10010011_00000001_10010100_0;
      patterns[37636] = 25'b10010011_00000010_10010101_0;
      patterns[37637] = 25'b10010011_00000011_10010110_0;
      patterns[37638] = 25'b10010011_00000100_10010111_0;
      patterns[37639] = 25'b10010011_00000101_10011000_0;
      patterns[37640] = 25'b10010011_00000110_10011001_0;
      patterns[37641] = 25'b10010011_00000111_10011010_0;
      patterns[37642] = 25'b10010011_00001000_10011011_0;
      patterns[37643] = 25'b10010011_00001001_10011100_0;
      patterns[37644] = 25'b10010011_00001010_10011101_0;
      patterns[37645] = 25'b10010011_00001011_10011110_0;
      patterns[37646] = 25'b10010011_00001100_10011111_0;
      patterns[37647] = 25'b10010011_00001101_10100000_0;
      patterns[37648] = 25'b10010011_00001110_10100001_0;
      patterns[37649] = 25'b10010011_00001111_10100010_0;
      patterns[37650] = 25'b10010011_00010000_10100011_0;
      patterns[37651] = 25'b10010011_00010001_10100100_0;
      patterns[37652] = 25'b10010011_00010010_10100101_0;
      patterns[37653] = 25'b10010011_00010011_10100110_0;
      patterns[37654] = 25'b10010011_00010100_10100111_0;
      patterns[37655] = 25'b10010011_00010101_10101000_0;
      patterns[37656] = 25'b10010011_00010110_10101001_0;
      patterns[37657] = 25'b10010011_00010111_10101010_0;
      patterns[37658] = 25'b10010011_00011000_10101011_0;
      patterns[37659] = 25'b10010011_00011001_10101100_0;
      patterns[37660] = 25'b10010011_00011010_10101101_0;
      patterns[37661] = 25'b10010011_00011011_10101110_0;
      patterns[37662] = 25'b10010011_00011100_10101111_0;
      patterns[37663] = 25'b10010011_00011101_10110000_0;
      patterns[37664] = 25'b10010011_00011110_10110001_0;
      patterns[37665] = 25'b10010011_00011111_10110010_0;
      patterns[37666] = 25'b10010011_00100000_10110011_0;
      patterns[37667] = 25'b10010011_00100001_10110100_0;
      patterns[37668] = 25'b10010011_00100010_10110101_0;
      patterns[37669] = 25'b10010011_00100011_10110110_0;
      patterns[37670] = 25'b10010011_00100100_10110111_0;
      patterns[37671] = 25'b10010011_00100101_10111000_0;
      patterns[37672] = 25'b10010011_00100110_10111001_0;
      patterns[37673] = 25'b10010011_00100111_10111010_0;
      patterns[37674] = 25'b10010011_00101000_10111011_0;
      patterns[37675] = 25'b10010011_00101001_10111100_0;
      patterns[37676] = 25'b10010011_00101010_10111101_0;
      patterns[37677] = 25'b10010011_00101011_10111110_0;
      patterns[37678] = 25'b10010011_00101100_10111111_0;
      patterns[37679] = 25'b10010011_00101101_11000000_0;
      patterns[37680] = 25'b10010011_00101110_11000001_0;
      patterns[37681] = 25'b10010011_00101111_11000010_0;
      patterns[37682] = 25'b10010011_00110000_11000011_0;
      patterns[37683] = 25'b10010011_00110001_11000100_0;
      patterns[37684] = 25'b10010011_00110010_11000101_0;
      patterns[37685] = 25'b10010011_00110011_11000110_0;
      patterns[37686] = 25'b10010011_00110100_11000111_0;
      patterns[37687] = 25'b10010011_00110101_11001000_0;
      patterns[37688] = 25'b10010011_00110110_11001001_0;
      patterns[37689] = 25'b10010011_00110111_11001010_0;
      patterns[37690] = 25'b10010011_00111000_11001011_0;
      patterns[37691] = 25'b10010011_00111001_11001100_0;
      patterns[37692] = 25'b10010011_00111010_11001101_0;
      patterns[37693] = 25'b10010011_00111011_11001110_0;
      patterns[37694] = 25'b10010011_00111100_11001111_0;
      patterns[37695] = 25'b10010011_00111101_11010000_0;
      patterns[37696] = 25'b10010011_00111110_11010001_0;
      patterns[37697] = 25'b10010011_00111111_11010010_0;
      patterns[37698] = 25'b10010011_01000000_11010011_0;
      patterns[37699] = 25'b10010011_01000001_11010100_0;
      patterns[37700] = 25'b10010011_01000010_11010101_0;
      patterns[37701] = 25'b10010011_01000011_11010110_0;
      patterns[37702] = 25'b10010011_01000100_11010111_0;
      patterns[37703] = 25'b10010011_01000101_11011000_0;
      patterns[37704] = 25'b10010011_01000110_11011001_0;
      patterns[37705] = 25'b10010011_01000111_11011010_0;
      patterns[37706] = 25'b10010011_01001000_11011011_0;
      patterns[37707] = 25'b10010011_01001001_11011100_0;
      patterns[37708] = 25'b10010011_01001010_11011101_0;
      patterns[37709] = 25'b10010011_01001011_11011110_0;
      patterns[37710] = 25'b10010011_01001100_11011111_0;
      patterns[37711] = 25'b10010011_01001101_11100000_0;
      patterns[37712] = 25'b10010011_01001110_11100001_0;
      patterns[37713] = 25'b10010011_01001111_11100010_0;
      patterns[37714] = 25'b10010011_01010000_11100011_0;
      patterns[37715] = 25'b10010011_01010001_11100100_0;
      patterns[37716] = 25'b10010011_01010010_11100101_0;
      patterns[37717] = 25'b10010011_01010011_11100110_0;
      patterns[37718] = 25'b10010011_01010100_11100111_0;
      patterns[37719] = 25'b10010011_01010101_11101000_0;
      patterns[37720] = 25'b10010011_01010110_11101001_0;
      patterns[37721] = 25'b10010011_01010111_11101010_0;
      patterns[37722] = 25'b10010011_01011000_11101011_0;
      patterns[37723] = 25'b10010011_01011001_11101100_0;
      patterns[37724] = 25'b10010011_01011010_11101101_0;
      patterns[37725] = 25'b10010011_01011011_11101110_0;
      patterns[37726] = 25'b10010011_01011100_11101111_0;
      patterns[37727] = 25'b10010011_01011101_11110000_0;
      patterns[37728] = 25'b10010011_01011110_11110001_0;
      patterns[37729] = 25'b10010011_01011111_11110010_0;
      patterns[37730] = 25'b10010011_01100000_11110011_0;
      patterns[37731] = 25'b10010011_01100001_11110100_0;
      patterns[37732] = 25'b10010011_01100010_11110101_0;
      patterns[37733] = 25'b10010011_01100011_11110110_0;
      patterns[37734] = 25'b10010011_01100100_11110111_0;
      patterns[37735] = 25'b10010011_01100101_11111000_0;
      patterns[37736] = 25'b10010011_01100110_11111001_0;
      patterns[37737] = 25'b10010011_01100111_11111010_0;
      patterns[37738] = 25'b10010011_01101000_11111011_0;
      patterns[37739] = 25'b10010011_01101001_11111100_0;
      patterns[37740] = 25'b10010011_01101010_11111101_0;
      patterns[37741] = 25'b10010011_01101011_11111110_0;
      patterns[37742] = 25'b10010011_01101100_11111111_0;
      patterns[37743] = 25'b10010011_01101101_00000000_1;
      patterns[37744] = 25'b10010011_01101110_00000001_1;
      patterns[37745] = 25'b10010011_01101111_00000010_1;
      patterns[37746] = 25'b10010011_01110000_00000011_1;
      patterns[37747] = 25'b10010011_01110001_00000100_1;
      patterns[37748] = 25'b10010011_01110010_00000101_1;
      patterns[37749] = 25'b10010011_01110011_00000110_1;
      patterns[37750] = 25'b10010011_01110100_00000111_1;
      patterns[37751] = 25'b10010011_01110101_00001000_1;
      patterns[37752] = 25'b10010011_01110110_00001001_1;
      patterns[37753] = 25'b10010011_01110111_00001010_1;
      patterns[37754] = 25'b10010011_01111000_00001011_1;
      patterns[37755] = 25'b10010011_01111001_00001100_1;
      patterns[37756] = 25'b10010011_01111010_00001101_1;
      patterns[37757] = 25'b10010011_01111011_00001110_1;
      patterns[37758] = 25'b10010011_01111100_00001111_1;
      patterns[37759] = 25'b10010011_01111101_00010000_1;
      patterns[37760] = 25'b10010011_01111110_00010001_1;
      patterns[37761] = 25'b10010011_01111111_00010010_1;
      patterns[37762] = 25'b10010011_10000000_00010011_1;
      patterns[37763] = 25'b10010011_10000001_00010100_1;
      patterns[37764] = 25'b10010011_10000010_00010101_1;
      patterns[37765] = 25'b10010011_10000011_00010110_1;
      patterns[37766] = 25'b10010011_10000100_00010111_1;
      patterns[37767] = 25'b10010011_10000101_00011000_1;
      patterns[37768] = 25'b10010011_10000110_00011001_1;
      patterns[37769] = 25'b10010011_10000111_00011010_1;
      patterns[37770] = 25'b10010011_10001000_00011011_1;
      patterns[37771] = 25'b10010011_10001001_00011100_1;
      patterns[37772] = 25'b10010011_10001010_00011101_1;
      patterns[37773] = 25'b10010011_10001011_00011110_1;
      patterns[37774] = 25'b10010011_10001100_00011111_1;
      patterns[37775] = 25'b10010011_10001101_00100000_1;
      patterns[37776] = 25'b10010011_10001110_00100001_1;
      patterns[37777] = 25'b10010011_10001111_00100010_1;
      patterns[37778] = 25'b10010011_10010000_00100011_1;
      patterns[37779] = 25'b10010011_10010001_00100100_1;
      patterns[37780] = 25'b10010011_10010010_00100101_1;
      patterns[37781] = 25'b10010011_10010011_00100110_1;
      patterns[37782] = 25'b10010011_10010100_00100111_1;
      patterns[37783] = 25'b10010011_10010101_00101000_1;
      patterns[37784] = 25'b10010011_10010110_00101001_1;
      patterns[37785] = 25'b10010011_10010111_00101010_1;
      patterns[37786] = 25'b10010011_10011000_00101011_1;
      patterns[37787] = 25'b10010011_10011001_00101100_1;
      patterns[37788] = 25'b10010011_10011010_00101101_1;
      patterns[37789] = 25'b10010011_10011011_00101110_1;
      patterns[37790] = 25'b10010011_10011100_00101111_1;
      patterns[37791] = 25'b10010011_10011101_00110000_1;
      patterns[37792] = 25'b10010011_10011110_00110001_1;
      patterns[37793] = 25'b10010011_10011111_00110010_1;
      patterns[37794] = 25'b10010011_10100000_00110011_1;
      patterns[37795] = 25'b10010011_10100001_00110100_1;
      patterns[37796] = 25'b10010011_10100010_00110101_1;
      patterns[37797] = 25'b10010011_10100011_00110110_1;
      patterns[37798] = 25'b10010011_10100100_00110111_1;
      patterns[37799] = 25'b10010011_10100101_00111000_1;
      patterns[37800] = 25'b10010011_10100110_00111001_1;
      patterns[37801] = 25'b10010011_10100111_00111010_1;
      patterns[37802] = 25'b10010011_10101000_00111011_1;
      patterns[37803] = 25'b10010011_10101001_00111100_1;
      patterns[37804] = 25'b10010011_10101010_00111101_1;
      patterns[37805] = 25'b10010011_10101011_00111110_1;
      patterns[37806] = 25'b10010011_10101100_00111111_1;
      patterns[37807] = 25'b10010011_10101101_01000000_1;
      patterns[37808] = 25'b10010011_10101110_01000001_1;
      patterns[37809] = 25'b10010011_10101111_01000010_1;
      patterns[37810] = 25'b10010011_10110000_01000011_1;
      patterns[37811] = 25'b10010011_10110001_01000100_1;
      patterns[37812] = 25'b10010011_10110010_01000101_1;
      patterns[37813] = 25'b10010011_10110011_01000110_1;
      patterns[37814] = 25'b10010011_10110100_01000111_1;
      patterns[37815] = 25'b10010011_10110101_01001000_1;
      patterns[37816] = 25'b10010011_10110110_01001001_1;
      patterns[37817] = 25'b10010011_10110111_01001010_1;
      patterns[37818] = 25'b10010011_10111000_01001011_1;
      patterns[37819] = 25'b10010011_10111001_01001100_1;
      patterns[37820] = 25'b10010011_10111010_01001101_1;
      patterns[37821] = 25'b10010011_10111011_01001110_1;
      patterns[37822] = 25'b10010011_10111100_01001111_1;
      patterns[37823] = 25'b10010011_10111101_01010000_1;
      patterns[37824] = 25'b10010011_10111110_01010001_1;
      patterns[37825] = 25'b10010011_10111111_01010010_1;
      patterns[37826] = 25'b10010011_11000000_01010011_1;
      patterns[37827] = 25'b10010011_11000001_01010100_1;
      patterns[37828] = 25'b10010011_11000010_01010101_1;
      patterns[37829] = 25'b10010011_11000011_01010110_1;
      patterns[37830] = 25'b10010011_11000100_01010111_1;
      patterns[37831] = 25'b10010011_11000101_01011000_1;
      patterns[37832] = 25'b10010011_11000110_01011001_1;
      patterns[37833] = 25'b10010011_11000111_01011010_1;
      patterns[37834] = 25'b10010011_11001000_01011011_1;
      patterns[37835] = 25'b10010011_11001001_01011100_1;
      patterns[37836] = 25'b10010011_11001010_01011101_1;
      patterns[37837] = 25'b10010011_11001011_01011110_1;
      patterns[37838] = 25'b10010011_11001100_01011111_1;
      patterns[37839] = 25'b10010011_11001101_01100000_1;
      patterns[37840] = 25'b10010011_11001110_01100001_1;
      patterns[37841] = 25'b10010011_11001111_01100010_1;
      patterns[37842] = 25'b10010011_11010000_01100011_1;
      patterns[37843] = 25'b10010011_11010001_01100100_1;
      patterns[37844] = 25'b10010011_11010010_01100101_1;
      patterns[37845] = 25'b10010011_11010011_01100110_1;
      patterns[37846] = 25'b10010011_11010100_01100111_1;
      patterns[37847] = 25'b10010011_11010101_01101000_1;
      patterns[37848] = 25'b10010011_11010110_01101001_1;
      patterns[37849] = 25'b10010011_11010111_01101010_1;
      patterns[37850] = 25'b10010011_11011000_01101011_1;
      patterns[37851] = 25'b10010011_11011001_01101100_1;
      patterns[37852] = 25'b10010011_11011010_01101101_1;
      patterns[37853] = 25'b10010011_11011011_01101110_1;
      patterns[37854] = 25'b10010011_11011100_01101111_1;
      patterns[37855] = 25'b10010011_11011101_01110000_1;
      patterns[37856] = 25'b10010011_11011110_01110001_1;
      patterns[37857] = 25'b10010011_11011111_01110010_1;
      patterns[37858] = 25'b10010011_11100000_01110011_1;
      patterns[37859] = 25'b10010011_11100001_01110100_1;
      patterns[37860] = 25'b10010011_11100010_01110101_1;
      patterns[37861] = 25'b10010011_11100011_01110110_1;
      patterns[37862] = 25'b10010011_11100100_01110111_1;
      patterns[37863] = 25'b10010011_11100101_01111000_1;
      patterns[37864] = 25'b10010011_11100110_01111001_1;
      patterns[37865] = 25'b10010011_11100111_01111010_1;
      patterns[37866] = 25'b10010011_11101000_01111011_1;
      patterns[37867] = 25'b10010011_11101001_01111100_1;
      patterns[37868] = 25'b10010011_11101010_01111101_1;
      patterns[37869] = 25'b10010011_11101011_01111110_1;
      patterns[37870] = 25'b10010011_11101100_01111111_1;
      patterns[37871] = 25'b10010011_11101101_10000000_1;
      patterns[37872] = 25'b10010011_11101110_10000001_1;
      patterns[37873] = 25'b10010011_11101111_10000010_1;
      patterns[37874] = 25'b10010011_11110000_10000011_1;
      patterns[37875] = 25'b10010011_11110001_10000100_1;
      patterns[37876] = 25'b10010011_11110010_10000101_1;
      patterns[37877] = 25'b10010011_11110011_10000110_1;
      patterns[37878] = 25'b10010011_11110100_10000111_1;
      patterns[37879] = 25'b10010011_11110101_10001000_1;
      patterns[37880] = 25'b10010011_11110110_10001001_1;
      patterns[37881] = 25'b10010011_11110111_10001010_1;
      patterns[37882] = 25'b10010011_11111000_10001011_1;
      patterns[37883] = 25'b10010011_11111001_10001100_1;
      patterns[37884] = 25'b10010011_11111010_10001101_1;
      patterns[37885] = 25'b10010011_11111011_10001110_1;
      patterns[37886] = 25'b10010011_11111100_10001111_1;
      patterns[37887] = 25'b10010011_11111101_10010000_1;
      patterns[37888] = 25'b10010011_11111110_10010001_1;
      patterns[37889] = 25'b10010011_11111111_10010010_1;
      patterns[37890] = 25'b10010100_00000000_10010100_0;
      patterns[37891] = 25'b10010100_00000001_10010101_0;
      patterns[37892] = 25'b10010100_00000010_10010110_0;
      patterns[37893] = 25'b10010100_00000011_10010111_0;
      patterns[37894] = 25'b10010100_00000100_10011000_0;
      patterns[37895] = 25'b10010100_00000101_10011001_0;
      patterns[37896] = 25'b10010100_00000110_10011010_0;
      patterns[37897] = 25'b10010100_00000111_10011011_0;
      patterns[37898] = 25'b10010100_00001000_10011100_0;
      patterns[37899] = 25'b10010100_00001001_10011101_0;
      patterns[37900] = 25'b10010100_00001010_10011110_0;
      patterns[37901] = 25'b10010100_00001011_10011111_0;
      patterns[37902] = 25'b10010100_00001100_10100000_0;
      patterns[37903] = 25'b10010100_00001101_10100001_0;
      patterns[37904] = 25'b10010100_00001110_10100010_0;
      patterns[37905] = 25'b10010100_00001111_10100011_0;
      patterns[37906] = 25'b10010100_00010000_10100100_0;
      patterns[37907] = 25'b10010100_00010001_10100101_0;
      patterns[37908] = 25'b10010100_00010010_10100110_0;
      patterns[37909] = 25'b10010100_00010011_10100111_0;
      patterns[37910] = 25'b10010100_00010100_10101000_0;
      patterns[37911] = 25'b10010100_00010101_10101001_0;
      patterns[37912] = 25'b10010100_00010110_10101010_0;
      patterns[37913] = 25'b10010100_00010111_10101011_0;
      patterns[37914] = 25'b10010100_00011000_10101100_0;
      patterns[37915] = 25'b10010100_00011001_10101101_0;
      patterns[37916] = 25'b10010100_00011010_10101110_0;
      patterns[37917] = 25'b10010100_00011011_10101111_0;
      patterns[37918] = 25'b10010100_00011100_10110000_0;
      patterns[37919] = 25'b10010100_00011101_10110001_0;
      patterns[37920] = 25'b10010100_00011110_10110010_0;
      patterns[37921] = 25'b10010100_00011111_10110011_0;
      patterns[37922] = 25'b10010100_00100000_10110100_0;
      patterns[37923] = 25'b10010100_00100001_10110101_0;
      patterns[37924] = 25'b10010100_00100010_10110110_0;
      patterns[37925] = 25'b10010100_00100011_10110111_0;
      patterns[37926] = 25'b10010100_00100100_10111000_0;
      patterns[37927] = 25'b10010100_00100101_10111001_0;
      patterns[37928] = 25'b10010100_00100110_10111010_0;
      patterns[37929] = 25'b10010100_00100111_10111011_0;
      patterns[37930] = 25'b10010100_00101000_10111100_0;
      patterns[37931] = 25'b10010100_00101001_10111101_0;
      patterns[37932] = 25'b10010100_00101010_10111110_0;
      patterns[37933] = 25'b10010100_00101011_10111111_0;
      patterns[37934] = 25'b10010100_00101100_11000000_0;
      patterns[37935] = 25'b10010100_00101101_11000001_0;
      patterns[37936] = 25'b10010100_00101110_11000010_0;
      patterns[37937] = 25'b10010100_00101111_11000011_0;
      patterns[37938] = 25'b10010100_00110000_11000100_0;
      patterns[37939] = 25'b10010100_00110001_11000101_0;
      patterns[37940] = 25'b10010100_00110010_11000110_0;
      patterns[37941] = 25'b10010100_00110011_11000111_0;
      patterns[37942] = 25'b10010100_00110100_11001000_0;
      patterns[37943] = 25'b10010100_00110101_11001001_0;
      patterns[37944] = 25'b10010100_00110110_11001010_0;
      patterns[37945] = 25'b10010100_00110111_11001011_0;
      patterns[37946] = 25'b10010100_00111000_11001100_0;
      patterns[37947] = 25'b10010100_00111001_11001101_0;
      patterns[37948] = 25'b10010100_00111010_11001110_0;
      patterns[37949] = 25'b10010100_00111011_11001111_0;
      patterns[37950] = 25'b10010100_00111100_11010000_0;
      patterns[37951] = 25'b10010100_00111101_11010001_0;
      patterns[37952] = 25'b10010100_00111110_11010010_0;
      patterns[37953] = 25'b10010100_00111111_11010011_0;
      patterns[37954] = 25'b10010100_01000000_11010100_0;
      patterns[37955] = 25'b10010100_01000001_11010101_0;
      patterns[37956] = 25'b10010100_01000010_11010110_0;
      patterns[37957] = 25'b10010100_01000011_11010111_0;
      patterns[37958] = 25'b10010100_01000100_11011000_0;
      patterns[37959] = 25'b10010100_01000101_11011001_0;
      patterns[37960] = 25'b10010100_01000110_11011010_0;
      patterns[37961] = 25'b10010100_01000111_11011011_0;
      patterns[37962] = 25'b10010100_01001000_11011100_0;
      patterns[37963] = 25'b10010100_01001001_11011101_0;
      patterns[37964] = 25'b10010100_01001010_11011110_0;
      patterns[37965] = 25'b10010100_01001011_11011111_0;
      patterns[37966] = 25'b10010100_01001100_11100000_0;
      patterns[37967] = 25'b10010100_01001101_11100001_0;
      patterns[37968] = 25'b10010100_01001110_11100010_0;
      patterns[37969] = 25'b10010100_01001111_11100011_0;
      patterns[37970] = 25'b10010100_01010000_11100100_0;
      patterns[37971] = 25'b10010100_01010001_11100101_0;
      patterns[37972] = 25'b10010100_01010010_11100110_0;
      patterns[37973] = 25'b10010100_01010011_11100111_0;
      patterns[37974] = 25'b10010100_01010100_11101000_0;
      patterns[37975] = 25'b10010100_01010101_11101001_0;
      patterns[37976] = 25'b10010100_01010110_11101010_0;
      patterns[37977] = 25'b10010100_01010111_11101011_0;
      patterns[37978] = 25'b10010100_01011000_11101100_0;
      patterns[37979] = 25'b10010100_01011001_11101101_0;
      patterns[37980] = 25'b10010100_01011010_11101110_0;
      patterns[37981] = 25'b10010100_01011011_11101111_0;
      patterns[37982] = 25'b10010100_01011100_11110000_0;
      patterns[37983] = 25'b10010100_01011101_11110001_0;
      patterns[37984] = 25'b10010100_01011110_11110010_0;
      patterns[37985] = 25'b10010100_01011111_11110011_0;
      patterns[37986] = 25'b10010100_01100000_11110100_0;
      patterns[37987] = 25'b10010100_01100001_11110101_0;
      patterns[37988] = 25'b10010100_01100010_11110110_0;
      patterns[37989] = 25'b10010100_01100011_11110111_0;
      patterns[37990] = 25'b10010100_01100100_11111000_0;
      patterns[37991] = 25'b10010100_01100101_11111001_0;
      patterns[37992] = 25'b10010100_01100110_11111010_0;
      patterns[37993] = 25'b10010100_01100111_11111011_0;
      patterns[37994] = 25'b10010100_01101000_11111100_0;
      patterns[37995] = 25'b10010100_01101001_11111101_0;
      patterns[37996] = 25'b10010100_01101010_11111110_0;
      patterns[37997] = 25'b10010100_01101011_11111111_0;
      patterns[37998] = 25'b10010100_01101100_00000000_1;
      patterns[37999] = 25'b10010100_01101101_00000001_1;
      patterns[38000] = 25'b10010100_01101110_00000010_1;
      patterns[38001] = 25'b10010100_01101111_00000011_1;
      patterns[38002] = 25'b10010100_01110000_00000100_1;
      patterns[38003] = 25'b10010100_01110001_00000101_1;
      patterns[38004] = 25'b10010100_01110010_00000110_1;
      patterns[38005] = 25'b10010100_01110011_00000111_1;
      patterns[38006] = 25'b10010100_01110100_00001000_1;
      patterns[38007] = 25'b10010100_01110101_00001001_1;
      patterns[38008] = 25'b10010100_01110110_00001010_1;
      patterns[38009] = 25'b10010100_01110111_00001011_1;
      patterns[38010] = 25'b10010100_01111000_00001100_1;
      patterns[38011] = 25'b10010100_01111001_00001101_1;
      patterns[38012] = 25'b10010100_01111010_00001110_1;
      patterns[38013] = 25'b10010100_01111011_00001111_1;
      patterns[38014] = 25'b10010100_01111100_00010000_1;
      patterns[38015] = 25'b10010100_01111101_00010001_1;
      patterns[38016] = 25'b10010100_01111110_00010010_1;
      patterns[38017] = 25'b10010100_01111111_00010011_1;
      patterns[38018] = 25'b10010100_10000000_00010100_1;
      patterns[38019] = 25'b10010100_10000001_00010101_1;
      patterns[38020] = 25'b10010100_10000010_00010110_1;
      patterns[38021] = 25'b10010100_10000011_00010111_1;
      patterns[38022] = 25'b10010100_10000100_00011000_1;
      patterns[38023] = 25'b10010100_10000101_00011001_1;
      patterns[38024] = 25'b10010100_10000110_00011010_1;
      patterns[38025] = 25'b10010100_10000111_00011011_1;
      patterns[38026] = 25'b10010100_10001000_00011100_1;
      patterns[38027] = 25'b10010100_10001001_00011101_1;
      patterns[38028] = 25'b10010100_10001010_00011110_1;
      patterns[38029] = 25'b10010100_10001011_00011111_1;
      patterns[38030] = 25'b10010100_10001100_00100000_1;
      patterns[38031] = 25'b10010100_10001101_00100001_1;
      patterns[38032] = 25'b10010100_10001110_00100010_1;
      patterns[38033] = 25'b10010100_10001111_00100011_1;
      patterns[38034] = 25'b10010100_10010000_00100100_1;
      patterns[38035] = 25'b10010100_10010001_00100101_1;
      patterns[38036] = 25'b10010100_10010010_00100110_1;
      patterns[38037] = 25'b10010100_10010011_00100111_1;
      patterns[38038] = 25'b10010100_10010100_00101000_1;
      patterns[38039] = 25'b10010100_10010101_00101001_1;
      patterns[38040] = 25'b10010100_10010110_00101010_1;
      patterns[38041] = 25'b10010100_10010111_00101011_1;
      patterns[38042] = 25'b10010100_10011000_00101100_1;
      patterns[38043] = 25'b10010100_10011001_00101101_1;
      patterns[38044] = 25'b10010100_10011010_00101110_1;
      patterns[38045] = 25'b10010100_10011011_00101111_1;
      patterns[38046] = 25'b10010100_10011100_00110000_1;
      patterns[38047] = 25'b10010100_10011101_00110001_1;
      patterns[38048] = 25'b10010100_10011110_00110010_1;
      patterns[38049] = 25'b10010100_10011111_00110011_1;
      patterns[38050] = 25'b10010100_10100000_00110100_1;
      patterns[38051] = 25'b10010100_10100001_00110101_1;
      patterns[38052] = 25'b10010100_10100010_00110110_1;
      patterns[38053] = 25'b10010100_10100011_00110111_1;
      patterns[38054] = 25'b10010100_10100100_00111000_1;
      patterns[38055] = 25'b10010100_10100101_00111001_1;
      patterns[38056] = 25'b10010100_10100110_00111010_1;
      patterns[38057] = 25'b10010100_10100111_00111011_1;
      patterns[38058] = 25'b10010100_10101000_00111100_1;
      patterns[38059] = 25'b10010100_10101001_00111101_1;
      patterns[38060] = 25'b10010100_10101010_00111110_1;
      patterns[38061] = 25'b10010100_10101011_00111111_1;
      patterns[38062] = 25'b10010100_10101100_01000000_1;
      patterns[38063] = 25'b10010100_10101101_01000001_1;
      patterns[38064] = 25'b10010100_10101110_01000010_1;
      patterns[38065] = 25'b10010100_10101111_01000011_1;
      patterns[38066] = 25'b10010100_10110000_01000100_1;
      patterns[38067] = 25'b10010100_10110001_01000101_1;
      patterns[38068] = 25'b10010100_10110010_01000110_1;
      patterns[38069] = 25'b10010100_10110011_01000111_1;
      patterns[38070] = 25'b10010100_10110100_01001000_1;
      patterns[38071] = 25'b10010100_10110101_01001001_1;
      patterns[38072] = 25'b10010100_10110110_01001010_1;
      patterns[38073] = 25'b10010100_10110111_01001011_1;
      patterns[38074] = 25'b10010100_10111000_01001100_1;
      patterns[38075] = 25'b10010100_10111001_01001101_1;
      patterns[38076] = 25'b10010100_10111010_01001110_1;
      patterns[38077] = 25'b10010100_10111011_01001111_1;
      patterns[38078] = 25'b10010100_10111100_01010000_1;
      patterns[38079] = 25'b10010100_10111101_01010001_1;
      patterns[38080] = 25'b10010100_10111110_01010010_1;
      patterns[38081] = 25'b10010100_10111111_01010011_1;
      patterns[38082] = 25'b10010100_11000000_01010100_1;
      patterns[38083] = 25'b10010100_11000001_01010101_1;
      patterns[38084] = 25'b10010100_11000010_01010110_1;
      patterns[38085] = 25'b10010100_11000011_01010111_1;
      patterns[38086] = 25'b10010100_11000100_01011000_1;
      patterns[38087] = 25'b10010100_11000101_01011001_1;
      patterns[38088] = 25'b10010100_11000110_01011010_1;
      patterns[38089] = 25'b10010100_11000111_01011011_1;
      patterns[38090] = 25'b10010100_11001000_01011100_1;
      patterns[38091] = 25'b10010100_11001001_01011101_1;
      patterns[38092] = 25'b10010100_11001010_01011110_1;
      patterns[38093] = 25'b10010100_11001011_01011111_1;
      patterns[38094] = 25'b10010100_11001100_01100000_1;
      patterns[38095] = 25'b10010100_11001101_01100001_1;
      patterns[38096] = 25'b10010100_11001110_01100010_1;
      patterns[38097] = 25'b10010100_11001111_01100011_1;
      patterns[38098] = 25'b10010100_11010000_01100100_1;
      patterns[38099] = 25'b10010100_11010001_01100101_1;
      patterns[38100] = 25'b10010100_11010010_01100110_1;
      patterns[38101] = 25'b10010100_11010011_01100111_1;
      patterns[38102] = 25'b10010100_11010100_01101000_1;
      patterns[38103] = 25'b10010100_11010101_01101001_1;
      patterns[38104] = 25'b10010100_11010110_01101010_1;
      patterns[38105] = 25'b10010100_11010111_01101011_1;
      patterns[38106] = 25'b10010100_11011000_01101100_1;
      patterns[38107] = 25'b10010100_11011001_01101101_1;
      patterns[38108] = 25'b10010100_11011010_01101110_1;
      patterns[38109] = 25'b10010100_11011011_01101111_1;
      patterns[38110] = 25'b10010100_11011100_01110000_1;
      patterns[38111] = 25'b10010100_11011101_01110001_1;
      patterns[38112] = 25'b10010100_11011110_01110010_1;
      patterns[38113] = 25'b10010100_11011111_01110011_1;
      patterns[38114] = 25'b10010100_11100000_01110100_1;
      patterns[38115] = 25'b10010100_11100001_01110101_1;
      patterns[38116] = 25'b10010100_11100010_01110110_1;
      patterns[38117] = 25'b10010100_11100011_01110111_1;
      patterns[38118] = 25'b10010100_11100100_01111000_1;
      patterns[38119] = 25'b10010100_11100101_01111001_1;
      patterns[38120] = 25'b10010100_11100110_01111010_1;
      patterns[38121] = 25'b10010100_11100111_01111011_1;
      patterns[38122] = 25'b10010100_11101000_01111100_1;
      patterns[38123] = 25'b10010100_11101001_01111101_1;
      patterns[38124] = 25'b10010100_11101010_01111110_1;
      patterns[38125] = 25'b10010100_11101011_01111111_1;
      patterns[38126] = 25'b10010100_11101100_10000000_1;
      patterns[38127] = 25'b10010100_11101101_10000001_1;
      patterns[38128] = 25'b10010100_11101110_10000010_1;
      patterns[38129] = 25'b10010100_11101111_10000011_1;
      patterns[38130] = 25'b10010100_11110000_10000100_1;
      patterns[38131] = 25'b10010100_11110001_10000101_1;
      patterns[38132] = 25'b10010100_11110010_10000110_1;
      patterns[38133] = 25'b10010100_11110011_10000111_1;
      patterns[38134] = 25'b10010100_11110100_10001000_1;
      patterns[38135] = 25'b10010100_11110101_10001001_1;
      patterns[38136] = 25'b10010100_11110110_10001010_1;
      patterns[38137] = 25'b10010100_11110111_10001011_1;
      patterns[38138] = 25'b10010100_11111000_10001100_1;
      patterns[38139] = 25'b10010100_11111001_10001101_1;
      patterns[38140] = 25'b10010100_11111010_10001110_1;
      patterns[38141] = 25'b10010100_11111011_10001111_1;
      patterns[38142] = 25'b10010100_11111100_10010000_1;
      patterns[38143] = 25'b10010100_11111101_10010001_1;
      patterns[38144] = 25'b10010100_11111110_10010010_1;
      patterns[38145] = 25'b10010100_11111111_10010011_1;
      patterns[38146] = 25'b10010101_00000000_10010101_0;
      patterns[38147] = 25'b10010101_00000001_10010110_0;
      patterns[38148] = 25'b10010101_00000010_10010111_0;
      patterns[38149] = 25'b10010101_00000011_10011000_0;
      patterns[38150] = 25'b10010101_00000100_10011001_0;
      patterns[38151] = 25'b10010101_00000101_10011010_0;
      patterns[38152] = 25'b10010101_00000110_10011011_0;
      patterns[38153] = 25'b10010101_00000111_10011100_0;
      patterns[38154] = 25'b10010101_00001000_10011101_0;
      patterns[38155] = 25'b10010101_00001001_10011110_0;
      patterns[38156] = 25'b10010101_00001010_10011111_0;
      patterns[38157] = 25'b10010101_00001011_10100000_0;
      patterns[38158] = 25'b10010101_00001100_10100001_0;
      patterns[38159] = 25'b10010101_00001101_10100010_0;
      patterns[38160] = 25'b10010101_00001110_10100011_0;
      patterns[38161] = 25'b10010101_00001111_10100100_0;
      patterns[38162] = 25'b10010101_00010000_10100101_0;
      patterns[38163] = 25'b10010101_00010001_10100110_0;
      patterns[38164] = 25'b10010101_00010010_10100111_0;
      patterns[38165] = 25'b10010101_00010011_10101000_0;
      patterns[38166] = 25'b10010101_00010100_10101001_0;
      patterns[38167] = 25'b10010101_00010101_10101010_0;
      patterns[38168] = 25'b10010101_00010110_10101011_0;
      patterns[38169] = 25'b10010101_00010111_10101100_0;
      patterns[38170] = 25'b10010101_00011000_10101101_0;
      patterns[38171] = 25'b10010101_00011001_10101110_0;
      patterns[38172] = 25'b10010101_00011010_10101111_0;
      patterns[38173] = 25'b10010101_00011011_10110000_0;
      patterns[38174] = 25'b10010101_00011100_10110001_0;
      patterns[38175] = 25'b10010101_00011101_10110010_0;
      patterns[38176] = 25'b10010101_00011110_10110011_0;
      patterns[38177] = 25'b10010101_00011111_10110100_0;
      patterns[38178] = 25'b10010101_00100000_10110101_0;
      patterns[38179] = 25'b10010101_00100001_10110110_0;
      patterns[38180] = 25'b10010101_00100010_10110111_0;
      patterns[38181] = 25'b10010101_00100011_10111000_0;
      patterns[38182] = 25'b10010101_00100100_10111001_0;
      patterns[38183] = 25'b10010101_00100101_10111010_0;
      patterns[38184] = 25'b10010101_00100110_10111011_0;
      patterns[38185] = 25'b10010101_00100111_10111100_0;
      patterns[38186] = 25'b10010101_00101000_10111101_0;
      patterns[38187] = 25'b10010101_00101001_10111110_0;
      patterns[38188] = 25'b10010101_00101010_10111111_0;
      patterns[38189] = 25'b10010101_00101011_11000000_0;
      patterns[38190] = 25'b10010101_00101100_11000001_0;
      patterns[38191] = 25'b10010101_00101101_11000010_0;
      patterns[38192] = 25'b10010101_00101110_11000011_0;
      patterns[38193] = 25'b10010101_00101111_11000100_0;
      patterns[38194] = 25'b10010101_00110000_11000101_0;
      patterns[38195] = 25'b10010101_00110001_11000110_0;
      patterns[38196] = 25'b10010101_00110010_11000111_0;
      patterns[38197] = 25'b10010101_00110011_11001000_0;
      patterns[38198] = 25'b10010101_00110100_11001001_0;
      patterns[38199] = 25'b10010101_00110101_11001010_0;
      patterns[38200] = 25'b10010101_00110110_11001011_0;
      patterns[38201] = 25'b10010101_00110111_11001100_0;
      patterns[38202] = 25'b10010101_00111000_11001101_0;
      patterns[38203] = 25'b10010101_00111001_11001110_0;
      patterns[38204] = 25'b10010101_00111010_11001111_0;
      patterns[38205] = 25'b10010101_00111011_11010000_0;
      patterns[38206] = 25'b10010101_00111100_11010001_0;
      patterns[38207] = 25'b10010101_00111101_11010010_0;
      patterns[38208] = 25'b10010101_00111110_11010011_0;
      patterns[38209] = 25'b10010101_00111111_11010100_0;
      patterns[38210] = 25'b10010101_01000000_11010101_0;
      patterns[38211] = 25'b10010101_01000001_11010110_0;
      patterns[38212] = 25'b10010101_01000010_11010111_0;
      patterns[38213] = 25'b10010101_01000011_11011000_0;
      patterns[38214] = 25'b10010101_01000100_11011001_0;
      patterns[38215] = 25'b10010101_01000101_11011010_0;
      patterns[38216] = 25'b10010101_01000110_11011011_0;
      patterns[38217] = 25'b10010101_01000111_11011100_0;
      patterns[38218] = 25'b10010101_01001000_11011101_0;
      patterns[38219] = 25'b10010101_01001001_11011110_0;
      patterns[38220] = 25'b10010101_01001010_11011111_0;
      patterns[38221] = 25'b10010101_01001011_11100000_0;
      patterns[38222] = 25'b10010101_01001100_11100001_0;
      patterns[38223] = 25'b10010101_01001101_11100010_0;
      patterns[38224] = 25'b10010101_01001110_11100011_0;
      patterns[38225] = 25'b10010101_01001111_11100100_0;
      patterns[38226] = 25'b10010101_01010000_11100101_0;
      patterns[38227] = 25'b10010101_01010001_11100110_0;
      patterns[38228] = 25'b10010101_01010010_11100111_0;
      patterns[38229] = 25'b10010101_01010011_11101000_0;
      patterns[38230] = 25'b10010101_01010100_11101001_0;
      patterns[38231] = 25'b10010101_01010101_11101010_0;
      patterns[38232] = 25'b10010101_01010110_11101011_0;
      patterns[38233] = 25'b10010101_01010111_11101100_0;
      patterns[38234] = 25'b10010101_01011000_11101101_0;
      patterns[38235] = 25'b10010101_01011001_11101110_0;
      patterns[38236] = 25'b10010101_01011010_11101111_0;
      patterns[38237] = 25'b10010101_01011011_11110000_0;
      patterns[38238] = 25'b10010101_01011100_11110001_0;
      patterns[38239] = 25'b10010101_01011101_11110010_0;
      patterns[38240] = 25'b10010101_01011110_11110011_0;
      patterns[38241] = 25'b10010101_01011111_11110100_0;
      patterns[38242] = 25'b10010101_01100000_11110101_0;
      patterns[38243] = 25'b10010101_01100001_11110110_0;
      patterns[38244] = 25'b10010101_01100010_11110111_0;
      patterns[38245] = 25'b10010101_01100011_11111000_0;
      patterns[38246] = 25'b10010101_01100100_11111001_0;
      patterns[38247] = 25'b10010101_01100101_11111010_0;
      patterns[38248] = 25'b10010101_01100110_11111011_0;
      patterns[38249] = 25'b10010101_01100111_11111100_0;
      patterns[38250] = 25'b10010101_01101000_11111101_0;
      patterns[38251] = 25'b10010101_01101001_11111110_0;
      patterns[38252] = 25'b10010101_01101010_11111111_0;
      patterns[38253] = 25'b10010101_01101011_00000000_1;
      patterns[38254] = 25'b10010101_01101100_00000001_1;
      patterns[38255] = 25'b10010101_01101101_00000010_1;
      patterns[38256] = 25'b10010101_01101110_00000011_1;
      patterns[38257] = 25'b10010101_01101111_00000100_1;
      patterns[38258] = 25'b10010101_01110000_00000101_1;
      patterns[38259] = 25'b10010101_01110001_00000110_1;
      patterns[38260] = 25'b10010101_01110010_00000111_1;
      patterns[38261] = 25'b10010101_01110011_00001000_1;
      patterns[38262] = 25'b10010101_01110100_00001001_1;
      patterns[38263] = 25'b10010101_01110101_00001010_1;
      patterns[38264] = 25'b10010101_01110110_00001011_1;
      patterns[38265] = 25'b10010101_01110111_00001100_1;
      patterns[38266] = 25'b10010101_01111000_00001101_1;
      patterns[38267] = 25'b10010101_01111001_00001110_1;
      patterns[38268] = 25'b10010101_01111010_00001111_1;
      patterns[38269] = 25'b10010101_01111011_00010000_1;
      patterns[38270] = 25'b10010101_01111100_00010001_1;
      patterns[38271] = 25'b10010101_01111101_00010010_1;
      patterns[38272] = 25'b10010101_01111110_00010011_1;
      patterns[38273] = 25'b10010101_01111111_00010100_1;
      patterns[38274] = 25'b10010101_10000000_00010101_1;
      patterns[38275] = 25'b10010101_10000001_00010110_1;
      patterns[38276] = 25'b10010101_10000010_00010111_1;
      patterns[38277] = 25'b10010101_10000011_00011000_1;
      patterns[38278] = 25'b10010101_10000100_00011001_1;
      patterns[38279] = 25'b10010101_10000101_00011010_1;
      patterns[38280] = 25'b10010101_10000110_00011011_1;
      patterns[38281] = 25'b10010101_10000111_00011100_1;
      patterns[38282] = 25'b10010101_10001000_00011101_1;
      patterns[38283] = 25'b10010101_10001001_00011110_1;
      patterns[38284] = 25'b10010101_10001010_00011111_1;
      patterns[38285] = 25'b10010101_10001011_00100000_1;
      patterns[38286] = 25'b10010101_10001100_00100001_1;
      patterns[38287] = 25'b10010101_10001101_00100010_1;
      patterns[38288] = 25'b10010101_10001110_00100011_1;
      patterns[38289] = 25'b10010101_10001111_00100100_1;
      patterns[38290] = 25'b10010101_10010000_00100101_1;
      patterns[38291] = 25'b10010101_10010001_00100110_1;
      patterns[38292] = 25'b10010101_10010010_00100111_1;
      patterns[38293] = 25'b10010101_10010011_00101000_1;
      patterns[38294] = 25'b10010101_10010100_00101001_1;
      patterns[38295] = 25'b10010101_10010101_00101010_1;
      patterns[38296] = 25'b10010101_10010110_00101011_1;
      patterns[38297] = 25'b10010101_10010111_00101100_1;
      patterns[38298] = 25'b10010101_10011000_00101101_1;
      patterns[38299] = 25'b10010101_10011001_00101110_1;
      patterns[38300] = 25'b10010101_10011010_00101111_1;
      patterns[38301] = 25'b10010101_10011011_00110000_1;
      patterns[38302] = 25'b10010101_10011100_00110001_1;
      patterns[38303] = 25'b10010101_10011101_00110010_1;
      patterns[38304] = 25'b10010101_10011110_00110011_1;
      patterns[38305] = 25'b10010101_10011111_00110100_1;
      patterns[38306] = 25'b10010101_10100000_00110101_1;
      patterns[38307] = 25'b10010101_10100001_00110110_1;
      patterns[38308] = 25'b10010101_10100010_00110111_1;
      patterns[38309] = 25'b10010101_10100011_00111000_1;
      patterns[38310] = 25'b10010101_10100100_00111001_1;
      patterns[38311] = 25'b10010101_10100101_00111010_1;
      patterns[38312] = 25'b10010101_10100110_00111011_1;
      patterns[38313] = 25'b10010101_10100111_00111100_1;
      patterns[38314] = 25'b10010101_10101000_00111101_1;
      patterns[38315] = 25'b10010101_10101001_00111110_1;
      patterns[38316] = 25'b10010101_10101010_00111111_1;
      patterns[38317] = 25'b10010101_10101011_01000000_1;
      patterns[38318] = 25'b10010101_10101100_01000001_1;
      patterns[38319] = 25'b10010101_10101101_01000010_1;
      patterns[38320] = 25'b10010101_10101110_01000011_1;
      patterns[38321] = 25'b10010101_10101111_01000100_1;
      patterns[38322] = 25'b10010101_10110000_01000101_1;
      patterns[38323] = 25'b10010101_10110001_01000110_1;
      patterns[38324] = 25'b10010101_10110010_01000111_1;
      patterns[38325] = 25'b10010101_10110011_01001000_1;
      patterns[38326] = 25'b10010101_10110100_01001001_1;
      patterns[38327] = 25'b10010101_10110101_01001010_1;
      patterns[38328] = 25'b10010101_10110110_01001011_1;
      patterns[38329] = 25'b10010101_10110111_01001100_1;
      patterns[38330] = 25'b10010101_10111000_01001101_1;
      patterns[38331] = 25'b10010101_10111001_01001110_1;
      patterns[38332] = 25'b10010101_10111010_01001111_1;
      patterns[38333] = 25'b10010101_10111011_01010000_1;
      patterns[38334] = 25'b10010101_10111100_01010001_1;
      patterns[38335] = 25'b10010101_10111101_01010010_1;
      patterns[38336] = 25'b10010101_10111110_01010011_1;
      patterns[38337] = 25'b10010101_10111111_01010100_1;
      patterns[38338] = 25'b10010101_11000000_01010101_1;
      patterns[38339] = 25'b10010101_11000001_01010110_1;
      patterns[38340] = 25'b10010101_11000010_01010111_1;
      patterns[38341] = 25'b10010101_11000011_01011000_1;
      patterns[38342] = 25'b10010101_11000100_01011001_1;
      patterns[38343] = 25'b10010101_11000101_01011010_1;
      patterns[38344] = 25'b10010101_11000110_01011011_1;
      patterns[38345] = 25'b10010101_11000111_01011100_1;
      patterns[38346] = 25'b10010101_11001000_01011101_1;
      patterns[38347] = 25'b10010101_11001001_01011110_1;
      patterns[38348] = 25'b10010101_11001010_01011111_1;
      patterns[38349] = 25'b10010101_11001011_01100000_1;
      patterns[38350] = 25'b10010101_11001100_01100001_1;
      patterns[38351] = 25'b10010101_11001101_01100010_1;
      patterns[38352] = 25'b10010101_11001110_01100011_1;
      patterns[38353] = 25'b10010101_11001111_01100100_1;
      patterns[38354] = 25'b10010101_11010000_01100101_1;
      patterns[38355] = 25'b10010101_11010001_01100110_1;
      patterns[38356] = 25'b10010101_11010010_01100111_1;
      patterns[38357] = 25'b10010101_11010011_01101000_1;
      patterns[38358] = 25'b10010101_11010100_01101001_1;
      patterns[38359] = 25'b10010101_11010101_01101010_1;
      patterns[38360] = 25'b10010101_11010110_01101011_1;
      patterns[38361] = 25'b10010101_11010111_01101100_1;
      patterns[38362] = 25'b10010101_11011000_01101101_1;
      patterns[38363] = 25'b10010101_11011001_01101110_1;
      patterns[38364] = 25'b10010101_11011010_01101111_1;
      patterns[38365] = 25'b10010101_11011011_01110000_1;
      patterns[38366] = 25'b10010101_11011100_01110001_1;
      patterns[38367] = 25'b10010101_11011101_01110010_1;
      patterns[38368] = 25'b10010101_11011110_01110011_1;
      patterns[38369] = 25'b10010101_11011111_01110100_1;
      patterns[38370] = 25'b10010101_11100000_01110101_1;
      patterns[38371] = 25'b10010101_11100001_01110110_1;
      patterns[38372] = 25'b10010101_11100010_01110111_1;
      patterns[38373] = 25'b10010101_11100011_01111000_1;
      patterns[38374] = 25'b10010101_11100100_01111001_1;
      patterns[38375] = 25'b10010101_11100101_01111010_1;
      patterns[38376] = 25'b10010101_11100110_01111011_1;
      patterns[38377] = 25'b10010101_11100111_01111100_1;
      patterns[38378] = 25'b10010101_11101000_01111101_1;
      patterns[38379] = 25'b10010101_11101001_01111110_1;
      patterns[38380] = 25'b10010101_11101010_01111111_1;
      patterns[38381] = 25'b10010101_11101011_10000000_1;
      patterns[38382] = 25'b10010101_11101100_10000001_1;
      patterns[38383] = 25'b10010101_11101101_10000010_1;
      patterns[38384] = 25'b10010101_11101110_10000011_1;
      patterns[38385] = 25'b10010101_11101111_10000100_1;
      patterns[38386] = 25'b10010101_11110000_10000101_1;
      patterns[38387] = 25'b10010101_11110001_10000110_1;
      patterns[38388] = 25'b10010101_11110010_10000111_1;
      patterns[38389] = 25'b10010101_11110011_10001000_1;
      patterns[38390] = 25'b10010101_11110100_10001001_1;
      patterns[38391] = 25'b10010101_11110101_10001010_1;
      patterns[38392] = 25'b10010101_11110110_10001011_1;
      patterns[38393] = 25'b10010101_11110111_10001100_1;
      patterns[38394] = 25'b10010101_11111000_10001101_1;
      patterns[38395] = 25'b10010101_11111001_10001110_1;
      patterns[38396] = 25'b10010101_11111010_10001111_1;
      patterns[38397] = 25'b10010101_11111011_10010000_1;
      patterns[38398] = 25'b10010101_11111100_10010001_1;
      patterns[38399] = 25'b10010101_11111101_10010010_1;
      patterns[38400] = 25'b10010101_11111110_10010011_1;
      patterns[38401] = 25'b10010101_11111111_10010100_1;
      patterns[38402] = 25'b10010110_00000000_10010110_0;
      patterns[38403] = 25'b10010110_00000001_10010111_0;
      patterns[38404] = 25'b10010110_00000010_10011000_0;
      patterns[38405] = 25'b10010110_00000011_10011001_0;
      patterns[38406] = 25'b10010110_00000100_10011010_0;
      patterns[38407] = 25'b10010110_00000101_10011011_0;
      patterns[38408] = 25'b10010110_00000110_10011100_0;
      patterns[38409] = 25'b10010110_00000111_10011101_0;
      patterns[38410] = 25'b10010110_00001000_10011110_0;
      patterns[38411] = 25'b10010110_00001001_10011111_0;
      patterns[38412] = 25'b10010110_00001010_10100000_0;
      patterns[38413] = 25'b10010110_00001011_10100001_0;
      patterns[38414] = 25'b10010110_00001100_10100010_0;
      patterns[38415] = 25'b10010110_00001101_10100011_0;
      patterns[38416] = 25'b10010110_00001110_10100100_0;
      patterns[38417] = 25'b10010110_00001111_10100101_0;
      patterns[38418] = 25'b10010110_00010000_10100110_0;
      patterns[38419] = 25'b10010110_00010001_10100111_0;
      patterns[38420] = 25'b10010110_00010010_10101000_0;
      patterns[38421] = 25'b10010110_00010011_10101001_0;
      patterns[38422] = 25'b10010110_00010100_10101010_0;
      patterns[38423] = 25'b10010110_00010101_10101011_0;
      patterns[38424] = 25'b10010110_00010110_10101100_0;
      patterns[38425] = 25'b10010110_00010111_10101101_0;
      patterns[38426] = 25'b10010110_00011000_10101110_0;
      patterns[38427] = 25'b10010110_00011001_10101111_0;
      patterns[38428] = 25'b10010110_00011010_10110000_0;
      patterns[38429] = 25'b10010110_00011011_10110001_0;
      patterns[38430] = 25'b10010110_00011100_10110010_0;
      patterns[38431] = 25'b10010110_00011101_10110011_0;
      patterns[38432] = 25'b10010110_00011110_10110100_0;
      patterns[38433] = 25'b10010110_00011111_10110101_0;
      patterns[38434] = 25'b10010110_00100000_10110110_0;
      patterns[38435] = 25'b10010110_00100001_10110111_0;
      patterns[38436] = 25'b10010110_00100010_10111000_0;
      patterns[38437] = 25'b10010110_00100011_10111001_0;
      patterns[38438] = 25'b10010110_00100100_10111010_0;
      patterns[38439] = 25'b10010110_00100101_10111011_0;
      patterns[38440] = 25'b10010110_00100110_10111100_0;
      patterns[38441] = 25'b10010110_00100111_10111101_0;
      patterns[38442] = 25'b10010110_00101000_10111110_0;
      patterns[38443] = 25'b10010110_00101001_10111111_0;
      patterns[38444] = 25'b10010110_00101010_11000000_0;
      patterns[38445] = 25'b10010110_00101011_11000001_0;
      patterns[38446] = 25'b10010110_00101100_11000010_0;
      patterns[38447] = 25'b10010110_00101101_11000011_0;
      patterns[38448] = 25'b10010110_00101110_11000100_0;
      patterns[38449] = 25'b10010110_00101111_11000101_0;
      patterns[38450] = 25'b10010110_00110000_11000110_0;
      patterns[38451] = 25'b10010110_00110001_11000111_0;
      patterns[38452] = 25'b10010110_00110010_11001000_0;
      patterns[38453] = 25'b10010110_00110011_11001001_0;
      patterns[38454] = 25'b10010110_00110100_11001010_0;
      patterns[38455] = 25'b10010110_00110101_11001011_0;
      patterns[38456] = 25'b10010110_00110110_11001100_0;
      patterns[38457] = 25'b10010110_00110111_11001101_0;
      patterns[38458] = 25'b10010110_00111000_11001110_0;
      patterns[38459] = 25'b10010110_00111001_11001111_0;
      patterns[38460] = 25'b10010110_00111010_11010000_0;
      patterns[38461] = 25'b10010110_00111011_11010001_0;
      patterns[38462] = 25'b10010110_00111100_11010010_0;
      patterns[38463] = 25'b10010110_00111101_11010011_0;
      patterns[38464] = 25'b10010110_00111110_11010100_0;
      patterns[38465] = 25'b10010110_00111111_11010101_0;
      patterns[38466] = 25'b10010110_01000000_11010110_0;
      patterns[38467] = 25'b10010110_01000001_11010111_0;
      patterns[38468] = 25'b10010110_01000010_11011000_0;
      patterns[38469] = 25'b10010110_01000011_11011001_0;
      patterns[38470] = 25'b10010110_01000100_11011010_0;
      patterns[38471] = 25'b10010110_01000101_11011011_0;
      patterns[38472] = 25'b10010110_01000110_11011100_0;
      patterns[38473] = 25'b10010110_01000111_11011101_0;
      patterns[38474] = 25'b10010110_01001000_11011110_0;
      patterns[38475] = 25'b10010110_01001001_11011111_0;
      patterns[38476] = 25'b10010110_01001010_11100000_0;
      patterns[38477] = 25'b10010110_01001011_11100001_0;
      patterns[38478] = 25'b10010110_01001100_11100010_0;
      patterns[38479] = 25'b10010110_01001101_11100011_0;
      patterns[38480] = 25'b10010110_01001110_11100100_0;
      patterns[38481] = 25'b10010110_01001111_11100101_0;
      patterns[38482] = 25'b10010110_01010000_11100110_0;
      patterns[38483] = 25'b10010110_01010001_11100111_0;
      patterns[38484] = 25'b10010110_01010010_11101000_0;
      patterns[38485] = 25'b10010110_01010011_11101001_0;
      patterns[38486] = 25'b10010110_01010100_11101010_0;
      patterns[38487] = 25'b10010110_01010101_11101011_0;
      patterns[38488] = 25'b10010110_01010110_11101100_0;
      patterns[38489] = 25'b10010110_01010111_11101101_0;
      patterns[38490] = 25'b10010110_01011000_11101110_0;
      patterns[38491] = 25'b10010110_01011001_11101111_0;
      patterns[38492] = 25'b10010110_01011010_11110000_0;
      patterns[38493] = 25'b10010110_01011011_11110001_0;
      patterns[38494] = 25'b10010110_01011100_11110010_0;
      patterns[38495] = 25'b10010110_01011101_11110011_0;
      patterns[38496] = 25'b10010110_01011110_11110100_0;
      patterns[38497] = 25'b10010110_01011111_11110101_0;
      patterns[38498] = 25'b10010110_01100000_11110110_0;
      patterns[38499] = 25'b10010110_01100001_11110111_0;
      patterns[38500] = 25'b10010110_01100010_11111000_0;
      patterns[38501] = 25'b10010110_01100011_11111001_0;
      patterns[38502] = 25'b10010110_01100100_11111010_0;
      patterns[38503] = 25'b10010110_01100101_11111011_0;
      patterns[38504] = 25'b10010110_01100110_11111100_0;
      patterns[38505] = 25'b10010110_01100111_11111101_0;
      patterns[38506] = 25'b10010110_01101000_11111110_0;
      patterns[38507] = 25'b10010110_01101001_11111111_0;
      patterns[38508] = 25'b10010110_01101010_00000000_1;
      patterns[38509] = 25'b10010110_01101011_00000001_1;
      patterns[38510] = 25'b10010110_01101100_00000010_1;
      patterns[38511] = 25'b10010110_01101101_00000011_1;
      patterns[38512] = 25'b10010110_01101110_00000100_1;
      patterns[38513] = 25'b10010110_01101111_00000101_1;
      patterns[38514] = 25'b10010110_01110000_00000110_1;
      patterns[38515] = 25'b10010110_01110001_00000111_1;
      patterns[38516] = 25'b10010110_01110010_00001000_1;
      patterns[38517] = 25'b10010110_01110011_00001001_1;
      patterns[38518] = 25'b10010110_01110100_00001010_1;
      patterns[38519] = 25'b10010110_01110101_00001011_1;
      patterns[38520] = 25'b10010110_01110110_00001100_1;
      patterns[38521] = 25'b10010110_01110111_00001101_1;
      patterns[38522] = 25'b10010110_01111000_00001110_1;
      patterns[38523] = 25'b10010110_01111001_00001111_1;
      patterns[38524] = 25'b10010110_01111010_00010000_1;
      patterns[38525] = 25'b10010110_01111011_00010001_1;
      patterns[38526] = 25'b10010110_01111100_00010010_1;
      patterns[38527] = 25'b10010110_01111101_00010011_1;
      patterns[38528] = 25'b10010110_01111110_00010100_1;
      patterns[38529] = 25'b10010110_01111111_00010101_1;
      patterns[38530] = 25'b10010110_10000000_00010110_1;
      patterns[38531] = 25'b10010110_10000001_00010111_1;
      patterns[38532] = 25'b10010110_10000010_00011000_1;
      patterns[38533] = 25'b10010110_10000011_00011001_1;
      patterns[38534] = 25'b10010110_10000100_00011010_1;
      patterns[38535] = 25'b10010110_10000101_00011011_1;
      patterns[38536] = 25'b10010110_10000110_00011100_1;
      patterns[38537] = 25'b10010110_10000111_00011101_1;
      patterns[38538] = 25'b10010110_10001000_00011110_1;
      patterns[38539] = 25'b10010110_10001001_00011111_1;
      patterns[38540] = 25'b10010110_10001010_00100000_1;
      patterns[38541] = 25'b10010110_10001011_00100001_1;
      patterns[38542] = 25'b10010110_10001100_00100010_1;
      patterns[38543] = 25'b10010110_10001101_00100011_1;
      patterns[38544] = 25'b10010110_10001110_00100100_1;
      patterns[38545] = 25'b10010110_10001111_00100101_1;
      patterns[38546] = 25'b10010110_10010000_00100110_1;
      patterns[38547] = 25'b10010110_10010001_00100111_1;
      patterns[38548] = 25'b10010110_10010010_00101000_1;
      patterns[38549] = 25'b10010110_10010011_00101001_1;
      patterns[38550] = 25'b10010110_10010100_00101010_1;
      patterns[38551] = 25'b10010110_10010101_00101011_1;
      patterns[38552] = 25'b10010110_10010110_00101100_1;
      patterns[38553] = 25'b10010110_10010111_00101101_1;
      patterns[38554] = 25'b10010110_10011000_00101110_1;
      patterns[38555] = 25'b10010110_10011001_00101111_1;
      patterns[38556] = 25'b10010110_10011010_00110000_1;
      patterns[38557] = 25'b10010110_10011011_00110001_1;
      patterns[38558] = 25'b10010110_10011100_00110010_1;
      patterns[38559] = 25'b10010110_10011101_00110011_1;
      patterns[38560] = 25'b10010110_10011110_00110100_1;
      patterns[38561] = 25'b10010110_10011111_00110101_1;
      patterns[38562] = 25'b10010110_10100000_00110110_1;
      patterns[38563] = 25'b10010110_10100001_00110111_1;
      patterns[38564] = 25'b10010110_10100010_00111000_1;
      patterns[38565] = 25'b10010110_10100011_00111001_1;
      patterns[38566] = 25'b10010110_10100100_00111010_1;
      patterns[38567] = 25'b10010110_10100101_00111011_1;
      patterns[38568] = 25'b10010110_10100110_00111100_1;
      patterns[38569] = 25'b10010110_10100111_00111101_1;
      patterns[38570] = 25'b10010110_10101000_00111110_1;
      patterns[38571] = 25'b10010110_10101001_00111111_1;
      patterns[38572] = 25'b10010110_10101010_01000000_1;
      patterns[38573] = 25'b10010110_10101011_01000001_1;
      patterns[38574] = 25'b10010110_10101100_01000010_1;
      patterns[38575] = 25'b10010110_10101101_01000011_1;
      patterns[38576] = 25'b10010110_10101110_01000100_1;
      patterns[38577] = 25'b10010110_10101111_01000101_1;
      patterns[38578] = 25'b10010110_10110000_01000110_1;
      patterns[38579] = 25'b10010110_10110001_01000111_1;
      patterns[38580] = 25'b10010110_10110010_01001000_1;
      patterns[38581] = 25'b10010110_10110011_01001001_1;
      patterns[38582] = 25'b10010110_10110100_01001010_1;
      patterns[38583] = 25'b10010110_10110101_01001011_1;
      patterns[38584] = 25'b10010110_10110110_01001100_1;
      patterns[38585] = 25'b10010110_10110111_01001101_1;
      patterns[38586] = 25'b10010110_10111000_01001110_1;
      patterns[38587] = 25'b10010110_10111001_01001111_1;
      patterns[38588] = 25'b10010110_10111010_01010000_1;
      patterns[38589] = 25'b10010110_10111011_01010001_1;
      patterns[38590] = 25'b10010110_10111100_01010010_1;
      patterns[38591] = 25'b10010110_10111101_01010011_1;
      patterns[38592] = 25'b10010110_10111110_01010100_1;
      patterns[38593] = 25'b10010110_10111111_01010101_1;
      patterns[38594] = 25'b10010110_11000000_01010110_1;
      patterns[38595] = 25'b10010110_11000001_01010111_1;
      patterns[38596] = 25'b10010110_11000010_01011000_1;
      patterns[38597] = 25'b10010110_11000011_01011001_1;
      patterns[38598] = 25'b10010110_11000100_01011010_1;
      patterns[38599] = 25'b10010110_11000101_01011011_1;
      patterns[38600] = 25'b10010110_11000110_01011100_1;
      patterns[38601] = 25'b10010110_11000111_01011101_1;
      patterns[38602] = 25'b10010110_11001000_01011110_1;
      patterns[38603] = 25'b10010110_11001001_01011111_1;
      patterns[38604] = 25'b10010110_11001010_01100000_1;
      patterns[38605] = 25'b10010110_11001011_01100001_1;
      patterns[38606] = 25'b10010110_11001100_01100010_1;
      patterns[38607] = 25'b10010110_11001101_01100011_1;
      patterns[38608] = 25'b10010110_11001110_01100100_1;
      patterns[38609] = 25'b10010110_11001111_01100101_1;
      patterns[38610] = 25'b10010110_11010000_01100110_1;
      patterns[38611] = 25'b10010110_11010001_01100111_1;
      patterns[38612] = 25'b10010110_11010010_01101000_1;
      patterns[38613] = 25'b10010110_11010011_01101001_1;
      patterns[38614] = 25'b10010110_11010100_01101010_1;
      patterns[38615] = 25'b10010110_11010101_01101011_1;
      patterns[38616] = 25'b10010110_11010110_01101100_1;
      patterns[38617] = 25'b10010110_11010111_01101101_1;
      patterns[38618] = 25'b10010110_11011000_01101110_1;
      patterns[38619] = 25'b10010110_11011001_01101111_1;
      patterns[38620] = 25'b10010110_11011010_01110000_1;
      patterns[38621] = 25'b10010110_11011011_01110001_1;
      patterns[38622] = 25'b10010110_11011100_01110010_1;
      patterns[38623] = 25'b10010110_11011101_01110011_1;
      patterns[38624] = 25'b10010110_11011110_01110100_1;
      patterns[38625] = 25'b10010110_11011111_01110101_1;
      patterns[38626] = 25'b10010110_11100000_01110110_1;
      patterns[38627] = 25'b10010110_11100001_01110111_1;
      patterns[38628] = 25'b10010110_11100010_01111000_1;
      patterns[38629] = 25'b10010110_11100011_01111001_1;
      patterns[38630] = 25'b10010110_11100100_01111010_1;
      patterns[38631] = 25'b10010110_11100101_01111011_1;
      patterns[38632] = 25'b10010110_11100110_01111100_1;
      patterns[38633] = 25'b10010110_11100111_01111101_1;
      patterns[38634] = 25'b10010110_11101000_01111110_1;
      patterns[38635] = 25'b10010110_11101001_01111111_1;
      patterns[38636] = 25'b10010110_11101010_10000000_1;
      patterns[38637] = 25'b10010110_11101011_10000001_1;
      patterns[38638] = 25'b10010110_11101100_10000010_1;
      patterns[38639] = 25'b10010110_11101101_10000011_1;
      patterns[38640] = 25'b10010110_11101110_10000100_1;
      patterns[38641] = 25'b10010110_11101111_10000101_1;
      patterns[38642] = 25'b10010110_11110000_10000110_1;
      patterns[38643] = 25'b10010110_11110001_10000111_1;
      patterns[38644] = 25'b10010110_11110010_10001000_1;
      patterns[38645] = 25'b10010110_11110011_10001001_1;
      patterns[38646] = 25'b10010110_11110100_10001010_1;
      patterns[38647] = 25'b10010110_11110101_10001011_1;
      patterns[38648] = 25'b10010110_11110110_10001100_1;
      patterns[38649] = 25'b10010110_11110111_10001101_1;
      patterns[38650] = 25'b10010110_11111000_10001110_1;
      patterns[38651] = 25'b10010110_11111001_10001111_1;
      patterns[38652] = 25'b10010110_11111010_10010000_1;
      patterns[38653] = 25'b10010110_11111011_10010001_1;
      patterns[38654] = 25'b10010110_11111100_10010010_1;
      patterns[38655] = 25'b10010110_11111101_10010011_1;
      patterns[38656] = 25'b10010110_11111110_10010100_1;
      patterns[38657] = 25'b10010110_11111111_10010101_1;
      patterns[38658] = 25'b10010111_00000000_10010111_0;
      patterns[38659] = 25'b10010111_00000001_10011000_0;
      patterns[38660] = 25'b10010111_00000010_10011001_0;
      patterns[38661] = 25'b10010111_00000011_10011010_0;
      patterns[38662] = 25'b10010111_00000100_10011011_0;
      patterns[38663] = 25'b10010111_00000101_10011100_0;
      patterns[38664] = 25'b10010111_00000110_10011101_0;
      patterns[38665] = 25'b10010111_00000111_10011110_0;
      patterns[38666] = 25'b10010111_00001000_10011111_0;
      patterns[38667] = 25'b10010111_00001001_10100000_0;
      patterns[38668] = 25'b10010111_00001010_10100001_0;
      patterns[38669] = 25'b10010111_00001011_10100010_0;
      patterns[38670] = 25'b10010111_00001100_10100011_0;
      patterns[38671] = 25'b10010111_00001101_10100100_0;
      patterns[38672] = 25'b10010111_00001110_10100101_0;
      patterns[38673] = 25'b10010111_00001111_10100110_0;
      patterns[38674] = 25'b10010111_00010000_10100111_0;
      patterns[38675] = 25'b10010111_00010001_10101000_0;
      patterns[38676] = 25'b10010111_00010010_10101001_0;
      patterns[38677] = 25'b10010111_00010011_10101010_0;
      patterns[38678] = 25'b10010111_00010100_10101011_0;
      patterns[38679] = 25'b10010111_00010101_10101100_0;
      patterns[38680] = 25'b10010111_00010110_10101101_0;
      patterns[38681] = 25'b10010111_00010111_10101110_0;
      patterns[38682] = 25'b10010111_00011000_10101111_0;
      patterns[38683] = 25'b10010111_00011001_10110000_0;
      patterns[38684] = 25'b10010111_00011010_10110001_0;
      patterns[38685] = 25'b10010111_00011011_10110010_0;
      patterns[38686] = 25'b10010111_00011100_10110011_0;
      patterns[38687] = 25'b10010111_00011101_10110100_0;
      patterns[38688] = 25'b10010111_00011110_10110101_0;
      patterns[38689] = 25'b10010111_00011111_10110110_0;
      patterns[38690] = 25'b10010111_00100000_10110111_0;
      patterns[38691] = 25'b10010111_00100001_10111000_0;
      patterns[38692] = 25'b10010111_00100010_10111001_0;
      patterns[38693] = 25'b10010111_00100011_10111010_0;
      patterns[38694] = 25'b10010111_00100100_10111011_0;
      patterns[38695] = 25'b10010111_00100101_10111100_0;
      patterns[38696] = 25'b10010111_00100110_10111101_0;
      patterns[38697] = 25'b10010111_00100111_10111110_0;
      patterns[38698] = 25'b10010111_00101000_10111111_0;
      patterns[38699] = 25'b10010111_00101001_11000000_0;
      patterns[38700] = 25'b10010111_00101010_11000001_0;
      patterns[38701] = 25'b10010111_00101011_11000010_0;
      patterns[38702] = 25'b10010111_00101100_11000011_0;
      patterns[38703] = 25'b10010111_00101101_11000100_0;
      patterns[38704] = 25'b10010111_00101110_11000101_0;
      patterns[38705] = 25'b10010111_00101111_11000110_0;
      patterns[38706] = 25'b10010111_00110000_11000111_0;
      patterns[38707] = 25'b10010111_00110001_11001000_0;
      patterns[38708] = 25'b10010111_00110010_11001001_0;
      patterns[38709] = 25'b10010111_00110011_11001010_0;
      patterns[38710] = 25'b10010111_00110100_11001011_0;
      patterns[38711] = 25'b10010111_00110101_11001100_0;
      patterns[38712] = 25'b10010111_00110110_11001101_0;
      patterns[38713] = 25'b10010111_00110111_11001110_0;
      patterns[38714] = 25'b10010111_00111000_11001111_0;
      patterns[38715] = 25'b10010111_00111001_11010000_0;
      patterns[38716] = 25'b10010111_00111010_11010001_0;
      patterns[38717] = 25'b10010111_00111011_11010010_0;
      patterns[38718] = 25'b10010111_00111100_11010011_0;
      patterns[38719] = 25'b10010111_00111101_11010100_0;
      patterns[38720] = 25'b10010111_00111110_11010101_0;
      patterns[38721] = 25'b10010111_00111111_11010110_0;
      patterns[38722] = 25'b10010111_01000000_11010111_0;
      patterns[38723] = 25'b10010111_01000001_11011000_0;
      patterns[38724] = 25'b10010111_01000010_11011001_0;
      patterns[38725] = 25'b10010111_01000011_11011010_0;
      patterns[38726] = 25'b10010111_01000100_11011011_0;
      patterns[38727] = 25'b10010111_01000101_11011100_0;
      patterns[38728] = 25'b10010111_01000110_11011101_0;
      patterns[38729] = 25'b10010111_01000111_11011110_0;
      patterns[38730] = 25'b10010111_01001000_11011111_0;
      patterns[38731] = 25'b10010111_01001001_11100000_0;
      patterns[38732] = 25'b10010111_01001010_11100001_0;
      patterns[38733] = 25'b10010111_01001011_11100010_0;
      patterns[38734] = 25'b10010111_01001100_11100011_0;
      patterns[38735] = 25'b10010111_01001101_11100100_0;
      patterns[38736] = 25'b10010111_01001110_11100101_0;
      patterns[38737] = 25'b10010111_01001111_11100110_0;
      patterns[38738] = 25'b10010111_01010000_11100111_0;
      patterns[38739] = 25'b10010111_01010001_11101000_0;
      patterns[38740] = 25'b10010111_01010010_11101001_0;
      patterns[38741] = 25'b10010111_01010011_11101010_0;
      patterns[38742] = 25'b10010111_01010100_11101011_0;
      patterns[38743] = 25'b10010111_01010101_11101100_0;
      patterns[38744] = 25'b10010111_01010110_11101101_0;
      patterns[38745] = 25'b10010111_01010111_11101110_0;
      patterns[38746] = 25'b10010111_01011000_11101111_0;
      patterns[38747] = 25'b10010111_01011001_11110000_0;
      patterns[38748] = 25'b10010111_01011010_11110001_0;
      patterns[38749] = 25'b10010111_01011011_11110010_0;
      patterns[38750] = 25'b10010111_01011100_11110011_0;
      patterns[38751] = 25'b10010111_01011101_11110100_0;
      patterns[38752] = 25'b10010111_01011110_11110101_0;
      patterns[38753] = 25'b10010111_01011111_11110110_0;
      patterns[38754] = 25'b10010111_01100000_11110111_0;
      patterns[38755] = 25'b10010111_01100001_11111000_0;
      patterns[38756] = 25'b10010111_01100010_11111001_0;
      patterns[38757] = 25'b10010111_01100011_11111010_0;
      patterns[38758] = 25'b10010111_01100100_11111011_0;
      patterns[38759] = 25'b10010111_01100101_11111100_0;
      patterns[38760] = 25'b10010111_01100110_11111101_0;
      patterns[38761] = 25'b10010111_01100111_11111110_0;
      patterns[38762] = 25'b10010111_01101000_11111111_0;
      patterns[38763] = 25'b10010111_01101001_00000000_1;
      patterns[38764] = 25'b10010111_01101010_00000001_1;
      patterns[38765] = 25'b10010111_01101011_00000010_1;
      patterns[38766] = 25'b10010111_01101100_00000011_1;
      patterns[38767] = 25'b10010111_01101101_00000100_1;
      patterns[38768] = 25'b10010111_01101110_00000101_1;
      patterns[38769] = 25'b10010111_01101111_00000110_1;
      patterns[38770] = 25'b10010111_01110000_00000111_1;
      patterns[38771] = 25'b10010111_01110001_00001000_1;
      patterns[38772] = 25'b10010111_01110010_00001001_1;
      patterns[38773] = 25'b10010111_01110011_00001010_1;
      patterns[38774] = 25'b10010111_01110100_00001011_1;
      patterns[38775] = 25'b10010111_01110101_00001100_1;
      patterns[38776] = 25'b10010111_01110110_00001101_1;
      patterns[38777] = 25'b10010111_01110111_00001110_1;
      patterns[38778] = 25'b10010111_01111000_00001111_1;
      patterns[38779] = 25'b10010111_01111001_00010000_1;
      patterns[38780] = 25'b10010111_01111010_00010001_1;
      patterns[38781] = 25'b10010111_01111011_00010010_1;
      patterns[38782] = 25'b10010111_01111100_00010011_1;
      patterns[38783] = 25'b10010111_01111101_00010100_1;
      patterns[38784] = 25'b10010111_01111110_00010101_1;
      patterns[38785] = 25'b10010111_01111111_00010110_1;
      patterns[38786] = 25'b10010111_10000000_00010111_1;
      patterns[38787] = 25'b10010111_10000001_00011000_1;
      patterns[38788] = 25'b10010111_10000010_00011001_1;
      patterns[38789] = 25'b10010111_10000011_00011010_1;
      patterns[38790] = 25'b10010111_10000100_00011011_1;
      patterns[38791] = 25'b10010111_10000101_00011100_1;
      patterns[38792] = 25'b10010111_10000110_00011101_1;
      patterns[38793] = 25'b10010111_10000111_00011110_1;
      patterns[38794] = 25'b10010111_10001000_00011111_1;
      patterns[38795] = 25'b10010111_10001001_00100000_1;
      patterns[38796] = 25'b10010111_10001010_00100001_1;
      patterns[38797] = 25'b10010111_10001011_00100010_1;
      patterns[38798] = 25'b10010111_10001100_00100011_1;
      patterns[38799] = 25'b10010111_10001101_00100100_1;
      patterns[38800] = 25'b10010111_10001110_00100101_1;
      patterns[38801] = 25'b10010111_10001111_00100110_1;
      patterns[38802] = 25'b10010111_10010000_00100111_1;
      patterns[38803] = 25'b10010111_10010001_00101000_1;
      patterns[38804] = 25'b10010111_10010010_00101001_1;
      patterns[38805] = 25'b10010111_10010011_00101010_1;
      patterns[38806] = 25'b10010111_10010100_00101011_1;
      patterns[38807] = 25'b10010111_10010101_00101100_1;
      patterns[38808] = 25'b10010111_10010110_00101101_1;
      patterns[38809] = 25'b10010111_10010111_00101110_1;
      patterns[38810] = 25'b10010111_10011000_00101111_1;
      patterns[38811] = 25'b10010111_10011001_00110000_1;
      patterns[38812] = 25'b10010111_10011010_00110001_1;
      patterns[38813] = 25'b10010111_10011011_00110010_1;
      patterns[38814] = 25'b10010111_10011100_00110011_1;
      patterns[38815] = 25'b10010111_10011101_00110100_1;
      patterns[38816] = 25'b10010111_10011110_00110101_1;
      patterns[38817] = 25'b10010111_10011111_00110110_1;
      patterns[38818] = 25'b10010111_10100000_00110111_1;
      patterns[38819] = 25'b10010111_10100001_00111000_1;
      patterns[38820] = 25'b10010111_10100010_00111001_1;
      patterns[38821] = 25'b10010111_10100011_00111010_1;
      patterns[38822] = 25'b10010111_10100100_00111011_1;
      patterns[38823] = 25'b10010111_10100101_00111100_1;
      patterns[38824] = 25'b10010111_10100110_00111101_1;
      patterns[38825] = 25'b10010111_10100111_00111110_1;
      patterns[38826] = 25'b10010111_10101000_00111111_1;
      patterns[38827] = 25'b10010111_10101001_01000000_1;
      patterns[38828] = 25'b10010111_10101010_01000001_1;
      patterns[38829] = 25'b10010111_10101011_01000010_1;
      patterns[38830] = 25'b10010111_10101100_01000011_1;
      patterns[38831] = 25'b10010111_10101101_01000100_1;
      patterns[38832] = 25'b10010111_10101110_01000101_1;
      patterns[38833] = 25'b10010111_10101111_01000110_1;
      patterns[38834] = 25'b10010111_10110000_01000111_1;
      patterns[38835] = 25'b10010111_10110001_01001000_1;
      patterns[38836] = 25'b10010111_10110010_01001001_1;
      patterns[38837] = 25'b10010111_10110011_01001010_1;
      patterns[38838] = 25'b10010111_10110100_01001011_1;
      patterns[38839] = 25'b10010111_10110101_01001100_1;
      patterns[38840] = 25'b10010111_10110110_01001101_1;
      patterns[38841] = 25'b10010111_10110111_01001110_1;
      patterns[38842] = 25'b10010111_10111000_01001111_1;
      patterns[38843] = 25'b10010111_10111001_01010000_1;
      patterns[38844] = 25'b10010111_10111010_01010001_1;
      patterns[38845] = 25'b10010111_10111011_01010010_1;
      patterns[38846] = 25'b10010111_10111100_01010011_1;
      patterns[38847] = 25'b10010111_10111101_01010100_1;
      patterns[38848] = 25'b10010111_10111110_01010101_1;
      patterns[38849] = 25'b10010111_10111111_01010110_1;
      patterns[38850] = 25'b10010111_11000000_01010111_1;
      patterns[38851] = 25'b10010111_11000001_01011000_1;
      patterns[38852] = 25'b10010111_11000010_01011001_1;
      patterns[38853] = 25'b10010111_11000011_01011010_1;
      patterns[38854] = 25'b10010111_11000100_01011011_1;
      patterns[38855] = 25'b10010111_11000101_01011100_1;
      patterns[38856] = 25'b10010111_11000110_01011101_1;
      patterns[38857] = 25'b10010111_11000111_01011110_1;
      patterns[38858] = 25'b10010111_11001000_01011111_1;
      patterns[38859] = 25'b10010111_11001001_01100000_1;
      patterns[38860] = 25'b10010111_11001010_01100001_1;
      patterns[38861] = 25'b10010111_11001011_01100010_1;
      patterns[38862] = 25'b10010111_11001100_01100011_1;
      patterns[38863] = 25'b10010111_11001101_01100100_1;
      patterns[38864] = 25'b10010111_11001110_01100101_1;
      patterns[38865] = 25'b10010111_11001111_01100110_1;
      patterns[38866] = 25'b10010111_11010000_01100111_1;
      patterns[38867] = 25'b10010111_11010001_01101000_1;
      patterns[38868] = 25'b10010111_11010010_01101001_1;
      patterns[38869] = 25'b10010111_11010011_01101010_1;
      patterns[38870] = 25'b10010111_11010100_01101011_1;
      patterns[38871] = 25'b10010111_11010101_01101100_1;
      patterns[38872] = 25'b10010111_11010110_01101101_1;
      patterns[38873] = 25'b10010111_11010111_01101110_1;
      patterns[38874] = 25'b10010111_11011000_01101111_1;
      patterns[38875] = 25'b10010111_11011001_01110000_1;
      patterns[38876] = 25'b10010111_11011010_01110001_1;
      patterns[38877] = 25'b10010111_11011011_01110010_1;
      patterns[38878] = 25'b10010111_11011100_01110011_1;
      patterns[38879] = 25'b10010111_11011101_01110100_1;
      patterns[38880] = 25'b10010111_11011110_01110101_1;
      patterns[38881] = 25'b10010111_11011111_01110110_1;
      patterns[38882] = 25'b10010111_11100000_01110111_1;
      patterns[38883] = 25'b10010111_11100001_01111000_1;
      patterns[38884] = 25'b10010111_11100010_01111001_1;
      patterns[38885] = 25'b10010111_11100011_01111010_1;
      patterns[38886] = 25'b10010111_11100100_01111011_1;
      patterns[38887] = 25'b10010111_11100101_01111100_1;
      patterns[38888] = 25'b10010111_11100110_01111101_1;
      patterns[38889] = 25'b10010111_11100111_01111110_1;
      patterns[38890] = 25'b10010111_11101000_01111111_1;
      patterns[38891] = 25'b10010111_11101001_10000000_1;
      patterns[38892] = 25'b10010111_11101010_10000001_1;
      patterns[38893] = 25'b10010111_11101011_10000010_1;
      patterns[38894] = 25'b10010111_11101100_10000011_1;
      patterns[38895] = 25'b10010111_11101101_10000100_1;
      patterns[38896] = 25'b10010111_11101110_10000101_1;
      patterns[38897] = 25'b10010111_11101111_10000110_1;
      patterns[38898] = 25'b10010111_11110000_10000111_1;
      patterns[38899] = 25'b10010111_11110001_10001000_1;
      patterns[38900] = 25'b10010111_11110010_10001001_1;
      patterns[38901] = 25'b10010111_11110011_10001010_1;
      patterns[38902] = 25'b10010111_11110100_10001011_1;
      patterns[38903] = 25'b10010111_11110101_10001100_1;
      patterns[38904] = 25'b10010111_11110110_10001101_1;
      patterns[38905] = 25'b10010111_11110111_10001110_1;
      patterns[38906] = 25'b10010111_11111000_10001111_1;
      patterns[38907] = 25'b10010111_11111001_10010000_1;
      patterns[38908] = 25'b10010111_11111010_10010001_1;
      patterns[38909] = 25'b10010111_11111011_10010010_1;
      patterns[38910] = 25'b10010111_11111100_10010011_1;
      patterns[38911] = 25'b10010111_11111101_10010100_1;
      patterns[38912] = 25'b10010111_11111110_10010101_1;
      patterns[38913] = 25'b10010111_11111111_10010110_1;
      patterns[38914] = 25'b10011000_00000000_10011000_0;
      patterns[38915] = 25'b10011000_00000001_10011001_0;
      patterns[38916] = 25'b10011000_00000010_10011010_0;
      patterns[38917] = 25'b10011000_00000011_10011011_0;
      patterns[38918] = 25'b10011000_00000100_10011100_0;
      patterns[38919] = 25'b10011000_00000101_10011101_0;
      patterns[38920] = 25'b10011000_00000110_10011110_0;
      patterns[38921] = 25'b10011000_00000111_10011111_0;
      patterns[38922] = 25'b10011000_00001000_10100000_0;
      patterns[38923] = 25'b10011000_00001001_10100001_0;
      patterns[38924] = 25'b10011000_00001010_10100010_0;
      patterns[38925] = 25'b10011000_00001011_10100011_0;
      patterns[38926] = 25'b10011000_00001100_10100100_0;
      patterns[38927] = 25'b10011000_00001101_10100101_0;
      patterns[38928] = 25'b10011000_00001110_10100110_0;
      patterns[38929] = 25'b10011000_00001111_10100111_0;
      patterns[38930] = 25'b10011000_00010000_10101000_0;
      patterns[38931] = 25'b10011000_00010001_10101001_0;
      patterns[38932] = 25'b10011000_00010010_10101010_0;
      patterns[38933] = 25'b10011000_00010011_10101011_0;
      patterns[38934] = 25'b10011000_00010100_10101100_0;
      patterns[38935] = 25'b10011000_00010101_10101101_0;
      patterns[38936] = 25'b10011000_00010110_10101110_0;
      patterns[38937] = 25'b10011000_00010111_10101111_0;
      patterns[38938] = 25'b10011000_00011000_10110000_0;
      patterns[38939] = 25'b10011000_00011001_10110001_0;
      patterns[38940] = 25'b10011000_00011010_10110010_0;
      patterns[38941] = 25'b10011000_00011011_10110011_0;
      patterns[38942] = 25'b10011000_00011100_10110100_0;
      patterns[38943] = 25'b10011000_00011101_10110101_0;
      patterns[38944] = 25'b10011000_00011110_10110110_0;
      patterns[38945] = 25'b10011000_00011111_10110111_0;
      patterns[38946] = 25'b10011000_00100000_10111000_0;
      patterns[38947] = 25'b10011000_00100001_10111001_0;
      patterns[38948] = 25'b10011000_00100010_10111010_0;
      patterns[38949] = 25'b10011000_00100011_10111011_0;
      patterns[38950] = 25'b10011000_00100100_10111100_0;
      patterns[38951] = 25'b10011000_00100101_10111101_0;
      patterns[38952] = 25'b10011000_00100110_10111110_0;
      patterns[38953] = 25'b10011000_00100111_10111111_0;
      patterns[38954] = 25'b10011000_00101000_11000000_0;
      patterns[38955] = 25'b10011000_00101001_11000001_0;
      patterns[38956] = 25'b10011000_00101010_11000010_0;
      patterns[38957] = 25'b10011000_00101011_11000011_0;
      patterns[38958] = 25'b10011000_00101100_11000100_0;
      patterns[38959] = 25'b10011000_00101101_11000101_0;
      patterns[38960] = 25'b10011000_00101110_11000110_0;
      patterns[38961] = 25'b10011000_00101111_11000111_0;
      patterns[38962] = 25'b10011000_00110000_11001000_0;
      patterns[38963] = 25'b10011000_00110001_11001001_0;
      patterns[38964] = 25'b10011000_00110010_11001010_0;
      patterns[38965] = 25'b10011000_00110011_11001011_0;
      patterns[38966] = 25'b10011000_00110100_11001100_0;
      patterns[38967] = 25'b10011000_00110101_11001101_0;
      patterns[38968] = 25'b10011000_00110110_11001110_0;
      patterns[38969] = 25'b10011000_00110111_11001111_0;
      patterns[38970] = 25'b10011000_00111000_11010000_0;
      patterns[38971] = 25'b10011000_00111001_11010001_0;
      patterns[38972] = 25'b10011000_00111010_11010010_0;
      patterns[38973] = 25'b10011000_00111011_11010011_0;
      patterns[38974] = 25'b10011000_00111100_11010100_0;
      patterns[38975] = 25'b10011000_00111101_11010101_0;
      patterns[38976] = 25'b10011000_00111110_11010110_0;
      patterns[38977] = 25'b10011000_00111111_11010111_0;
      patterns[38978] = 25'b10011000_01000000_11011000_0;
      patterns[38979] = 25'b10011000_01000001_11011001_0;
      patterns[38980] = 25'b10011000_01000010_11011010_0;
      patterns[38981] = 25'b10011000_01000011_11011011_0;
      patterns[38982] = 25'b10011000_01000100_11011100_0;
      patterns[38983] = 25'b10011000_01000101_11011101_0;
      patterns[38984] = 25'b10011000_01000110_11011110_0;
      patterns[38985] = 25'b10011000_01000111_11011111_0;
      patterns[38986] = 25'b10011000_01001000_11100000_0;
      patterns[38987] = 25'b10011000_01001001_11100001_0;
      patterns[38988] = 25'b10011000_01001010_11100010_0;
      patterns[38989] = 25'b10011000_01001011_11100011_0;
      patterns[38990] = 25'b10011000_01001100_11100100_0;
      patterns[38991] = 25'b10011000_01001101_11100101_0;
      patterns[38992] = 25'b10011000_01001110_11100110_0;
      patterns[38993] = 25'b10011000_01001111_11100111_0;
      patterns[38994] = 25'b10011000_01010000_11101000_0;
      patterns[38995] = 25'b10011000_01010001_11101001_0;
      patterns[38996] = 25'b10011000_01010010_11101010_0;
      patterns[38997] = 25'b10011000_01010011_11101011_0;
      patterns[38998] = 25'b10011000_01010100_11101100_0;
      patterns[38999] = 25'b10011000_01010101_11101101_0;
      patterns[39000] = 25'b10011000_01010110_11101110_0;
      patterns[39001] = 25'b10011000_01010111_11101111_0;
      patterns[39002] = 25'b10011000_01011000_11110000_0;
      patterns[39003] = 25'b10011000_01011001_11110001_0;
      patterns[39004] = 25'b10011000_01011010_11110010_0;
      patterns[39005] = 25'b10011000_01011011_11110011_0;
      patterns[39006] = 25'b10011000_01011100_11110100_0;
      patterns[39007] = 25'b10011000_01011101_11110101_0;
      patterns[39008] = 25'b10011000_01011110_11110110_0;
      patterns[39009] = 25'b10011000_01011111_11110111_0;
      patterns[39010] = 25'b10011000_01100000_11111000_0;
      patterns[39011] = 25'b10011000_01100001_11111001_0;
      patterns[39012] = 25'b10011000_01100010_11111010_0;
      patterns[39013] = 25'b10011000_01100011_11111011_0;
      patterns[39014] = 25'b10011000_01100100_11111100_0;
      patterns[39015] = 25'b10011000_01100101_11111101_0;
      patterns[39016] = 25'b10011000_01100110_11111110_0;
      patterns[39017] = 25'b10011000_01100111_11111111_0;
      patterns[39018] = 25'b10011000_01101000_00000000_1;
      patterns[39019] = 25'b10011000_01101001_00000001_1;
      patterns[39020] = 25'b10011000_01101010_00000010_1;
      patterns[39021] = 25'b10011000_01101011_00000011_1;
      patterns[39022] = 25'b10011000_01101100_00000100_1;
      patterns[39023] = 25'b10011000_01101101_00000101_1;
      patterns[39024] = 25'b10011000_01101110_00000110_1;
      patterns[39025] = 25'b10011000_01101111_00000111_1;
      patterns[39026] = 25'b10011000_01110000_00001000_1;
      patterns[39027] = 25'b10011000_01110001_00001001_1;
      patterns[39028] = 25'b10011000_01110010_00001010_1;
      patterns[39029] = 25'b10011000_01110011_00001011_1;
      patterns[39030] = 25'b10011000_01110100_00001100_1;
      patterns[39031] = 25'b10011000_01110101_00001101_1;
      patterns[39032] = 25'b10011000_01110110_00001110_1;
      patterns[39033] = 25'b10011000_01110111_00001111_1;
      patterns[39034] = 25'b10011000_01111000_00010000_1;
      patterns[39035] = 25'b10011000_01111001_00010001_1;
      patterns[39036] = 25'b10011000_01111010_00010010_1;
      patterns[39037] = 25'b10011000_01111011_00010011_1;
      patterns[39038] = 25'b10011000_01111100_00010100_1;
      patterns[39039] = 25'b10011000_01111101_00010101_1;
      patterns[39040] = 25'b10011000_01111110_00010110_1;
      patterns[39041] = 25'b10011000_01111111_00010111_1;
      patterns[39042] = 25'b10011000_10000000_00011000_1;
      patterns[39043] = 25'b10011000_10000001_00011001_1;
      patterns[39044] = 25'b10011000_10000010_00011010_1;
      patterns[39045] = 25'b10011000_10000011_00011011_1;
      patterns[39046] = 25'b10011000_10000100_00011100_1;
      patterns[39047] = 25'b10011000_10000101_00011101_1;
      patterns[39048] = 25'b10011000_10000110_00011110_1;
      patterns[39049] = 25'b10011000_10000111_00011111_1;
      patterns[39050] = 25'b10011000_10001000_00100000_1;
      patterns[39051] = 25'b10011000_10001001_00100001_1;
      patterns[39052] = 25'b10011000_10001010_00100010_1;
      patterns[39053] = 25'b10011000_10001011_00100011_1;
      patterns[39054] = 25'b10011000_10001100_00100100_1;
      patterns[39055] = 25'b10011000_10001101_00100101_1;
      patterns[39056] = 25'b10011000_10001110_00100110_1;
      patterns[39057] = 25'b10011000_10001111_00100111_1;
      patterns[39058] = 25'b10011000_10010000_00101000_1;
      patterns[39059] = 25'b10011000_10010001_00101001_1;
      patterns[39060] = 25'b10011000_10010010_00101010_1;
      patterns[39061] = 25'b10011000_10010011_00101011_1;
      patterns[39062] = 25'b10011000_10010100_00101100_1;
      patterns[39063] = 25'b10011000_10010101_00101101_1;
      patterns[39064] = 25'b10011000_10010110_00101110_1;
      patterns[39065] = 25'b10011000_10010111_00101111_1;
      patterns[39066] = 25'b10011000_10011000_00110000_1;
      patterns[39067] = 25'b10011000_10011001_00110001_1;
      patterns[39068] = 25'b10011000_10011010_00110010_1;
      patterns[39069] = 25'b10011000_10011011_00110011_1;
      patterns[39070] = 25'b10011000_10011100_00110100_1;
      patterns[39071] = 25'b10011000_10011101_00110101_1;
      patterns[39072] = 25'b10011000_10011110_00110110_1;
      patterns[39073] = 25'b10011000_10011111_00110111_1;
      patterns[39074] = 25'b10011000_10100000_00111000_1;
      patterns[39075] = 25'b10011000_10100001_00111001_1;
      patterns[39076] = 25'b10011000_10100010_00111010_1;
      patterns[39077] = 25'b10011000_10100011_00111011_1;
      patterns[39078] = 25'b10011000_10100100_00111100_1;
      patterns[39079] = 25'b10011000_10100101_00111101_1;
      patterns[39080] = 25'b10011000_10100110_00111110_1;
      patterns[39081] = 25'b10011000_10100111_00111111_1;
      patterns[39082] = 25'b10011000_10101000_01000000_1;
      patterns[39083] = 25'b10011000_10101001_01000001_1;
      patterns[39084] = 25'b10011000_10101010_01000010_1;
      patterns[39085] = 25'b10011000_10101011_01000011_1;
      patterns[39086] = 25'b10011000_10101100_01000100_1;
      patterns[39087] = 25'b10011000_10101101_01000101_1;
      patterns[39088] = 25'b10011000_10101110_01000110_1;
      patterns[39089] = 25'b10011000_10101111_01000111_1;
      patterns[39090] = 25'b10011000_10110000_01001000_1;
      patterns[39091] = 25'b10011000_10110001_01001001_1;
      patterns[39092] = 25'b10011000_10110010_01001010_1;
      patterns[39093] = 25'b10011000_10110011_01001011_1;
      patterns[39094] = 25'b10011000_10110100_01001100_1;
      patterns[39095] = 25'b10011000_10110101_01001101_1;
      patterns[39096] = 25'b10011000_10110110_01001110_1;
      patterns[39097] = 25'b10011000_10110111_01001111_1;
      patterns[39098] = 25'b10011000_10111000_01010000_1;
      patterns[39099] = 25'b10011000_10111001_01010001_1;
      patterns[39100] = 25'b10011000_10111010_01010010_1;
      patterns[39101] = 25'b10011000_10111011_01010011_1;
      patterns[39102] = 25'b10011000_10111100_01010100_1;
      patterns[39103] = 25'b10011000_10111101_01010101_1;
      patterns[39104] = 25'b10011000_10111110_01010110_1;
      patterns[39105] = 25'b10011000_10111111_01010111_1;
      patterns[39106] = 25'b10011000_11000000_01011000_1;
      patterns[39107] = 25'b10011000_11000001_01011001_1;
      patterns[39108] = 25'b10011000_11000010_01011010_1;
      patterns[39109] = 25'b10011000_11000011_01011011_1;
      patterns[39110] = 25'b10011000_11000100_01011100_1;
      patterns[39111] = 25'b10011000_11000101_01011101_1;
      patterns[39112] = 25'b10011000_11000110_01011110_1;
      patterns[39113] = 25'b10011000_11000111_01011111_1;
      patterns[39114] = 25'b10011000_11001000_01100000_1;
      patterns[39115] = 25'b10011000_11001001_01100001_1;
      patterns[39116] = 25'b10011000_11001010_01100010_1;
      patterns[39117] = 25'b10011000_11001011_01100011_1;
      patterns[39118] = 25'b10011000_11001100_01100100_1;
      patterns[39119] = 25'b10011000_11001101_01100101_1;
      patterns[39120] = 25'b10011000_11001110_01100110_1;
      patterns[39121] = 25'b10011000_11001111_01100111_1;
      patterns[39122] = 25'b10011000_11010000_01101000_1;
      patterns[39123] = 25'b10011000_11010001_01101001_1;
      patterns[39124] = 25'b10011000_11010010_01101010_1;
      patterns[39125] = 25'b10011000_11010011_01101011_1;
      patterns[39126] = 25'b10011000_11010100_01101100_1;
      patterns[39127] = 25'b10011000_11010101_01101101_1;
      patterns[39128] = 25'b10011000_11010110_01101110_1;
      patterns[39129] = 25'b10011000_11010111_01101111_1;
      patterns[39130] = 25'b10011000_11011000_01110000_1;
      patterns[39131] = 25'b10011000_11011001_01110001_1;
      patterns[39132] = 25'b10011000_11011010_01110010_1;
      patterns[39133] = 25'b10011000_11011011_01110011_1;
      patterns[39134] = 25'b10011000_11011100_01110100_1;
      patterns[39135] = 25'b10011000_11011101_01110101_1;
      patterns[39136] = 25'b10011000_11011110_01110110_1;
      patterns[39137] = 25'b10011000_11011111_01110111_1;
      patterns[39138] = 25'b10011000_11100000_01111000_1;
      patterns[39139] = 25'b10011000_11100001_01111001_1;
      patterns[39140] = 25'b10011000_11100010_01111010_1;
      patterns[39141] = 25'b10011000_11100011_01111011_1;
      patterns[39142] = 25'b10011000_11100100_01111100_1;
      patterns[39143] = 25'b10011000_11100101_01111101_1;
      patterns[39144] = 25'b10011000_11100110_01111110_1;
      patterns[39145] = 25'b10011000_11100111_01111111_1;
      patterns[39146] = 25'b10011000_11101000_10000000_1;
      patterns[39147] = 25'b10011000_11101001_10000001_1;
      patterns[39148] = 25'b10011000_11101010_10000010_1;
      patterns[39149] = 25'b10011000_11101011_10000011_1;
      patterns[39150] = 25'b10011000_11101100_10000100_1;
      patterns[39151] = 25'b10011000_11101101_10000101_1;
      patterns[39152] = 25'b10011000_11101110_10000110_1;
      patterns[39153] = 25'b10011000_11101111_10000111_1;
      patterns[39154] = 25'b10011000_11110000_10001000_1;
      patterns[39155] = 25'b10011000_11110001_10001001_1;
      patterns[39156] = 25'b10011000_11110010_10001010_1;
      patterns[39157] = 25'b10011000_11110011_10001011_1;
      patterns[39158] = 25'b10011000_11110100_10001100_1;
      patterns[39159] = 25'b10011000_11110101_10001101_1;
      patterns[39160] = 25'b10011000_11110110_10001110_1;
      patterns[39161] = 25'b10011000_11110111_10001111_1;
      patterns[39162] = 25'b10011000_11111000_10010000_1;
      patterns[39163] = 25'b10011000_11111001_10010001_1;
      patterns[39164] = 25'b10011000_11111010_10010010_1;
      patterns[39165] = 25'b10011000_11111011_10010011_1;
      patterns[39166] = 25'b10011000_11111100_10010100_1;
      patterns[39167] = 25'b10011000_11111101_10010101_1;
      patterns[39168] = 25'b10011000_11111110_10010110_1;
      patterns[39169] = 25'b10011000_11111111_10010111_1;
      patterns[39170] = 25'b10011001_00000000_10011001_0;
      patterns[39171] = 25'b10011001_00000001_10011010_0;
      patterns[39172] = 25'b10011001_00000010_10011011_0;
      patterns[39173] = 25'b10011001_00000011_10011100_0;
      patterns[39174] = 25'b10011001_00000100_10011101_0;
      patterns[39175] = 25'b10011001_00000101_10011110_0;
      patterns[39176] = 25'b10011001_00000110_10011111_0;
      patterns[39177] = 25'b10011001_00000111_10100000_0;
      patterns[39178] = 25'b10011001_00001000_10100001_0;
      patterns[39179] = 25'b10011001_00001001_10100010_0;
      patterns[39180] = 25'b10011001_00001010_10100011_0;
      patterns[39181] = 25'b10011001_00001011_10100100_0;
      patterns[39182] = 25'b10011001_00001100_10100101_0;
      patterns[39183] = 25'b10011001_00001101_10100110_0;
      patterns[39184] = 25'b10011001_00001110_10100111_0;
      patterns[39185] = 25'b10011001_00001111_10101000_0;
      patterns[39186] = 25'b10011001_00010000_10101001_0;
      patterns[39187] = 25'b10011001_00010001_10101010_0;
      patterns[39188] = 25'b10011001_00010010_10101011_0;
      patterns[39189] = 25'b10011001_00010011_10101100_0;
      patterns[39190] = 25'b10011001_00010100_10101101_0;
      patterns[39191] = 25'b10011001_00010101_10101110_0;
      patterns[39192] = 25'b10011001_00010110_10101111_0;
      patterns[39193] = 25'b10011001_00010111_10110000_0;
      patterns[39194] = 25'b10011001_00011000_10110001_0;
      patterns[39195] = 25'b10011001_00011001_10110010_0;
      patterns[39196] = 25'b10011001_00011010_10110011_0;
      patterns[39197] = 25'b10011001_00011011_10110100_0;
      patterns[39198] = 25'b10011001_00011100_10110101_0;
      patterns[39199] = 25'b10011001_00011101_10110110_0;
      patterns[39200] = 25'b10011001_00011110_10110111_0;
      patterns[39201] = 25'b10011001_00011111_10111000_0;
      patterns[39202] = 25'b10011001_00100000_10111001_0;
      patterns[39203] = 25'b10011001_00100001_10111010_0;
      patterns[39204] = 25'b10011001_00100010_10111011_0;
      patterns[39205] = 25'b10011001_00100011_10111100_0;
      patterns[39206] = 25'b10011001_00100100_10111101_0;
      patterns[39207] = 25'b10011001_00100101_10111110_0;
      patterns[39208] = 25'b10011001_00100110_10111111_0;
      patterns[39209] = 25'b10011001_00100111_11000000_0;
      patterns[39210] = 25'b10011001_00101000_11000001_0;
      patterns[39211] = 25'b10011001_00101001_11000010_0;
      patterns[39212] = 25'b10011001_00101010_11000011_0;
      patterns[39213] = 25'b10011001_00101011_11000100_0;
      patterns[39214] = 25'b10011001_00101100_11000101_0;
      patterns[39215] = 25'b10011001_00101101_11000110_0;
      patterns[39216] = 25'b10011001_00101110_11000111_0;
      patterns[39217] = 25'b10011001_00101111_11001000_0;
      patterns[39218] = 25'b10011001_00110000_11001001_0;
      patterns[39219] = 25'b10011001_00110001_11001010_0;
      patterns[39220] = 25'b10011001_00110010_11001011_0;
      patterns[39221] = 25'b10011001_00110011_11001100_0;
      patterns[39222] = 25'b10011001_00110100_11001101_0;
      patterns[39223] = 25'b10011001_00110101_11001110_0;
      patterns[39224] = 25'b10011001_00110110_11001111_0;
      patterns[39225] = 25'b10011001_00110111_11010000_0;
      patterns[39226] = 25'b10011001_00111000_11010001_0;
      patterns[39227] = 25'b10011001_00111001_11010010_0;
      patterns[39228] = 25'b10011001_00111010_11010011_0;
      patterns[39229] = 25'b10011001_00111011_11010100_0;
      patterns[39230] = 25'b10011001_00111100_11010101_0;
      patterns[39231] = 25'b10011001_00111101_11010110_0;
      patterns[39232] = 25'b10011001_00111110_11010111_0;
      patterns[39233] = 25'b10011001_00111111_11011000_0;
      patterns[39234] = 25'b10011001_01000000_11011001_0;
      patterns[39235] = 25'b10011001_01000001_11011010_0;
      patterns[39236] = 25'b10011001_01000010_11011011_0;
      patterns[39237] = 25'b10011001_01000011_11011100_0;
      patterns[39238] = 25'b10011001_01000100_11011101_0;
      patterns[39239] = 25'b10011001_01000101_11011110_0;
      patterns[39240] = 25'b10011001_01000110_11011111_0;
      patterns[39241] = 25'b10011001_01000111_11100000_0;
      patterns[39242] = 25'b10011001_01001000_11100001_0;
      patterns[39243] = 25'b10011001_01001001_11100010_0;
      patterns[39244] = 25'b10011001_01001010_11100011_0;
      patterns[39245] = 25'b10011001_01001011_11100100_0;
      patterns[39246] = 25'b10011001_01001100_11100101_0;
      patterns[39247] = 25'b10011001_01001101_11100110_0;
      patterns[39248] = 25'b10011001_01001110_11100111_0;
      patterns[39249] = 25'b10011001_01001111_11101000_0;
      patterns[39250] = 25'b10011001_01010000_11101001_0;
      patterns[39251] = 25'b10011001_01010001_11101010_0;
      patterns[39252] = 25'b10011001_01010010_11101011_0;
      patterns[39253] = 25'b10011001_01010011_11101100_0;
      patterns[39254] = 25'b10011001_01010100_11101101_0;
      patterns[39255] = 25'b10011001_01010101_11101110_0;
      patterns[39256] = 25'b10011001_01010110_11101111_0;
      patterns[39257] = 25'b10011001_01010111_11110000_0;
      patterns[39258] = 25'b10011001_01011000_11110001_0;
      patterns[39259] = 25'b10011001_01011001_11110010_0;
      patterns[39260] = 25'b10011001_01011010_11110011_0;
      patterns[39261] = 25'b10011001_01011011_11110100_0;
      patterns[39262] = 25'b10011001_01011100_11110101_0;
      patterns[39263] = 25'b10011001_01011101_11110110_0;
      patterns[39264] = 25'b10011001_01011110_11110111_0;
      patterns[39265] = 25'b10011001_01011111_11111000_0;
      patterns[39266] = 25'b10011001_01100000_11111001_0;
      patterns[39267] = 25'b10011001_01100001_11111010_0;
      patterns[39268] = 25'b10011001_01100010_11111011_0;
      patterns[39269] = 25'b10011001_01100011_11111100_0;
      patterns[39270] = 25'b10011001_01100100_11111101_0;
      patterns[39271] = 25'b10011001_01100101_11111110_0;
      patterns[39272] = 25'b10011001_01100110_11111111_0;
      patterns[39273] = 25'b10011001_01100111_00000000_1;
      patterns[39274] = 25'b10011001_01101000_00000001_1;
      patterns[39275] = 25'b10011001_01101001_00000010_1;
      patterns[39276] = 25'b10011001_01101010_00000011_1;
      patterns[39277] = 25'b10011001_01101011_00000100_1;
      patterns[39278] = 25'b10011001_01101100_00000101_1;
      patterns[39279] = 25'b10011001_01101101_00000110_1;
      patterns[39280] = 25'b10011001_01101110_00000111_1;
      patterns[39281] = 25'b10011001_01101111_00001000_1;
      patterns[39282] = 25'b10011001_01110000_00001001_1;
      patterns[39283] = 25'b10011001_01110001_00001010_1;
      patterns[39284] = 25'b10011001_01110010_00001011_1;
      patterns[39285] = 25'b10011001_01110011_00001100_1;
      patterns[39286] = 25'b10011001_01110100_00001101_1;
      patterns[39287] = 25'b10011001_01110101_00001110_1;
      patterns[39288] = 25'b10011001_01110110_00001111_1;
      patterns[39289] = 25'b10011001_01110111_00010000_1;
      patterns[39290] = 25'b10011001_01111000_00010001_1;
      patterns[39291] = 25'b10011001_01111001_00010010_1;
      patterns[39292] = 25'b10011001_01111010_00010011_1;
      patterns[39293] = 25'b10011001_01111011_00010100_1;
      patterns[39294] = 25'b10011001_01111100_00010101_1;
      patterns[39295] = 25'b10011001_01111101_00010110_1;
      patterns[39296] = 25'b10011001_01111110_00010111_1;
      patterns[39297] = 25'b10011001_01111111_00011000_1;
      patterns[39298] = 25'b10011001_10000000_00011001_1;
      patterns[39299] = 25'b10011001_10000001_00011010_1;
      patterns[39300] = 25'b10011001_10000010_00011011_1;
      patterns[39301] = 25'b10011001_10000011_00011100_1;
      patterns[39302] = 25'b10011001_10000100_00011101_1;
      patterns[39303] = 25'b10011001_10000101_00011110_1;
      patterns[39304] = 25'b10011001_10000110_00011111_1;
      patterns[39305] = 25'b10011001_10000111_00100000_1;
      patterns[39306] = 25'b10011001_10001000_00100001_1;
      patterns[39307] = 25'b10011001_10001001_00100010_1;
      patterns[39308] = 25'b10011001_10001010_00100011_1;
      patterns[39309] = 25'b10011001_10001011_00100100_1;
      patterns[39310] = 25'b10011001_10001100_00100101_1;
      patterns[39311] = 25'b10011001_10001101_00100110_1;
      patterns[39312] = 25'b10011001_10001110_00100111_1;
      patterns[39313] = 25'b10011001_10001111_00101000_1;
      patterns[39314] = 25'b10011001_10010000_00101001_1;
      patterns[39315] = 25'b10011001_10010001_00101010_1;
      patterns[39316] = 25'b10011001_10010010_00101011_1;
      patterns[39317] = 25'b10011001_10010011_00101100_1;
      patterns[39318] = 25'b10011001_10010100_00101101_1;
      patterns[39319] = 25'b10011001_10010101_00101110_1;
      patterns[39320] = 25'b10011001_10010110_00101111_1;
      patterns[39321] = 25'b10011001_10010111_00110000_1;
      patterns[39322] = 25'b10011001_10011000_00110001_1;
      patterns[39323] = 25'b10011001_10011001_00110010_1;
      patterns[39324] = 25'b10011001_10011010_00110011_1;
      patterns[39325] = 25'b10011001_10011011_00110100_1;
      patterns[39326] = 25'b10011001_10011100_00110101_1;
      patterns[39327] = 25'b10011001_10011101_00110110_1;
      patterns[39328] = 25'b10011001_10011110_00110111_1;
      patterns[39329] = 25'b10011001_10011111_00111000_1;
      patterns[39330] = 25'b10011001_10100000_00111001_1;
      patterns[39331] = 25'b10011001_10100001_00111010_1;
      patterns[39332] = 25'b10011001_10100010_00111011_1;
      patterns[39333] = 25'b10011001_10100011_00111100_1;
      patterns[39334] = 25'b10011001_10100100_00111101_1;
      patterns[39335] = 25'b10011001_10100101_00111110_1;
      patterns[39336] = 25'b10011001_10100110_00111111_1;
      patterns[39337] = 25'b10011001_10100111_01000000_1;
      patterns[39338] = 25'b10011001_10101000_01000001_1;
      patterns[39339] = 25'b10011001_10101001_01000010_1;
      patterns[39340] = 25'b10011001_10101010_01000011_1;
      patterns[39341] = 25'b10011001_10101011_01000100_1;
      patterns[39342] = 25'b10011001_10101100_01000101_1;
      patterns[39343] = 25'b10011001_10101101_01000110_1;
      patterns[39344] = 25'b10011001_10101110_01000111_1;
      patterns[39345] = 25'b10011001_10101111_01001000_1;
      patterns[39346] = 25'b10011001_10110000_01001001_1;
      patterns[39347] = 25'b10011001_10110001_01001010_1;
      patterns[39348] = 25'b10011001_10110010_01001011_1;
      patterns[39349] = 25'b10011001_10110011_01001100_1;
      patterns[39350] = 25'b10011001_10110100_01001101_1;
      patterns[39351] = 25'b10011001_10110101_01001110_1;
      patterns[39352] = 25'b10011001_10110110_01001111_1;
      patterns[39353] = 25'b10011001_10110111_01010000_1;
      patterns[39354] = 25'b10011001_10111000_01010001_1;
      patterns[39355] = 25'b10011001_10111001_01010010_1;
      patterns[39356] = 25'b10011001_10111010_01010011_1;
      patterns[39357] = 25'b10011001_10111011_01010100_1;
      patterns[39358] = 25'b10011001_10111100_01010101_1;
      patterns[39359] = 25'b10011001_10111101_01010110_1;
      patterns[39360] = 25'b10011001_10111110_01010111_1;
      patterns[39361] = 25'b10011001_10111111_01011000_1;
      patterns[39362] = 25'b10011001_11000000_01011001_1;
      patterns[39363] = 25'b10011001_11000001_01011010_1;
      patterns[39364] = 25'b10011001_11000010_01011011_1;
      patterns[39365] = 25'b10011001_11000011_01011100_1;
      patterns[39366] = 25'b10011001_11000100_01011101_1;
      patterns[39367] = 25'b10011001_11000101_01011110_1;
      patterns[39368] = 25'b10011001_11000110_01011111_1;
      patterns[39369] = 25'b10011001_11000111_01100000_1;
      patterns[39370] = 25'b10011001_11001000_01100001_1;
      patterns[39371] = 25'b10011001_11001001_01100010_1;
      patterns[39372] = 25'b10011001_11001010_01100011_1;
      patterns[39373] = 25'b10011001_11001011_01100100_1;
      patterns[39374] = 25'b10011001_11001100_01100101_1;
      patterns[39375] = 25'b10011001_11001101_01100110_1;
      patterns[39376] = 25'b10011001_11001110_01100111_1;
      patterns[39377] = 25'b10011001_11001111_01101000_1;
      patterns[39378] = 25'b10011001_11010000_01101001_1;
      patterns[39379] = 25'b10011001_11010001_01101010_1;
      patterns[39380] = 25'b10011001_11010010_01101011_1;
      patterns[39381] = 25'b10011001_11010011_01101100_1;
      patterns[39382] = 25'b10011001_11010100_01101101_1;
      patterns[39383] = 25'b10011001_11010101_01101110_1;
      patterns[39384] = 25'b10011001_11010110_01101111_1;
      patterns[39385] = 25'b10011001_11010111_01110000_1;
      patterns[39386] = 25'b10011001_11011000_01110001_1;
      patterns[39387] = 25'b10011001_11011001_01110010_1;
      patterns[39388] = 25'b10011001_11011010_01110011_1;
      patterns[39389] = 25'b10011001_11011011_01110100_1;
      patterns[39390] = 25'b10011001_11011100_01110101_1;
      patterns[39391] = 25'b10011001_11011101_01110110_1;
      patterns[39392] = 25'b10011001_11011110_01110111_1;
      patterns[39393] = 25'b10011001_11011111_01111000_1;
      patterns[39394] = 25'b10011001_11100000_01111001_1;
      patterns[39395] = 25'b10011001_11100001_01111010_1;
      patterns[39396] = 25'b10011001_11100010_01111011_1;
      patterns[39397] = 25'b10011001_11100011_01111100_1;
      patterns[39398] = 25'b10011001_11100100_01111101_1;
      patterns[39399] = 25'b10011001_11100101_01111110_1;
      patterns[39400] = 25'b10011001_11100110_01111111_1;
      patterns[39401] = 25'b10011001_11100111_10000000_1;
      patterns[39402] = 25'b10011001_11101000_10000001_1;
      patterns[39403] = 25'b10011001_11101001_10000010_1;
      patterns[39404] = 25'b10011001_11101010_10000011_1;
      patterns[39405] = 25'b10011001_11101011_10000100_1;
      patterns[39406] = 25'b10011001_11101100_10000101_1;
      patterns[39407] = 25'b10011001_11101101_10000110_1;
      patterns[39408] = 25'b10011001_11101110_10000111_1;
      patterns[39409] = 25'b10011001_11101111_10001000_1;
      patterns[39410] = 25'b10011001_11110000_10001001_1;
      patterns[39411] = 25'b10011001_11110001_10001010_1;
      patterns[39412] = 25'b10011001_11110010_10001011_1;
      patterns[39413] = 25'b10011001_11110011_10001100_1;
      patterns[39414] = 25'b10011001_11110100_10001101_1;
      patterns[39415] = 25'b10011001_11110101_10001110_1;
      patterns[39416] = 25'b10011001_11110110_10001111_1;
      patterns[39417] = 25'b10011001_11110111_10010000_1;
      patterns[39418] = 25'b10011001_11111000_10010001_1;
      patterns[39419] = 25'b10011001_11111001_10010010_1;
      patterns[39420] = 25'b10011001_11111010_10010011_1;
      patterns[39421] = 25'b10011001_11111011_10010100_1;
      patterns[39422] = 25'b10011001_11111100_10010101_1;
      patterns[39423] = 25'b10011001_11111101_10010110_1;
      patterns[39424] = 25'b10011001_11111110_10010111_1;
      patterns[39425] = 25'b10011001_11111111_10011000_1;
      patterns[39426] = 25'b10011010_00000000_10011010_0;
      patterns[39427] = 25'b10011010_00000001_10011011_0;
      patterns[39428] = 25'b10011010_00000010_10011100_0;
      patterns[39429] = 25'b10011010_00000011_10011101_0;
      patterns[39430] = 25'b10011010_00000100_10011110_0;
      patterns[39431] = 25'b10011010_00000101_10011111_0;
      patterns[39432] = 25'b10011010_00000110_10100000_0;
      patterns[39433] = 25'b10011010_00000111_10100001_0;
      patterns[39434] = 25'b10011010_00001000_10100010_0;
      patterns[39435] = 25'b10011010_00001001_10100011_0;
      patterns[39436] = 25'b10011010_00001010_10100100_0;
      patterns[39437] = 25'b10011010_00001011_10100101_0;
      patterns[39438] = 25'b10011010_00001100_10100110_0;
      patterns[39439] = 25'b10011010_00001101_10100111_0;
      patterns[39440] = 25'b10011010_00001110_10101000_0;
      patterns[39441] = 25'b10011010_00001111_10101001_0;
      patterns[39442] = 25'b10011010_00010000_10101010_0;
      patterns[39443] = 25'b10011010_00010001_10101011_0;
      patterns[39444] = 25'b10011010_00010010_10101100_0;
      patterns[39445] = 25'b10011010_00010011_10101101_0;
      patterns[39446] = 25'b10011010_00010100_10101110_0;
      patterns[39447] = 25'b10011010_00010101_10101111_0;
      patterns[39448] = 25'b10011010_00010110_10110000_0;
      patterns[39449] = 25'b10011010_00010111_10110001_0;
      patterns[39450] = 25'b10011010_00011000_10110010_0;
      patterns[39451] = 25'b10011010_00011001_10110011_0;
      patterns[39452] = 25'b10011010_00011010_10110100_0;
      patterns[39453] = 25'b10011010_00011011_10110101_0;
      patterns[39454] = 25'b10011010_00011100_10110110_0;
      patterns[39455] = 25'b10011010_00011101_10110111_0;
      patterns[39456] = 25'b10011010_00011110_10111000_0;
      patterns[39457] = 25'b10011010_00011111_10111001_0;
      patterns[39458] = 25'b10011010_00100000_10111010_0;
      patterns[39459] = 25'b10011010_00100001_10111011_0;
      patterns[39460] = 25'b10011010_00100010_10111100_0;
      patterns[39461] = 25'b10011010_00100011_10111101_0;
      patterns[39462] = 25'b10011010_00100100_10111110_0;
      patterns[39463] = 25'b10011010_00100101_10111111_0;
      patterns[39464] = 25'b10011010_00100110_11000000_0;
      patterns[39465] = 25'b10011010_00100111_11000001_0;
      patterns[39466] = 25'b10011010_00101000_11000010_0;
      patterns[39467] = 25'b10011010_00101001_11000011_0;
      patterns[39468] = 25'b10011010_00101010_11000100_0;
      patterns[39469] = 25'b10011010_00101011_11000101_0;
      patterns[39470] = 25'b10011010_00101100_11000110_0;
      patterns[39471] = 25'b10011010_00101101_11000111_0;
      patterns[39472] = 25'b10011010_00101110_11001000_0;
      patterns[39473] = 25'b10011010_00101111_11001001_0;
      patterns[39474] = 25'b10011010_00110000_11001010_0;
      patterns[39475] = 25'b10011010_00110001_11001011_0;
      patterns[39476] = 25'b10011010_00110010_11001100_0;
      patterns[39477] = 25'b10011010_00110011_11001101_0;
      patterns[39478] = 25'b10011010_00110100_11001110_0;
      patterns[39479] = 25'b10011010_00110101_11001111_0;
      patterns[39480] = 25'b10011010_00110110_11010000_0;
      patterns[39481] = 25'b10011010_00110111_11010001_0;
      patterns[39482] = 25'b10011010_00111000_11010010_0;
      patterns[39483] = 25'b10011010_00111001_11010011_0;
      patterns[39484] = 25'b10011010_00111010_11010100_0;
      patterns[39485] = 25'b10011010_00111011_11010101_0;
      patterns[39486] = 25'b10011010_00111100_11010110_0;
      patterns[39487] = 25'b10011010_00111101_11010111_0;
      patterns[39488] = 25'b10011010_00111110_11011000_0;
      patterns[39489] = 25'b10011010_00111111_11011001_0;
      patterns[39490] = 25'b10011010_01000000_11011010_0;
      patterns[39491] = 25'b10011010_01000001_11011011_0;
      patterns[39492] = 25'b10011010_01000010_11011100_0;
      patterns[39493] = 25'b10011010_01000011_11011101_0;
      patterns[39494] = 25'b10011010_01000100_11011110_0;
      patterns[39495] = 25'b10011010_01000101_11011111_0;
      patterns[39496] = 25'b10011010_01000110_11100000_0;
      patterns[39497] = 25'b10011010_01000111_11100001_0;
      patterns[39498] = 25'b10011010_01001000_11100010_0;
      patterns[39499] = 25'b10011010_01001001_11100011_0;
      patterns[39500] = 25'b10011010_01001010_11100100_0;
      patterns[39501] = 25'b10011010_01001011_11100101_0;
      patterns[39502] = 25'b10011010_01001100_11100110_0;
      patterns[39503] = 25'b10011010_01001101_11100111_0;
      patterns[39504] = 25'b10011010_01001110_11101000_0;
      patterns[39505] = 25'b10011010_01001111_11101001_0;
      patterns[39506] = 25'b10011010_01010000_11101010_0;
      patterns[39507] = 25'b10011010_01010001_11101011_0;
      patterns[39508] = 25'b10011010_01010010_11101100_0;
      patterns[39509] = 25'b10011010_01010011_11101101_0;
      patterns[39510] = 25'b10011010_01010100_11101110_0;
      patterns[39511] = 25'b10011010_01010101_11101111_0;
      patterns[39512] = 25'b10011010_01010110_11110000_0;
      patterns[39513] = 25'b10011010_01010111_11110001_0;
      patterns[39514] = 25'b10011010_01011000_11110010_0;
      patterns[39515] = 25'b10011010_01011001_11110011_0;
      patterns[39516] = 25'b10011010_01011010_11110100_0;
      patterns[39517] = 25'b10011010_01011011_11110101_0;
      patterns[39518] = 25'b10011010_01011100_11110110_0;
      patterns[39519] = 25'b10011010_01011101_11110111_0;
      patterns[39520] = 25'b10011010_01011110_11111000_0;
      patterns[39521] = 25'b10011010_01011111_11111001_0;
      patterns[39522] = 25'b10011010_01100000_11111010_0;
      patterns[39523] = 25'b10011010_01100001_11111011_0;
      patterns[39524] = 25'b10011010_01100010_11111100_0;
      patterns[39525] = 25'b10011010_01100011_11111101_0;
      patterns[39526] = 25'b10011010_01100100_11111110_0;
      patterns[39527] = 25'b10011010_01100101_11111111_0;
      patterns[39528] = 25'b10011010_01100110_00000000_1;
      patterns[39529] = 25'b10011010_01100111_00000001_1;
      patterns[39530] = 25'b10011010_01101000_00000010_1;
      patterns[39531] = 25'b10011010_01101001_00000011_1;
      patterns[39532] = 25'b10011010_01101010_00000100_1;
      patterns[39533] = 25'b10011010_01101011_00000101_1;
      patterns[39534] = 25'b10011010_01101100_00000110_1;
      patterns[39535] = 25'b10011010_01101101_00000111_1;
      patterns[39536] = 25'b10011010_01101110_00001000_1;
      patterns[39537] = 25'b10011010_01101111_00001001_1;
      patterns[39538] = 25'b10011010_01110000_00001010_1;
      patterns[39539] = 25'b10011010_01110001_00001011_1;
      patterns[39540] = 25'b10011010_01110010_00001100_1;
      patterns[39541] = 25'b10011010_01110011_00001101_1;
      patterns[39542] = 25'b10011010_01110100_00001110_1;
      patterns[39543] = 25'b10011010_01110101_00001111_1;
      patterns[39544] = 25'b10011010_01110110_00010000_1;
      patterns[39545] = 25'b10011010_01110111_00010001_1;
      patterns[39546] = 25'b10011010_01111000_00010010_1;
      patterns[39547] = 25'b10011010_01111001_00010011_1;
      patterns[39548] = 25'b10011010_01111010_00010100_1;
      patterns[39549] = 25'b10011010_01111011_00010101_1;
      patterns[39550] = 25'b10011010_01111100_00010110_1;
      patterns[39551] = 25'b10011010_01111101_00010111_1;
      patterns[39552] = 25'b10011010_01111110_00011000_1;
      patterns[39553] = 25'b10011010_01111111_00011001_1;
      patterns[39554] = 25'b10011010_10000000_00011010_1;
      patterns[39555] = 25'b10011010_10000001_00011011_1;
      patterns[39556] = 25'b10011010_10000010_00011100_1;
      patterns[39557] = 25'b10011010_10000011_00011101_1;
      patterns[39558] = 25'b10011010_10000100_00011110_1;
      patterns[39559] = 25'b10011010_10000101_00011111_1;
      patterns[39560] = 25'b10011010_10000110_00100000_1;
      patterns[39561] = 25'b10011010_10000111_00100001_1;
      patterns[39562] = 25'b10011010_10001000_00100010_1;
      patterns[39563] = 25'b10011010_10001001_00100011_1;
      patterns[39564] = 25'b10011010_10001010_00100100_1;
      patterns[39565] = 25'b10011010_10001011_00100101_1;
      patterns[39566] = 25'b10011010_10001100_00100110_1;
      patterns[39567] = 25'b10011010_10001101_00100111_1;
      patterns[39568] = 25'b10011010_10001110_00101000_1;
      patterns[39569] = 25'b10011010_10001111_00101001_1;
      patterns[39570] = 25'b10011010_10010000_00101010_1;
      patterns[39571] = 25'b10011010_10010001_00101011_1;
      patterns[39572] = 25'b10011010_10010010_00101100_1;
      patterns[39573] = 25'b10011010_10010011_00101101_1;
      patterns[39574] = 25'b10011010_10010100_00101110_1;
      patterns[39575] = 25'b10011010_10010101_00101111_1;
      patterns[39576] = 25'b10011010_10010110_00110000_1;
      patterns[39577] = 25'b10011010_10010111_00110001_1;
      patterns[39578] = 25'b10011010_10011000_00110010_1;
      patterns[39579] = 25'b10011010_10011001_00110011_1;
      patterns[39580] = 25'b10011010_10011010_00110100_1;
      patterns[39581] = 25'b10011010_10011011_00110101_1;
      patterns[39582] = 25'b10011010_10011100_00110110_1;
      patterns[39583] = 25'b10011010_10011101_00110111_1;
      patterns[39584] = 25'b10011010_10011110_00111000_1;
      patterns[39585] = 25'b10011010_10011111_00111001_1;
      patterns[39586] = 25'b10011010_10100000_00111010_1;
      patterns[39587] = 25'b10011010_10100001_00111011_1;
      patterns[39588] = 25'b10011010_10100010_00111100_1;
      patterns[39589] = 25'b10011010_10100011_00111101_1;
      patterns[39590] = 25'b10011010_10100100_00111110_1;
      patterns[39591] = 25'b10011010_10100101_00111111_1;
      patterns[39592] = 25'b10011010_10100110_01000000_1;
      patterns[39593] = 25'b10011010_10100111_01000001_1;
      patterns[39594] = 25'b10011010_10101000_01000010_1;
      patterns[39595] = 25'b10011010_10101001_01000011_1;
      patterns[39596] = 25'b10011010_10101010_01000100_1;
      patterns[39597] = 25'b10011010_10101011_01000101_1;
      patterns[39598] = 25'b10011010_10101100_01000110_1;
      patterns[39599] = 25'b10011010_10101101_01000111_1;
      patterns[39600] = 25'b10011010_10101110_01001000_1;
      patterns[39601] = 25'b10011010_10101111_01001001_1;
      patterns[39602] = 25'b10011010_10110000_01001010_1;
      patterns[39603] = 25'b10011010_10110001_01001011_1;
      patterns[39604] = 25'b10011010_10110010_01001100_1;
      patterns[39605] = 25'b10011010_10110011_01001101_1;
      patterns[39606] = 25'b10011010_10110100_01001110_1;
      patterns[39607] = 25'b10011010_10110101_01001111_1;
      patterns[39608] = 25'b10011010_10110110_01010000_1;
      patterns[39609] = 25'b10011010_10110111_01010001_1;
      patterns[39610] = 25'b10011010_10111000_01010010_1;
      patterns[39611] = 25'b10011010_10111001_01010011_1;
      patterns[39612] = 25'b10011010_10111010_01010100_1;
      patterns[39613] = 25'b10011010_10111011_01010101_1;
      patterns[39614] = 25'b10011010_10111100_01010110_1;
      patterns[39615] = 25'b10011010_10111101_01010111_1;
      patterns[39616] = 25'b10011010_10111110_01011000_1;
      patterns[39617] = 25'b10011010_10111111_01011001_1;
      patterns[39618] = 25'b10011010_11000000_01011010_1;
      patterns[39619] = 25'b10011010_11000001_01011011_1;
      patterns[39620] = 25'b10011010_11000010_01011100_1;
      patterns[39621] = 25'b10011010_11000011_01011101_1;
      patterns[39622] = 25'b10011010_11000100_01011110_1;
      patterns[39623] = 25'b10011010_11000101_01011111_1;
      patterns[39624] = 25'b10011010_11000110_01100000_1;
      patterns[39625] = 25'b10011010_11000111_01100001_1;
      patterns[39626] = 25'b10011010_11001000_01100010_1;
      patterns[39627] = 25'b10011010_11001001_01100011_1;
      patterns[39628] = 25'b10011010_11001010_01100100_1;
      patterns[39629] = 25'b10011010_11001011_01100101_1;
      patterns[39630] = 25'b10011010_11001100_01100110_1;
      patterns[39631] = 25'b10011010_11001101_01100111_1;
      patterns[39632] = 25'b10011010_11001110_01101000_1;
      patterns[39633] = 25'b10011010_11001111_01101001_1;
      patterns[39634] = 25'b10011010_11010000_01101010_1;
      patterns[39635] = 25'b10011010_11010001_01101011_1;
      patterns[39636] = 25'b10011010_11010010_01101100_1;
      patterns[39637] = 25'b10011010_11010011_01101101_1;
      patterns[39638] = 25'b10011010_11010100_01101110_1;
      patterns[39639] = 25'b10011010_11010101_01101111_1;
      patterns[39640] = 25'b10011010_11010110_01110000_1;
      patterns[39641] = 25'b10011010_11010111_01110001_1;
      patterns[39642] = 25'b10011010_11011000_01110010_1;
      patterns[39643] = 25'b10011010_11011001_01110011_1;
      patterns[39644] = 25'b10011010_11011010_01110100_1;
      patterns[39645] = 25'b10011010_11011011_01110101_1;
      patterns[39646] = 25'b10011010_11011100_01110110_1;
      patterns[39647] = 25'b10011010_11011101_01110111_1;
      patterns[39648] = 25'b10011010_11011110_01111000_1;
      patterns[39649] = 25'b10011010_11011111_01111001_1;
      patterns[39650] = 25'b10011010_11100000_01111010_1;
      patterns[39651] = 25'b10011010_11100001_01111011_1;
      patterns[39652] = 25'b10011010_11100010_01111100_1;
      patterns[39653] = 25'b10011010_11100011_01111101_1;
      patterns[39654] = 25'b10011010_11100100_01111110_1;
      patterns[39655] = 25'b10011010_11100101_01111111_1;
      patterns[39656] = 25'b10011010_11100110_10000000_1;
      patterns[39657] = 25'b10011010_11100111_10000001_1;
      patterns[39658] = 25'b10011010_11101000_10000010_1;
      patterns[39659] = 25'b10011010_11101001_10000011_1;
      patterns[39660] = 25'b10011010_11101010_10000100_1;
      patterns[39661] = 25'b10011010_11101011_10000101_1;
      patterns[39662] = 25'b10011010_11101100_10000110_1;
      patterns[39663] = 25'b10011010_11101101_10000111_1;
      patterns[39664] = 25'b10011010_11101110_10001000_1;
      patterns[39665] = 25'b10011010_11101111_10001001_1;
      patterns[39666] = 25'b10011010_11110000_10001010_1;
      patterns[39667] = 25'b10011010_11110001_10001011_1;
      patterns[39668] = 25'b10011010_11110010_10001100_1;
      patterns[39669] = 25'b10011010_11110011_10001101_1;
      patterns[39670] = 25'b10011010_11110100_10001110_1;
      patterns[39671] = 25'b10011010_11110101_10001111_1;
      patterns[39672] = 25'b10011010_11110110_10010000_1;
      patterns[39673] = 25'b10011010_11110111_10010001_1;
      patterns[39674] = 25'b10011010_11111000_10010010_1;
      patterns[39675] = 25'b10011010_11111001_10010011_1;
      patterns[39676] = 25'b10011010_11111010_10010100_1;
      patterns[39677] = 25'b10011010_11111011_10010101_1;
      patterns[39678] = 25'b10011010_11111100_10010110_1;
      patterns[39679] = 25'b10011010_11111101_10010111_1;
      patterns[39680] = 25'b10011010_11111110_10011000_1;
      patterns[39681] = 25'b10011010_11111111_10011001_1;
      patterns[39682] = 25'b10011011_00000000_10011011_0;
      patterns[39683] = 25'b10011011_00000001_10011100_0;
      patterns[39684] = 25'b10011011_00000010_10011101_0;
      patterns[39685] = 25'b10011011_00000011_10011110_0;
      patterns[39686] = 25'b10011011_00000100_10011111_0;
      patterns[39687] = 25'b10011011_00000101_10100000_0;
      patterns[39688] = 25'b10011011_00000110_10100001_0;
      patterns[39689] = 25'b10011011_00000111_10100010_0;
      patterns[39690] = 25'b10011011_00001000_10100011_0;
      patterns[39691] = 25'b10011011_00001001_10100100_0;
      patterns[39692] = 25'b10011011_00001010_10100101_0;
      patterns[39693] = 25'b10011011_00001011_10100110_0;
      patterns[39694] = 25'b10011011_00001100_10100111_0;
      patterns[39695] = 25'b10011011_00001101_10101000_0;
      patterns[39696] = 25'b10011011_00001110_10101001_0;
      patterns[39697] = 25'b10011011_00001111_10101010_0;
      patterns[39698] = 25'b10011011_00010000_10101011_0;
      patterns[39699] = 25'b10011011_00010001_10101100_0;
      patterns[39700] = 25'b10011011_00010010_10101101_0;
      patterns[39701] = 25'b10011011_00010011_10101110_0;
      patterns[39702] = 25'b10011011_00010100_10101111_0;
      patterns[39703] = 25'b10011011_00010101_10110000_0;
      patterns[39704] = 25'b10011011_00010110_10110001_0;
      patterns[39705] = 25'b10011011_00010111_10110010_0;
      patterns[39706] = 25'b10011011_00011000_10110011_0;
      patterns[39707] = 25'b10011011_00011001_10110100_0;
      patterns[39708] = 25'b10011011_00011010_10110101_0;
      patterns[39709] = 25'b10011011_00011011_10110110_0;
      patterns[39710] = 25'b10011011_00011100_10110111_0;
      patterns[39711] = 25'b10011011_00011101_10111000_0;
      patterns[39712] = 25'b10011011_00011110_10111001_0;
      patterns[39713] = 25'b10011011_00011111_10111010_0;
      patterns[39714] = 25'b10011011_00100000_10111011_0;
      patterns[39715] = 25'b10011011_00100001_10111100_0;
      patterns[39716] = 25'b10011011_00100010_10111101_0;
      patterns[39717] = 25'b10011011_00100011_10111110_0;
      patterns[39718] = 25'b10011011_00100100_10111111_0;
      patterns[39719] = 25'b10011011_00100101_11000000_0;
      patterns[39720] = 25'b10011011_00100110_11000001_0;
      patterns[39721] = 25'b10011011_00100111_11000010_0;
      patterns[39722] = 25'b10011011_00101000_11000011_0;
      patterns[39723] = 25'b10011011_00101001_11000100_0;
      patterns[39724] = 25'b10011011_00101010_11000101_0;
      patterns[39725] = 25'b10011011_00101011_11000110_0;
      patterns[39726] = 25'b10011011_00101100_11000111_0;
      patterns[39727] = 25'b10011011_00101101_11001000_0;
      patterns[39728] = 25'b10011011_00101110_11001001_0;
      patterns[39729] = 25'b10011011_00101111_11001010_0;
      patterns[39730] = 25'b10011011_00110000_11001011_0;
      patterns[39731] = 25'b10011011_00110001_11001100_0;
      patterns[39732] = 25'b10011011_00110010_11001101_0;
      patterns[39733] = 25'b10011011_00110011_11001110_0;
      patterns[39734] = 25'b10011011_00110100_11001111_0;
      patterns[39735] = 25'b10011011_00110101_11010000_0;
      patterns[39736] = 25'b10011011_00110110_11010001_0;
      patterns[39737] = 25'b10011011_00110111_11010010_0;
      patterns[39738] = 25'b10011011_00111000_11010011_0;
      patterns[39739] = 25'b10011011_00111001_11010100_0;
      patterns[39740] = 25'b10011011_00111010_11010101_0;
      patterns[39741] = 25'b10011011_00111011_11010110_0;
      patterns[39742] = 25'b10011011_00111100_11010111_0;
      patterns[39743] = 25'b10011011_00111101_11011000_0;
      patterns[39744] = 25'b10011011_00111110_11011001_0;
      patterns[39745] = 25'b10011011_00111111_11011010_0;
      patterns[39746] = 25'b10011011_01000000_11011011_0;
      patterns[39747] = 25'b10011011_01000001_11011100_0;
      patterns[39748] = 25'b10011011_01000010_11011101_0;
      patterns[39749] = 25'b10011011_01000011_11011110_0;
      patterns[39750] = 25'b10011011_01000100_11011111_0;
      patterns[39751] = 25'b10011011_01000101_11100000_0;
      patterns[39752] = 25'b10011011_01000110_11100001_0;
      patterns[39753] = 25'b10011011_01000111_11100010_0;
      patterns[39754] = 25'b10011011_01001000_11100011_0;
      patterns[39755] = 25'b10011011_01001001_11100100_0;
      patterns[39756] = 25'b10011011_01001010_11100101_0;
      patterns[39757] = 25'b10011011_01001011_11100110_0;
      patterns[39758] = 25'b10011011_01001100_11100111_0;
      patterns[39759] = 25'b10011011_01001101_11101000_0;
      patterns[39760] = 25'b10011011_01001110_11101001_0;
      patterns[39761] = 25'b10011011_01001111_11101010_0;
      patterns[39762] = 25'b10011011_01010000_11101011_0;
      patterns[39763] = 25'b10011011_01010001_11101100_0;
      patterns[39764] = 25'b10011011_01010010_11101101_0;
      patterns[39765] = 25'b10011011_01010011_11101110_0;
      patterns[39766] = 25'b10011011_01010100_11101111_0;
      patterns[39767] = 25'b10011011_01010101_11110000_0;
      patterns[39768] = 25'b10011011_01010110_11110001_0;
      patterns[39769] = 25'b10011011_01010111_11110010_0;
      patterns[39770] = 25'b10011011_01011000_11110011_0;
      patterns[39771] = 25'b10011011_01011001_11110100_0;
      patterns[39772] = 25'b10011011_01011010_11110101_0;
      patterns[39773] = 25'b10011011_01011011_11110110_0;
      patterns[39774] = 25'b10011011_01011100_11110111_0;
      patterns[39775] = 25'b10011011_01011101_11111000_0;
      patterns[39776] = 25'b10011011_01011110_11111001_0;
      patterns[39777] = 25'b10011011_01011111_11111010_0;
      patterns[39778] = 25'b10011011_01100000_11111011_0;
      patterns[39779] = 25'b10011011_01100001_11111100_0;
      patterns[39780] = 25'b10011011_01100010_11111101_0;
      patterns[39781] = 25'b10011011_01100011_11111110_0;
      patterns[39782] = 25'b10011011_01100100_11111111_0;
      patterns[39783] = 25'b10011011_01100101_00000000_1;
      patterns[39784] = 25'b10011011_01100110_00000001_1;
      patterns[39785] = 25'b10011011_01100111_00000010_1;
      patterns[39786] = 25'b10011011_01101000_00000011_1;
      patterns[39787] = 25'b10011011_01101001_00000100_1;
      patterns[39788] = 25'b10011011_01101010_00000101_1;
      patterns[39789] = 25'b10011011_01101011_00000110_1;
      patterns[39790] = 25'b10011011_01101100_00000111_1;
      patterns[39791] = 25'b10011011_01101101_00001000_1;
      patterns[39792] = 25'b10011011_01101110_00001001_1;
      patterns[39793] = 25'b10011011_01101111_00001010_1;
      patterns[39794] = 25'b10011011_01110000_00001011_1;
      patterns[39795] = 25'b10011011_01110001_00001100_1;
      patterns[39796] = 25'b10011011_01110010_00001101_1;
      patterns[39797] = 25'b10011011_01110011_00001110_1;
      patterns[39798] = 25'b10011011_01110100_00001111_1;
      patterns[39799] = 25'b10011011_01110101_00010000_1;
      patterns[39800] = 25'b10011011_01110110_00010001_1;
      patterns[39801] = 25'b10011011_01110111_00010010_1;
      patterns[39802] = 25'b10011011_01111000_00010011_1;
      patterns[39803] = 25'b10011011_01111001_00010100_1;
      patterns[39804] = 25'b10011011_01111010_00010101_1;
      patterns[39805] = 25'b10011011_01111011_00010110_1;
      patterns[39806] = 25'b10011011_01111100_00010111_1;
      patterns[39807] = 25'b10011011_01111101_00011000_1;
      patterns[39808] = 25'b10011011_01111110_00011001_1;
      patterns[39809] = 25'b10011011_01111111_00011010_1;
      patterns[39810] = 25'b10011011_10000000_00011011_1;
      patterns[39811] = 25'b10011011_10000001_00011100_1;
      patterns[39812] = 25'b10011011_10000010_00011101_1;
      patterns[39813] = 25'b10011011_10000011_00011110_1;
      patterns[39814] = 25'b10011011_10000100_00011111_1;
      patterns[39815] = 25'b10011011_10000101_00100000_1;
      patterns[39816] = 25'b10011011_10000110_00100001_1;
      patterns[39817] = 25'b10011011_10000111_00100010_1;
      patterns[39818] = 25'b10011011_10001000_00100011_1;
      patterns[39819] = 25'b10011011_10001001_00100100_1;
      patterns[39820] = 25'b10011011_10001010_00100101_1;
      patterns[39821] = 25'b10011011_10001011_00100110_1;
      patterns[39822] = 25'b10011011_10001100_00100111_1;
      patterns[39823] = 25'b10011011_10001101_00101000_1;
      patterns[39824] = 25'b10011011_10001110_00101001_1;
      patterns[39825] = 25'b10011011_10001111_00101010_1;
      patterns[39826] = 25'b10011011_10010000_00101011_1;
      patterns[39827] = 25'b10011011_10010001_00101100_1;
      patterns[39828] = 25'b10011011_10010010_00101101_1;
      patterns[39829] = 25'b10011011_10010011_00101110_1;
      patterns[39830] = 25'b10011011_10010100_00101111_1;
      patterns[39831] = 25'b10011011_10010101_00110000_1;
      patterns[39832] = 25'b10011011_10010110_00110001_1;
      patterns[39833] = 25'b10011011_10010111_00110010_1;
      patterns[39834] = 25'b10011011_10011000_00110011_1;
      patterns[39835] = 25'b10011011_10011001_00110100_1;
      patterns[39836] = 25'b10011011_10011010_00110101_1;
      patterns[39837] = 25'b10011011_10011011_00110110_1;
      patterns[39838] = 25'b10011011_10011100_00110111_1;
      patterns[39839] = 25'b10011011_10011101_00111000_1;
      patterns[39840] = 25'b10011011_10011110_00111001_1;
      patterns[39841] = 25'b10011011_10011111_00111010_1;
      patterns[39842] = 25'b10011011_10100000_00111011_1;
      patterns[39843] = 25'b10011011_10100001_00111100_1;
      patterns[39844] = 25'b10011011_10100010_00111101_1;
      patterns[39845] = 25'b10011011_10100011_00111110_1;
      patterns[39846] = 25'b10011011_10100100_00111111_1;
      patterns[39847] = 25'b10011011_10100101_01000000_1;
      patterns[39848] = 25'b10011011_10100110_01000001_1;
      patterns[39849] = 25'b10011011_10100111_01000010_1;
      patterns[39850] = 25'b10011011_10101000_01000011_1;
      patterns[39851] = 25'b10011011_10101001_01000100_1;
      patterns[39852] = 25'b10011011_10101010_01000101_1;
      patterns[39853] = 25'b10011011_10101011_01000110_1;
      patterns[39854] = 25'b10011011_10101100_01000111_1;
      patterns[39855] = 25'b10011011_10101101_01001000_1;
      patterns[39856] = 25'b10011011_10101110_01001001_1;
      patterns[39857] = 25'b10011011_10101111_01001010_1;
      patterns[39858] = 25'b10011011_10110000_01001011_1;
      patterns[39859] = 25'b10011011_10110001_01001100_1;
      patterns[39860] = 25'b10011011_10110010_01001101_1;
      patterns[39861] = 25'b10011011_10110011_01001110_1;
      patterns[39862] = 25'b10011011_10110100_01001111_1;
      patterns[39863] = 25'b10011011_10110101_01010000_1;
      patterns[39864] = 25'b10011011_10110110_01010001_1;
      patterns[39865] = 25'b10011011_10110111_01010010_1;
      patterns[39866] = 25'b10011011_10111000_01010011_1;
      patterns[39867] = 25'b10011011_10111001_01010100_1;
      patterns[39868] = 25'b10011011_10111010_01010101_1;
      patterns[39869] = 25'b10011011_10111011_01010110_1;
      patterns[39870] = 25'b10011011_10111100_01010111_1;
      patterns[39871] = 25'b10011011_10111101_01011000_1;
      patterns[39872] = 25'b10011011_10111110_01011001_1;
      patterns[39873] = 25'b10011011_10111111_01011010_1;
      patterns[39874] = 25'b10011011_11000000_01011011_1;
      patterns[39875] = 25'b10011011_11000001_01011100_1;
      patterns[39876] = 25'b10011011_11000010_01011101_1;
      patterns[39877] = 25'b10011011_11000011_01011110_1;
      patterns[39878] = 25'b10011011_11000100_01011111_1;
      patterns[39879] = 25'b10011011_11000101_01100000_1;
      patterns[39880] = 25'b10011011_11000110_01100001_1;
      patterns[39881] = 25'b10011011_11000111_01100010_1;
      patterns[39882] = 25'b10011011_11001000_01100011_1;
      patterns[39883] = 25'b10011011_11001001_01100100_1;
      patterns[39884] = 25'b10011011_11001010_01100101_1;
      patterns[39885] = 25'b10011011_11001011_01100110_1;
      patterns[39886] = 25'b10011011_11001100_01100111_1;
      patterns[39887] = 25'b10011011_11001101_01101000_1;
      patterns[39888] = 25'b10011011_11001110_01101001_1;
      patterns[39889] = 25'b10011011_11001111_01101010_1;
      patterns[39890] = 25'b10011011_11010000_01101011_1;
      patterns[39891] = 25'b10011011_11010001_01101100_1;
      patterns[39892] = 25'b10011011_11010010_01101101_1;
      patterns[39893] = 25'b10011011_11010011_01101110_1;
      patterns[39894] = 25'b10011011_11010100_01101111_1;
      patterns[39895] = 25'b10011011_11010101_01110000_1;
      patterns[39896] = 25'b10011011_11010110_01110001_1;
      patterns[39897] = 25'b10011011_11010111_01110010_1;
      patterns[39898] = 25'b10011011_11011000_01110011_1;
      patterns[39899] = 25'b10011011_11011001_01110100_1;
      patterns[39900] = 25'b10011011_11011010_01110101_1;
      patterns[39901] = 25'b10011011_11011011_01110110_1;
      patterns[39902] = 25'b10011011_11011100_01110111_1;
      patterns[39903] = 25'b10011011_11011101_01111000_1;
      patterns[39904] = 25'b10011011_11011110_01111001_1;
      patterns[39905] = 25'b10011011_11011111_01111010_1;
      patterns[39906] = 25'b10011011_11100000_01111011_1;
      patterns[39907] = 25'b10011011_11100001_01111100_1;
      patterns[39908] = 25'b10011011_11100010_01111101_1;
      patterns[39909] = 25'b10011011_11100011_01111110_1;
      patterns[39910] = 25'b10011011_11100100_01111111_1;
      patterns[39911] = 25'b10011011_11100101_10000000_1;
      patterns[39912] = 25'b10011011_11100110_10000001_1;
      patterns[39913] = 25'b10011011_11100111_10000010_1;
      patterns[39914] = 25'b10011011_11101000_10000011_1;
      patterns[39915] = 25'b10011011_11101001_10000100_1;
      patterns[39916] = 25'b10011011_11101010_10000101_1;
      patterns[39917] = 25'b10011011_11101011_10000110_1;
      patterns[39918] = 25'b10011011_11101100_10000111_1;
      patterns[39919] = 25'b10011011_11101101_10001000_1;
      patterns[39920] = 25'b10011011_11101110_10001001_1;
      patterns[39921] = 25'b10011011_11101111_10001010_1;
      patterns[39922] = 25'b10011011_11110000_10001011_1;
      patterns[39923] = 25'b10011011_11110001_10001100_1;
      patterns[39924] = 25'b10011011_11110010_10001101_1;
      patterns[39925] = 25'b10011011_11110011_10001110_1;
      patterns[39926] = 25'b10011011_11110100_10001111_1;
      patterns[39927] = 25'b10011011_11110101_10010000_1;
      patterns[39928] = 25'b10011011_11110110_10010001_1;
      patterns[39929] = 25'b10011011_11110111_10010010_1;
      patterns[39930] = 25'b10011011_11111000_10010011_1;
      patterns[39931] = 25'b10011011_11111001_10010100_1;
      patterns[39932] = 25'b10011011_11111010_10010101_1;
      patterns[39933] = 25'b10011011_11111011_10010110_1;
      patterns[39934] = 25'b10011011_11111100_10010111_1;
      patterns[39935] = 25'b10011011_11111101_10011000_1;
      patterns[39936] = 25'b10011011_11111110_10011001_1;
      patterns[39937] = 25'b10011011_11111111_10011010_1;
      patterns[39938] = 25'b10011100_00000000_10011100_0;
      patterns[39939] = 25'b10011100_00000001_10011101_0;
      patterns[39940] = 25'b10011100_00000010_10011110_0;
      patterns[39941] = 25'b10011100_00000011_10011111_0;
      patterns[39942] = 25'b10011100_00000100_10100000_0;
      patterns[39943] = 25'b10011100_00000101_10100001_0;
      patterns[39944] = 25'b10011100_00000110_10100010_0;
      patterns[39945] = 25'b10011100_00000111_10100011_0;
      patterns[39946] = 25'b10011100_00001000_10100100_0;
      patterns[39947] = 25'b10011100_00001001_10100101_0;
      patterns[39948] = 25'b10011100_00001010_10100110_0;
      patterns[39949] = 25'b10011100_00001011_10100111_0;
      patterns[39950] = 25'b10011100_00001100_10101000_0;
      patterns[39951] = 25'b10011100_00001101_10101001_0;
      patterns[39952] = 25'b10011100_00001110_10101010_0;
      patterns[39953] = 25'b10011100_00001111_10101011_0;
      patterns[39954] = 25'b10011100_00010000_10101100_0;
      patterns[39955] = 25'b10011100_00010001_10101101_0;
      patterns[39956] = 25'b10011100_00010010_10101110_0;
      patterns[39957] = 25'b10011100_00010011_10101111_0;
      patterns[39958] = 25'b10011100_00010100_10110000_0;
      patterns[39959] = 25'b10011100_00010101_10110001_0;
      patterns[39960] = 25'b10011100_00010110_10110010_0;
      patterns[39961] = 25'b10011100_00010111_10110011_0;
      patterns[39962] = 25'b10011100_00011000_10110100_0;
      patterns[39963] = 25'b10011100_00011001_10110101_0;
      patterns[39964] = 25'b10011100_00011010_10110110_0;
      patterns[39965] = 25'b10011100_00011011_10110111_0;
      patterns[39966] = 25'b10011100_00011100_10111000_0;
      patterns[39967] = 25'b10011100_00011101_10111001_0;
      patterns[39968] = 25'b10011100_00011110_10111010_0;
      patterns[39969] = 25'b10011100_00011111_10111011_0;
      patterns[39970] = 25'b10011100_00100000_10111100_0;
      patterns[39971] = 25'b10011100_00100001_10111101_0;
      patterns[39972] = 25'b10011100_00100010_10111110_0;
      patterns[39973] = 25'b10011100_00100011_10111111_0;
      patterns[39974] = 25'b10011100_00100100_11000000_0;
      patterns[39975] = 25'b10011100_00100101_11000001_0;
      patterns[39976] = 25'b10011100_00100110_11000010_0;
      patterns[39977] = 25'b10011100_00100111_11000011_0;
      patterns[39978] = 25'b10011100_00101000_11000100_0;
      patterns[39979] = 25'b10011100_00101001_11000101_0;
      patterns[39980] = 25'b10011100_00101010_11000110_0;
      patterns[39981] = 25'b10011100_00101011_11000111_0;
      patterns[39982] = 25'b10011100_00101100_11001000_0;
      patterns[39983] = 25'b10011100_00101101_11001001_0;
      patterns[39984] = 25'b10011100_00101110_11001010_0;
      patterns[39985] = 25'b10011100_00101111_11001011_0;
      patterns[39986] = 25'b10011100_00110000_11001100_0;
      patterns[39987] = 25'b10011100_00110001_11001101_0;
      patterns[39988] = 25'b10011100_00110010_11001110_0;
      patterns[39989] = 25'b10011100_00110011_11001111_0;
      patterns[39990] = 25'b10011100_00110100_11010000_0;
      patterns[39991] = 25'b10011100_00110101_11010001_0;
      patterns[39992] = 25'b10011100_00110110_11010010_0;
      patterns[39993] = 25'b10011100_00110111_11010011_0;
      patterns[39994] = 25'b10011100_00111000_11010100_0;
      patterns[39995] = 25'b10011100_00111001_11010101_0;
      patterns[39996] = 25'b10011100_00111010_11010110_0;
      patterns[39997] = 25'b10011100_00111011_11010111_0;
      patterns[39998] = 25'b10011100_00111100_11011000_0;
      patterns[39999] = 25'b10011100_00111101_11011001_0;
      patterns[40000] = 25'b10011100_00111110_11011010_0;
      patterns[40001] = 25'b10011100_00111111_11011011_0;
      patterns[40002] = 25'b10011100_01000000_11011100_0;
      patterns[40003] = 25'b10011100_01000001_11011101_0;
      patterns[40004] = 25'b10011100_01000010_11011110_0;
      patterns[40005] = 25'b10011100_01000011_11011111_0;
      patterns[40006] = 25'b10011100_01000100_11100000_0;
      patterns[40007] = 25'b10011100_01000101_11100001_0;
      patterns[40008] = 25'b10011100_01000110_11100010_0;
      patterns[40009] = 25'b10011100_01000111_11100011_0;
      patterns[40010] = 25'b10011100_01001000_11100100_0;
      patterns[40011] = 25'b10011100_01001001_11100101_0;
      patterns[40012] = 25'b10011100_01001010_11100110_0;
      patterns[40013] = 25'b10011100_01001011_11100111_0;
      patterns[40014] = 25'b10011100_01001100_11101000_0;
      patterns[40015] = 25'b10011100_01001101_11101001_0;
      patterns[40016] = 25'b10011100_01001110_11101010_0;
      patterns[40017] = 25'b10011100_01001111_11101011_0;
      patterns[40018] = 25'b10011100_01010000_11101100_0;
      patterns[40019] = 25'b10011100_01010001_11101101_0;
      patterns[40020] = 25'b10011100_01010010_11101110_0;
      patterns[40021] = 25'b10011100_01010011_11101111_0;
      patterns[40022] = 25'b10011100_01010100_11110000_0;
      patterns[40023] = 25'b10011100_01010101_11110001_0;
      patterns[40024] = 25'b10011100_01010110_11110010_0;
      patterns[40025] = 25'b10011100_01010111_11110011_0;
      patterns[40026] = 25'b10011100_01011000_11110100_0;
      patterns[40027] = 25'b10011100_01011001_11110101_0;
      patterns[40028] = 25'b10011100_01011010_11110110_0;
      patterns[40029] = 25'b10011100_01011011_11110111_0;
      patterns[40030] = 25'b10011100_01011100_11111000_0;
      patterns[40031] = 25'b10011100_01011101_11111001_0;
      patterns[40032] = 25'b10011100_01011110_11111010_0;
      patterns[40033] = 25'b10011100_01011111_11111011_0;
      patterns[40034] = 25'b10011100_01100000_11111100_0;
      patterns[40035] = 25'b10011100_01100001_11111101_0;
      patterns[40036] = 25'b10011100_01100010_11111110_0;
      patterns[40037] = 25'b10011100_01100011_11111111_0;
      patterns[40038] = 25'b10011100_01100100_00000000_1;
      patterns[40039] = 25'b10011100_01100101_00000001_1;
      patterns[40040] = 25'b10011100_01100110_00000010_1;
      patterns[40041] = 25'b10011100_01100111_00000011_1;
      patterns[40042] = 25'b10011100_01101000_00000100_1;
      patterns[40043] = 25'b10011100_01101001_00000101_1;
      patterns[40044] = 25'b10011100_01101010_00000110_1;
      patterns[40045] = 25'b10011100_01101011_00000111_1;
      patterns[40046] = 25'b10011100_01101100_00001000_1;
      patterns[40047] = 25'b10011100_01101101_00001001_1;
      patterns[40048] = 25'b10011100_01101110_00001010_1;
      patterns[40049] = 25'b10011100_01101111_00001011_1;
      patterns[40050] = 25'b10011100_01110000_00001100_1;
      patterns[40051] = 25'b10011100_01110001_00001101_1;
      patterns[40052] = 25'b10011100_01110010_00001110_1;
      patterns[40053] = 25'b10011100_01110011_00001111_1;
      patterns[40054] = 25'b10011100_01110100_00010000_1;
      patterns[40055] = 25'b10011100_01110101_00010001_1;
      patterns[40056] = 25'b10011100_01110110_00010010_1;
      patterns[40057] = 25'b10011100_01110111_00010011_1;
      patterns[40058] = 25'b10011100_01111000_00010100_1;
      patterns[40059] = 25'b10011100_01111001_00010101_1;
      patterns[40060] = 25'b10011100_01111010_00010110_1;
      patterns[40061] = 25'b10011100_01111011_00010111_1;
      patterns[40062] = 25'b10011100_01111100_00011000_1;
      patterns[40063] = 25'b10011100_01111101_00011001_1;
      patterns[40064] = 25'b10011100_01111110_00011010_1;
      patterns[40065] = 25'b10011100_01111111_00011011_1;
      patterns[40066] = 25'b10011100_10000000_00011100_1;
      patterns[40067] = 25'b10011100_10000001_00011101_1;
      patterns[40068] = 25'b10011100_10000010_00011110_1;
      patterns[40069] = 25'b10011100_10000011_00011111_1;
      patterns[40070] = 25'b10011100_10000100_00100000_1;
      patterns[40071] = 25'b10011100_10000101_00100001_1;
      patterns[40072] = 25'b10011100_10000110_00100010_1;
      patterns[40073] = 25'b10011100_10000111_00100011_1;
      patterns[40074] = 25'b10011100_10001000_00100100_1;
      patterns[40075] = 25'b10011100_10001001_00100101_1;
      patterns[40076] = 25'b10011100_10001010_00100110_1;
      patterns[40077] = 25'b10011100_10001011_00100111_1;
      patterns[40078] = 25'b10011100_10001100_00101000_1;
      patterns[40079] = 25'b10011100_10001101_00101001_1;
      patterns[40080] = 25'b10011100_10001110_00101010_1;
      patterns[40081] = 25'b10011100_10001111_00101011_1;
      patterns[40082] = 25'b10011100_10010000_00101100_1;
      patterns[40083] = 25'b10011100_10010001_00101101_1;
      patterns[40084] = 25'b10011100_10010010_00101110_1;
      patterns[40085] = 25'b10011100_10010011_00101111_1;
      patterns[40086] = 25'b10011100_10010100_00110000_1;
      patterns[40087] = 25'b10011100_10010101_00110001_1;
      patterns[40088] = 25'b10011100_10010110_00110010_1;
      patterns[40089] = 25'b10011100_10010111_00110011_1;
      patterns[40090] = 25'b10011100_10011000_00110100_1;
      patterns[40091] = 25'b10011100_10011001_00110101_1;
      patterns[40092] = 25'b10011100_10011010_00110110_1;
      patterns[40093] = 25'b10011100_10011011_00110111_1;
      patterns[40094] = 25'b10011100_10011100_00111000_1;
      patterns[40095] = 25'b10011100_10011101_00111001_1;
      patterns[40096] = 25'b10011100_10011110_00111010_1;
      patterns[40097] = 25'b10011100_10011111_00111011_1;
      patterns[40098] = 25'b10011100_10100000_00111100_1;
      patterns[40099] = 25'b10011100_10100001_00111101_1;
      patterns[40100] = 25'b10011100_10100010_00111110_1;
      patterns[40101] = 25'b10011100_10100011_00111111_1;
      patterns[40102] = 25'b10011100_10100100_01000000_1;
      patterns[40103] = 25'b10011100_10100101_01000001_1;
      patterns[40104] = 25'b10011100_10100110_01000010_1;
      patterns[40105] = 25'b10011100_10100111_01000011_1;
      patterns[40106] = 25'b10011100_10101000_01000100_1;
      patterns[40107] = 25'b10011100_10101001_01000101_1;
      patterns[40108] = 25'b10011100_10101010_01000110_1;
      patterns[40109] = 25'b10011100_10101011_01000111_1;
      patterns[40110] = 25'b10011100_10101100_01001000_1;
      patterns[40111] = 25'b10011100_10101101_01001001_1;
      patterns[40112] = 25'b10011100_10101110_01001010_1;
      patterns[40113] = 25'b10011100_10101111_01001011_1;
      patterns[40114] = 25'b10011100_10110000_01001100_1;
      patterns[40115] = 25'b10011100_10110001_01001101_1;
      patterns[40116] = 25'b10011100_10110010_01001110_1;
      patterns[40117] = 25'b10011100_10110011_01001111_1;
      patterns[40118] = 25'b10011100_10110100_01010000_1;
      patterns[40119] = 25'b10011100_10110101_01010001_1;
      patterns[40120] = 25'b10011100_10110110_01010010_1;
      patterns[40121] = 25'b10011100_10110111_01010011_1;
      patterns[40122] = 25'b10011100_10111000_01010100_1;
      patterns[40123] = 25'b10011100_10111001_01010101_1;
      patterns[40124] = 25'b10011100_10111010_01010110_1;
      patterns[40125] = 25'b10011100_10111011_01010111_1;
      patterns[40126] = 25'b10011100_10111100_01011000_1;
      patterns[40127] = 25'b10011100_10111101_01011001_1;
      patterns[40128] = 25'b10011100_10111110_01011010_1;
      patterns[40129] = 25'b10011100_10111111_01011011_1;
      patterns[40130] = 25'b10011100_11000000_01011100_1;
      patterns[40131] = 25'b10011100_11000001_01011101_1;
      patterns[40132] = 25'b10011100_11000010_01011110_1;
      patterns[40133] = 25'b10011100_11000011_01011111_1;
      patterns[40134] = 25'b10011100_11000100_01100000_1;
      patterns[40135] = 25'b10011100_11000101_01100001_1;
      patterns[40136] = 25'b10011100_11000110_01100010_1;
      patterns[40137] = 25'b10011100_11000111_01100011_1;
      patterns[40138] = 25'b10011100_11001000_01100100_1;
      patterns[40139] = 25'b10011100_11001001_01100101_1;
      patterns[40140] = 25'b10011100_11001010_01100110_1;
      patterns[40141] = 25'b10011100_11001011_01100111_1;
      patterns[40142] = 25'b10011100_11001100_01101000_1;
      patterns[40143] = 25'b10011100_11001101_01101001_1;
      patterns[40144] = 25'b10011100_11001110_01101010_1;
      patterns[40145] = 25'b10011100_11001111_01101011_1;
      patterns[40146] = 25'b10011100_11010000_01101100_1;
      patterns[40147] = 25'b10011100_11010001_01101101_1;
      patterns[40148] = 25'b10011100_11010010_01101110_1;
      patterns[40149] = 25'b10011100_11010011_01101111_1;
      patterns[40150] = 25'b10011100_11010100_01110000_1;
      patterns[40151] = 25'b10011100_11010101_01110001_1;
      patterns[40152] = 25'b10011100_11010110_01110010_1;
      patterns[40153] = 25'b10011100_11010111_01110011_1;
      patterns[40154] = 25'b10011100_11011000_01110100_1;
      patterns[40155] = 25'b10011100_11011001_01110101_1;
      patterns[40156] = 25'b10011100_11011010_01110110_1;
      patterns[40157] = 25'b10011100_11011011_01110111_1;
      patterns[40158] = 25'b10011100_11011100_01111000_1;
      patterns[40159] = 25'b10011100_11011101_01111001_1;
      patterns[40160] = 25'b10011100_11011110_01111010_1;
      patterns[40161] = 25'b10011100_11011111_01111011_1;
      patterns[40162] = 25'b10011100_11100000_01111100_1;
      patterns[40163] = 25'b10011100_11100001_01111101_1;
      patterns[40164] = 25'b10011100_11100010_01111110_1;
      patterns[40165] = 25'b10011100_11100011_01111111_1;
      patterns[40166] = 25'b10011100_11100100_10000000_1;
      patterns[40167] = 25'b10011100_11100101_10000001_1;
      patterns[40168] = 25'b10011100_11100110_10000010_1;
      patterns[40169] = 25'b10011100_11100111_10000011_1;
      patterns[40170] = 25'b10011100_11101000_10000100_1;
      patterns[40171] = 25'b10011100_11101001_10000101_1;
      patterns[40172] = 25'b10011100_11101010_10000110_1;
      patterns[40173] = 25'b10011100_11101011_10000111_1;
      patterns[40174] = 25'b10011100_11101100_10001000_1;
      patterns[40175] = 25'b10011100_11101101_10001001_1;
      patterns[40176] = 25'b10011100_11101110_10001010_1;
      patterns[40177] = 25'b10011100_11101111_10001011_1;
      patterns[40178] = 25'b10011100_11110000_10001100_1;
      patterns[40179] = 25'b10011100_11110001_10001101_1;
      patterns[40180] = 25'b10011100_11110010_10001110_1;
      patterns[40181] = 25'b10011100_11110011_10001111_1;
      patterns[40182] = 25'b10011100_11110100_10010000_1;
      patterns[40183] = 25'b10011100_11110101_10010001_1;
      patterns[40184] = 25'b10011100_11110110_10010010_1;
      patterns[40185] = 25'b10011100_11110111_10010011_1;
      patterns[40186] = 25'b10011100_11111000_10010100_1;
      patterns[40187] = 25'b10011100_11111001_10010101_1;
      patterns[40188] = 25'b10011100_11111010_10010110_1;
      patterns[40189] = 25'b10011100_11111011_10010111_1;
      patterns[40190] = 25'b10011100_11111100_10011000_1;
      patterns[40191] = 25'b10011100_11111101_10011001_1;
      patterns[40192] = 25'b10011100_11111110_10011010_1;
      patterns[40193] = 25'b10011100_11111111_10011011_1;
      patterns[40194] = 25'b10011101_00000000_10011101_0;
      patterns[40195] = 25'b10011101_00000001_10011110_0;
      patterns[40196] = 25'b10011101_00000010_10011111_0;
      patterns[40197] = 25'b10011101_00000011_10100000_0;
      patterns[40198] = 25'b10011101_00000100_10100001_0;
      patterns[40199] = 25'b10011101_00000101_10100010_0;
      patterns[40200] = 25'b10011101_00000110_10100011_0;
      patterns[40201] = 25'b10011101_00000111_10100100_0;
      patterns[40202] = 25'b10011101_00001000_10100101_0;
      patterns[40203] = 25'b10011101_00001001_10100110_0;
      patterns[40204] = 25'b10011101_00001010_10100111_0;
      patterns[40205] = 25'b10011101_00001011_10101000_0;
      patterns[40206] = 25'b10011101_00001100_10101001_0;
      patterns[40207] = 25'b10011101_00001101_10101010_0;
      patterns[40208] = 25'b10011101_00001110_10101011_0;
      patterns[40209] = 25'b10011101_00001111_10101100_0;
      patterns[40210] = 25'b10011101_00010000_10101101_0;
      patterns[40211] = 25'b10011101_00010001_10101110_0;
      patterns[40212] = 25'b10011101_00010010_10101111_0;
      patterns[40213] = 25'b10011101_00010011_10110000_0;
      patterns[40214] = 25'b10011101_00010100_10110001_0;
      patterns[40215] = 25'b10011101_00010101_10110010_0;
      patterns[40216] = 25'b10011101_00010110_10110011_0;
      patterns[40217] = 25'b10011101_00010111_10110100_0;
      patterns[40218] = 25'b10011101_00011000_10110101_0;
      patterns[40219] = 25'b10011101_00011001_10110110_0;
      patterns[40220] = 25'b10011101_00011010_10110111_0;
      patterns[40221] = 25'b10011101_00011011_10111000_0;
      patterns[40222] = 25'b10011101_00011100_10111001_0;
      patterns[40223] = 25'b10011101_00011101_10111010_0;
      patterns[40224] = 25'b10011101_00011110_10111011_0;
      patterns[40225] = 25'b10011101_00011111_10111100_0;
      patterns[40226] = 25'b10011101_00100000_10111101_0;
      patterns[40227] = 25'b10011101_00100001_10111110_0;
      patterns[40228] = 25'b10011101_00100010_10111111_0;
      patterns[40229] = 25'b10011101_00100011_11000000_0;
      patterns[40230] = 25'b10011101_00100100_11000001_0;
      patterns[40231] = 25'b10011101_00100101_11000010_0;
      patterns[40232] = 25'b10011101_00100110_11000011_0;
      patterns[40233] = 25'b10011101_00100111_11000100_0;
      patterns[40234] = 25'b10011101_00101000_11000101_0;
      patterns[40235] = 25'b10011101_00101001_11000110_0;
      patterns[40236] = 25'b10011101_00101010_11000111_0;
      patterns[40237] = 25'b10011101_00101011_11001000_0;
      patterns[40238] = 25'b10011101_00101100_11001001_0;
      patterns[40239] = 25'b10011101_00101101_11001010_0;
      patterns[40240] = 25'b10011101_00101110_11001011_0;
      patterns[40241] = 25'b10011101_00101111_11001100_0;
      patterns[40242] = 25'b10011101_00110000_11001101_0;
      patterns[40243] = 25'b10011101_00110001_11001110_0;
      patterns[40244] = 25'b10011101_00110010_11001111_0;
      patterns[40245] = 25'b10011101_00110011_11010000_0;
      patterns[40246] = 25'b10011101_00110100_11010001_0;
      patterns[40247] = 25'b10011101_00110101_11010010_0;
      patterns[40248] = 25'b10011101_00110110_11010011_0;
      patterns[40249] = 25'b10011101_00110111_11010100_0;
      patterns[40250] = 25'b10011101_00111000_11010101_0;
      patterns[40251] = 25'b10011101_00111001_11010110_0;
      patterns[40252] = 25'b10011101_00111010_11010111_0;
      patterns[40253] = 25'b10011101_00111011_11011000_0;
      patterns[40254] = 25'b10011101_00111100_11011001_0;
      patterns[40255] = 25'b10011101_00111101_11011010_0;
      patterns[40256] = 25'b10011101_00111110_11011011_0;
      patterns[40257] = 25'b10011101_00111111_11011100_0;
      patterns[40258] = 25'b10011101_01000000_11011101_0;
      patterns[40259] = 25'b10011101_01000001_11011110_0;
      patterns[40260] = 25'b10011101_01000010_11011111_0;
      patterns[40261] = 25'b10011101_01000011_11100000_0;
      patterns[40262] = 25'b10011101_01000100_11100001_0;
      patterns[40263] = 25'b10011101_01000101_11100010_0;
      patterns[40264] = 25'b10011101_01000110_11100011_0;
      patterns[40265] = 25'b10011101_01000111_11100100_0;
      patterns[40266] = 25'b10011101_01001000_11100101_0;
      patterns[40267] = 25'b10011101_01001001_11100110_0;
      patterns[40268] = 25'b10011101_01001010_11100111_0;
      patterns[40269] = 25'b10011101_01001011_11101000_0;
      patterns[40270] = 25'b10011101_01001100_11101001_0;
      patterns[40271] = 25'b10011101_01001101_11101010_0;
      patterns[40272] = 25'b10011101_01001110_11101011_0;
      patterns[40273] = 25'b10011101_01001111_11101100_0;
      patterns[40274] = 25'b10011101_01010000_11101101_0;
      patterns[40275] = 25'b10011101_01010001_11101110_0;
      patterns[40276] = 25'b10011101_01010010_11101111_0;
      patterns[40277] = 25'b10011101_01010011_11110000_0;
      patterns[40278] = 25'b10011101_01010100_11110001_0;
      patterns[40279] = 25'b10011101_01010101_11110010_0;
      patterns[40280] = 25'b10011101_01010110_11110011_0;
      patterns[40281] = 25'b10011101_01010111_11110100_0;
      patterns[40282] = 25'b10011101_01011000_11110101_0;
      patterns[40283] = 25'b10011101_01011001_11110110_0;
      patterns[40284] = 25'b10011101_01011010_11110111_0;
      patterns[40285] = 25'b10011101_01011011_11111000_0;
      patterns[40286] = 25'b10011101_01011100_11111001_0;
      patterns[40287] = 25'b10011101_01011101_11111010_0;
      patterns[40288] = 25'b10011101_01011110_11111011_0;
      patterns[40289] = 25'b10011101_01011111_11111100_0;
      patterns[40290] = 25'b10011101_01100000_11111101_0;
      patterns[40291] = 25'b10011101_01100001_11111110_0;
      patterns[40292] = 25'b10011101_01100010_11111111_0;
      patterns[40293] = 25'b10011101_01100011_00000000_1;
      patterns[40294] = 25'b10011101_01100100_00000001_1;
      patterns[40295] = 25'b10011101_01100101_00000010_1;
      patterns[40296] = 25'b10011101_01100110_00000011_1;
      patterns[40297] = 25'b10011101_01100111_00000100_1;
      patterns[40298] = 25'b10011101_01101000_00000101_1;
      patterns[40299] = 25'b10011101_01101001_00000110_1;
      patterns[40300] = 25'b10011101_01101010_00000111_1;
      patterns[40301] = 25'b10011101_01101011_00001000_1;
      patterns[40302] = 25'b10011101_01101100_00001001_1;
      patterns[40303] = 25'b10011101_01101101_00001010_1;
      patterns[40304] = 25'b10011101_01101110_00001011_1;
      patterns[40305] = 25'b10011101_01101111_00001100_1;
      patterns[40306] = 25'b10011101_01110000_00001101_1;
      patterns[40307] = 25'b10011101_01110001_00001110_1;
      patterns[40308] = 25'b10011101_01110010_00001111_1;
      patterns[40309] = 25'b10011101_01110011_00010000_1;
      patterns[40310] = 25'b10011101_01110100_00010001_1;
      patterns[40311] = 25'b10011101_01110101_00010010_1;
      patterns[40312] = 25'b10011101_01110110_00010011_1;
      patterns[40313] = 25'b10011101_01110111_00010100_1;
      patterns[40314] = 25'b10011101_01111000_00010101_1;
      patterns[40315] = 25'b10011101_01111001_00010110_1;
      patterns[40316] = 25'b10011101_01111010_00010111_1;
      patterns[40317] = 25'b10011101_01111011_00011000_1;
      patterns[40318] = 25'b10011101_01111100_00011001_1;
      patterns[40319] = 25'b10011101_01111101_00011010_1;
      patterns[40320] = 25'b10011101_01111110_00011011_1;
      patterns[40321] = 25'b10011101_01111111_00011100_1;
      patterns[40322] = 25'b10011101_10000000_00011101_1;
      patterns[40323] = 25'b10011101_10000001_00011110_1;
      patterns[40324] = 25'b10011101_10000010_00011111_1;
      patterns[40325] = 25'b10011101_10000011_00100000_1;
      patterns[40326] = 25'b10011101_10000100_00100001_1;
      patterns[40327] = 25'b10011101_10000101_00100010_1;
      patterns[40328] = 25'b10011101_10000110_00100011_1;
      patterns[40329] = 25'b10011101_10000111_00100100_1;
      patterns[40330] = 25'b10011101_10001000_00100101_1;
      patterns[40331] = 25'b10011101_10001001_00100110_1;
      patterns[40332] = 25'b10011101_10001010_00100111_1;
      patterns[40333] = 25'b10011101_10001011_00101000_1;
      patterns[40334] = 25'b10011101_10001100_00101001_1;
      patterns[40335] = 25'b10011101_10001101_00101010_1;
      patterns[40336] = 25'b10011101_10001110_00101011_1;
      patterns[40337] = 25'b10011101_10001111_00101100_1;
      patterns[40338] = 25'b10011101_10010000_00101101_1;
      patterns[40339] = 25'b10011101_10010001_00101110_1;
      patterns[40340] = 25'b10011101_10010010_00101111_1;
      patterns[40341] = 25'b10011101_10010011_00110000_1;
      patterns[40342] = 25'b10011101_10010100_00110001_1;
      patterns[40343] = 25'b10011101_10010101_00110010_1;
      patterns[40344] = 25'b10011101_10010110_00110011_1;
      patterns[40345] = 25'b10011101_10010111_00110100_1;
      patterns[40346] = 25'b10011101_10011000_00110101_1;
      patterns[40347] = 25'b10011101_10011001_00110110_1;
      patterns[40348] = 25'b10011101_10011010_00110111_1;
      patterns[40349] = 25'b10011101_10011011_00111000_1;
      patterns[40350] = 25'b10011101_10011100_00111001_1;
      patterns[40351] = 25'b10011101_10011101_00111010_1;
      patterns[40352] = 25'b10011101_10011110_00111011_1;
      patterns[40353] = 25'b10011101_10011111_00111100_1;
      patterns[40354] = 25'b10011101_10100000_00111101_1;
      patterns[40355] = 25'b10011101_10100001_00111110_1;
      patterns[40356] = 25'b10011101_10100010_00111111_1;
      patterns[40357] = 25'b10011101_10100011_01000000_1;
      patterns[40358] = 25'b10011101_10100100_01000001_1;
      patterns[40359] = 25'b10011101_10100101_01000010_1;
      patterns[40360] = 25'b10011101_10100110_01000011_1;
      patterns[40361] = 25'b10011101_10100111_01000100_1;
      patterns[40362] = 25'b10011101_10101000_01000101_1;
      patterns[40363] = 25'b10011101_10101001_01000110_1;
      patterns[40364] = 25'b10011101_10101010_01000111_1;
      patterns[40365] = 25'b10011101_10101011_01001000_1;
      patterns[40366] = 25'b10011101_10101100_01001001_1;
      patterns[40367] = 25'b10011101_10101101_01001010_1;
      patterns[40368] = 25'b10011101_10101110_01001011_1;
      patterns[40369] = 25'b10011101_10101111_01001100_1;
      patterns[40370] = 25'b10011101_10110000_01001101_1;
      patterns[40371] = 25'b10011101_10110001_01001110_1;
      patterns[40372] = 25'b10011101_10110010_01001111_1;
      patterns[40373] = 25'b10011101_10110011_01010000_1;
      patterns[40374] = 25'b10011101_10110100_01010001_1;
      patterns[40375] = 25'b10011101_10110101_01010010_1;
      patterns[40376] = 25'b10011101_10110110_01010011_1;
      patterns[40377] = 25'b10011101_10110111_01010100_1;
      patterns[40378] = 25'b10011101_10111000_01010101_1;
      patterns[40379] = 25'b10011101_10111001_01010110_1;
      patterns[40380] = 25'b10011101_10111010_01010111_1;
      patterns[40381] = 25'b10011101_10111011_01011000_1;
      patterns[40382] = 25'b10011101_10111100_01011001_1;
      patterns[40383] = 25'b10011101_10111101_01011010_1;
      patterns[40384] = 25'b10011101_10111110_01011011_1;
      patterns[40385] = 25'b10011101_10111111_01011100_1;
      patterns[40386] = 25'b10011101_11000000_01011101_1;
      patterns[40387] = 25'b10011101_11000001_01011110_1;
      patterns[40388] = 25'b10011101_11000010_01011111_1;
      patterns[40389] = 25'b10011101_11000011_01100000_1;
      patterns[40390] = 25'b10011101_11000100_01100001_1;
      patterns[40391] = 25'b10011101_11000101_01100010_1;
      patterns[40392] = 25'b10011101_11000110_01100011_1;
      patterns[40393] = 25'b10011101_11000111_01100100_1;
      patterns[40394] = 25'b10011101_11001000_01100101_1;
      patterns[40395] = 25'b10011101_11001001_01100110_1;
      patterns[40396] = 25'b10011101_11001010_01100111_1;
      patterns[40397] = 25'b10011101_11001011_01101000_1;
      patterns[40398] = 25'b10011101_11001100_01101001_1;
      patterns[40399] = 25'b10011101_11001101_01101010_1;
      patterns[40400] = 25'b10011101_11001110_01101011_1;
      patterns[40401] = 25'b10011101_11001111_01101100_1;
      patterns[40402] = 25'b10011101_11010000_01101101_1;
      patterns[40403] = 25'b10011101_11010001_01101110_1;
      patterns[40404] = 25'b10011101_11010010_01101111_1;
      patterns[40405] = 25'b10011101_11010011_01110000_1;
      patterns[40406] = 25'b10011101_11010100_01110001_1;
      patterns[40407] = 25'b10011101_11010101_01110010_1;
      patterns[40408] = 25'b10011101_11010110_01110011_1;
      patterns[40409] = 25'b10011101_11010111_01110100_1;
      patterns[40410] = 25'b10011101_11011000_01110101_1;
      patterns[40411] = 25'b10011101_11011001_01110110_1;
      patterns[40412] = 25'b10011101_11011010_01110111_1;
      patterns[40413] = 25'b10011101_11011011_01111000_1;
      patterns[40414] = 25'b10011101_11011100_01111001_1;
      patterns[40415] = 25'b10011101_11011101_01111010_1;
      patterns[40416] = 25'b10011101_11011110_01111011_1;
      patterns[40417] = 25'b10011101_11011111_01111100_1;
      patterns[40418] = 25'b10011101_11100000_01111101_1;
      patterns[40419] = 25'b10011101_11100001_01111110_1;
      patterns[40420] = 25'b10011101_11100010_01111111_1;
      patterns[40421] = 25'b10011101_11100011_10000000_1;
      patterns[40422] = 25'b10011101_11100100_10000001_1;
      patterns[40423] = 25'b10011101_11100101_10000010_1;
      patterns[40424] = 25'b10011101_11100110_10000011_1;
      patterns[40425] = 25'b10011101_11100111_10000100_1;
      patterns[40426] = 25'b10011101_11101000_10000101_1;
      patterns[40427] = 25'b10011101_11101001_10000110_1;
      patterns[40428] = 25'b10011101_11101010_10000111_1;
      patterns[40429] = 25'b10011101_11101011_10001000_1;
      patterns[40430] = 25'b10011101_11101100_10001001_1;
      patterns[40431] = 25'b10011101_11101101_10001010_1;
      patterns[40432] = 25'b10011101_11101110_10001011_1;
      patterns[40433] = 25'b10011101_11101111_10001100_1;
      patterns[40434] = 25'b10011101_11110000_10001101_1;
      patterns[40435] = 25'b10011101_11110001_10001110_1;
      patterns[40436] = 25'b10011101_11110010_10001111_1;
      patterns[40437] = 25'b10011101_11110011_10010000_1;
      patterns[40438] = 25'b10011101_11110100_10010001_1;
      patterns[40439] = 25'b10011101_11110101_10010010_1;
      patterns[40440] = 25'b10011101_11110110_10010011_1;
      patterns[40441] = 25'b10011101_11110111_10010100_1;
      patterns[40442] = 25'b10011101_11111000_10010101_1;
      patterns[40443] = 25'b10011101_11111001_10010110_1;
      patterns[40444] = 25'b10011101_11111010_10010111_1;
      patterns[40445] = 25'b10011101_11111011_10011000_1;
      patterns[40446] = 25'b10011101_11111100_10011001_1;
      patterns[40447] = 25'b10011101_11111101_10011010_1;
      patterns[40448] = 25'b10011101_11111110_10011011_1;
      patterns[40449] = 25'b10011101_11111111_10011100_1;
      patterns[40450] = 25'b10011110_00000000_10011110_0;
      patterns[40451] = 25'b10011110_00000001_10011111_0;
      patterns[40452] = 25'b10011110_00000010_10100000_0;
      patterns[40453] = 25'b10011110_00000011_10100001_0;
      patterns[40454] = 25'b10011110_00000100_10100010_0;
      patterns[40455] = 25'b10011110_00000101_10100011_0;
      patterns[40456] = 25'b10011110_00000110_10100100_0;
      patterns[40457] = 25'b10011110_00000111_10100101_0;
      patterns[40458] = 25'b10011110_00001000_10100110_0;
      patterns[40459] = 25'b10011110_00001001_10100111_0;
      patterns[40460] = 25'b10011110_00001010_10101000_0;
      patterns[40461] = 25'b10011110_00001011_10101001_0;
      patterns[40462] = 25'b10011110_00001100_10101010_0;
      patterns[40463] = 25'b10011110_00001101_10101011_0;
      patterns[40464] = 25'b10011110_00001110_10101100_0;
      patterns[40465] = 25'b10011110_00001111_10101101_0;
      patterns[40466] = 25'b10011110_00010000_10101110_0;
      patterns[40467] = 25'b10011110_00010001_10101111_0;
      patterns[40468] = 25'b10011110_00010010_10110000_0;
      patterns[40469] = 25'b10011110_00010011_10110001_0;
      patterns[40470] = 25'b10011110_00010100_10110010_0;
      patterns[40471] = 25'b10011110_00010101_10110011_0;
      patterns[40472] = 25'b10011110_00010110_10110100_0;
      patterns[40473] = 25'b10011110_00010111_10110101_0;
      patterns[40474] = 25'b10011110_00011000_10110110_0;
      patterns[40475] = 25'b10011110_00011001_10110111_0;
      patterns[40476] = 25'b10011110_00011010_10111000_0;
      patterns[40477] = 25'b10011110_00011011_10111001_0;
      patterns[40478] = 25'b10011110_00011100_10111010_0;
      patterns[40479] = 25'b10011110_00011101_10111011_0;
      patterns[40480] = 25'b10011110_00011110_10111100_0;
      patterns[40481] = 25'b10011110_00011111_10111101_0;
      patterns[40482] = 25'b10011110_00100000_10111110_0;
      patterns[40483] = 25'b10011110_00100001_10111111_0;
      patterns[40484] = 25'b10011110_00100010_11000000_0;
      patterns[40485] = 25'b10011110_00100011_11000001_0;
      patterns[40486] = 25'b10011110_00100100_11000010_0;
      patterns[40487] = 25'b10011110_00100101_11000011_0;
      patterns[40488] = 25'b10011110_00100110_11000100_0;
      patterns[40489] = 25'b10011110_00100111_11000101_0;
      patterns[40490] = 25'b10011110_00101000_11000110_0;
      patterns[40491] = 25'b10011110_00101001_11000111_0;
      patterns[40492] = 25'b10011110_00101010_11001000_0;
      patterns[40493] = 25'b10011110_00101011_11001001_0;
      patterns[40494] = 25'b10011110_00101100_11001010_0;
      patterns[40495] = 25'b10011110_00101101_11001011_0;
      patterns[40496] = 25'b10011110_00101110_11001100_0;
      patterns[40497] = 25'b10011110_00101111_11001101_0;
      patterns[40498] = 25'b10011110_00110000_11001110_0;
      patterns[40499] = 25'b10011110_00110001_11001111_0;
      patterns[40500] = 25'b10011110_00110010_11010000_0;
      patterns[40501] = 25'b10011110_00110011_11010001_0;
      patterns[40502] = 25'b10011110_00110100_11010010_0;
      patterns[40503] = 25'b10011110_00110101_11010011_0;
      patterns[40504] = 25'b10011110_00110110_11010100_0;
      patterns[40505] = 25'b10011110_00110111_11010101_0;
      patterns[40506] = 25'b10011110_00111000_11010110_0;
      patterns[40507] = 25'b10011110_00111001_11010111_0;
      patterns[40508] = 25'b10011110_00111010_11011000_0;
      patterns[40509] = 25'b10011110_00111011_11011001_0;
      patterns[40510] = 25'b10011110_00111100_11011010_0;
      patterns[40511] = 25'b10011110_00111101_11011011_0;
      patterns[40512] = 25'b10011110_00111110_11011100_0;
      patterns[40513] = 25'b10011110_00111111_11011101_0;
      patterns[40514] = 25'b10011110_01000000_11011110_0;
      patterns[40515] = 25'b10011110_01000001_11011111_0;
      patterns[40516] = 25'b10011110_01000010_11100000_0;
      patterns[40517] = 25'b10011110_01000011_11100001_0;
      patterns[40518] = 25'b10011110_01000100_11100010_0;
      patterns[40519] = 25'b10011110_01000101_11100011_0;
      patterns[40520] = 25'b10011110_01000110_11100100_0;
      patterns[40521] = 25'b10011110_01000111_11100101_0;
      patterns[40522] = 25'b10011110_01001000_11100110_0;
      patterns[40523] = 25'b10011110_01001001_11100111_0;
      patterns[40524] = 25'b10011110_01001010_11101000_0;
      patterns[40525] = 25'b10011110_01001011_11101001_0;
      patterns[40526] = 25'b10011110_01001100_11101010_0;
      patterns[40527] = 25'b10011110_01001101_11101011_0;
      patterns[40528] = 25'b10011110_01001110_11101100_0;
      patterns[40529] = 25'b10011110_01001111_11101101_0;
      patterns[40530] = 25'b10011110_01010000_11101110_0;
      patterns[40531] = 25'b10011110_01010001_11101111_0;
      patterns[40532] = 25'b10011110_01010010_11110000_0;
      patterns[40533] = 25'b10011110_01010011_11110001_0;
      patterns[40534] = 25'b10011110_01010100_11110010_0;
      patterns[40535] = 25'b10011110_01010101_11110011_0;
      patterns[40536] = 25'b10011110_01010110_11110100_0;
      patterns[40537] = 25'b10011110_01010111_11110101_0;
      patterns[40538] = 25'b10011110_01011000_11110110_0;
      patterns[40539] = 25'b10011110_01011001_11110111_0;
      patterns[40540] = 25'b10011110_01011010_11111000_0;
      patterns[40541] = 25'b10011110_01011011_11111001_0;
      patterns[40542] = 25'b10011110_01011100_11111010_0;
      patterns[40543] = 25'b10011110_01011101_11111011_0;
      patterns[40544] = 25'b10011110_01011110_11111100_0;
      patterns[40545] = 25'b10011110_01011111_11111101_0;
      patterns[40546] = 25'b10011110_01100000_11111110_0;
      patterns[40547] = 25'b10011110_01100001_11111111_0;
      patterns[40548] = 25'b10011110_01100010_00000000_1;
      patterns[40549] = 25'b10011110_01100011_00000001_1;
      patterns[40550] = 25'b10011110_01100100_00000010_1;
      patterns[40551] = 25'b10011110_01100101_00000011_1;
      patterns[40552] = 25'b10011110_01100110_00000100_1;
      patterns[40553] = 25'b10011110_01100111_00000101_1;
      patterns[40554] = 25'b10011110_01101000_00000110_1;
      patterns[40555] = 25'b10011110_01101001_00000111_1;
      patterns[40556] = 25'b10011110_01101010_00001000_1;
      patterns[40557] = 25'b10011110_01101011_00001001_1;
      patterns[40558] = 25'b10011110_01101100_00001010_1;
      patterns[40559] = 25'b10011110_01101101_00001011_1;
      patterns[40560] = 25'b10011110_01101110_00001100_1;
      patterns[40561] = 25'b10011110_01101111_00001101_1;
      patterns[40562] = 25'b10011110_01110000_00001110_1;
      patterns[40563] = 25'b10011110_01110001_00001111_1;
      patterns[40564] = 25'b10011110_01110010_00010000_1;
      patterns[40565] = 25'b10011110_01110011_00010001_1;
      patterns[40566] = 25'b10011110_01110100_00010010_1;
      patterns[40567] = 25'b10011110_01110101_00010011_1;
      patterns[40568] = 25'b10011110_01110110_00010100_1;
      patterns[40569] = 25'b10011110_01110111_00010101_1;
      patterns[40570] = 25'b10011110_01111000_00010110_1;
      patterns[40571] = 25'b10011110_01111001_00010111_1;
      patterns[40572] = 25'b10011110_01111010_00011000_1;
      patterns[40573] = 25'b10011110_01111011_00011001_1;
      patterns[40574] = 25'b10011110_01111100_00011010_1;
      patterns[40575] = 25'b10011110_01111101_00011011_1;
      patterns[40576] = 25'b10011110_01111110_00011100_1;
      patterns[40577] = 25'b10011110_01111111_00011101_1;
      patterns[40578] = 25'b10011110_10000000_00011110_1;
      patterns[40579] = 25'b10011110_10000001_00011111_1;
      patterns[40580] = 25'b10011110_10000010_00100000_1;
      patterns[40581] = 25'b10011110_10000011_00100001_1;
      patterns[40582] = 25'b10011110_10000100_00100010_1;
      patterns[40583] = 25'b10011110_10000101_00100011_1;
      patterns[40584] = 25'b10011110_10000110_00100100_1;
      patterns[40585] = 25'b10011110_10000111_00100101_1;
      patterns[40586] = 25'b10011110_10001000_00100110_1;
      patterns[40587] = 25'b10011110_10001001_00100111_1;
      patterns[40588] = 25'b10011110_10001010_00101000_1;
      patterns[40589] = 25'b10011110_10001011_00101001_1;
      patterns[40590] = 25'b10011110_10001100_00101010_1;
      patterns[40591] = 25'b10011110_10001101_00101011_1;
      patterns[40592] = 25'b10011110_10001110_00101100_1;
      patterns[40593] = 25'b10011110_10001111_00101101_1;
      patterns[40594] = 25'b10011110_10010000_00101110_1;
      patterns[40595] = 25'b10011110_10010001_00101111_1;
      patterns[40596] = 25'b10011110_10010010_00110000_1;
      patterns[40597] = 25'b10011110_10010011_00110001_1;
      patterns[40598] = 25'b10011110_10010100_00110010_1;
      patterns[40599] = 25'b10011110_10010101_00110011_1;
      patterns[40600] = 25'b10011110_10010110_00110100_1;
      patterns[40601] = 25'b10011110_10010111_00110101_1;
      patterns[40602] = 25'b10011110_10011000_00110110_1;
      patterns[40603] = 25'b10011110_10011001_00110111_1;
      patterns[40604] = 25'b10011110_10011010_00111000_1;
      patterns[40605] = 25'b10011110_10011011_00111001_1;
      patterns[40606] = 25'b10011110_10011100_00111010_1;
      patterns[40607] = 25'b10011110_10011101_00111011_1;
      patterns[40608] = 25'b10011110_10011110_00111100_1;
      patterns[40609] = 25'b10011110_10011111_00111101_1;
      patterns[40610] = 25'b10011110_10100000_00111110_1;
      patterns[40611] = 25'b10011110_10100001_00111111_1;
      patterns[40612] = 25'b10011110_10100010_01000000_1;
      patterns[40613] = 25'b10011110_10100011_01000001_1;
      patterns[40614] = 25'b10011110_10100100_01000010_1;
      patterns[40615] = 25'b10011110_10100101_01000011_1;
      patterns[40616] = 25'b10011110_10100110_01000100_1;
      patterns[40617] = 25'b10011110_10100111_01000101_1;
      patterns[40618] = 25'b10011110_10101000_01000110_1;
      patterns[40619] = 25'b10011110_10101001_01000111_1;
      patterns[40620] = 25'b10011110_10101010_01001000_1;
      patterns[40621] = 25'b10011110_10101011_01001001_1;
      patterns[40622] = 25'b10011110_10101100_01001010_1;
      patterns[40623] = 25'b10011110_10101101_01001011_1;
      patterns[40624] = 25'b10011110_10101110_01001100_1;
      patterns[40625] = 25'b10011110_10101111_01001101_1;
      patterns[40626] = 25'b10011110_10110000_01001110_1;
      patterns[40627] = 25'b10011110_10110001_01001111_1;
      patterns[40628] = 25'b10011110_10110010_01010000_1;
      patterns[40629] = 25'b10011110_10110011_01010001_1;
      patterns[40630] = 25'b10011110_10110100_01010010_1;
      patterns[40631] = 25'b10011110_10110101_01010011_1;
      patterns[40632] = 25'b10011110_10110110_01010100_1;
      patterns[40633] = 25'b10011110_10110111_01010101_1;
      patterns[40634] = 25'b10011110_10111000_01010110_1;
      patterns[40635] = 25'b10011110_10111001_01010111_1;
      patterns[40636] = 25'b10011110_10111010_01011000_1;
      patterns[40637] = 25'b10011110_10111011_01011001_1;
      patterns[40638] = 25'b10011110_10111100_01011010_1;
      patterns[40639] = 25'b10011110_10111101_01011011_1;
      patterns[40640] = 25'b10011110_10111110_01011100_1;
      patterns[40641] = 25'b10011110_10111111_01011101_1;
      patterns[40642] = 25'b10011110_11000000_01011110_1;
      patterns[40643] = 25'b10011110_11000001_01011111_1;
      patterns[40644] = 25'b10011110_11000010_01100000_1;
      patterns[40645] = 25'b10011110_11000011_01100001_1;
      patterns[40646] = 25'b10011110_11000100_01100010_1;
      patterns[40647] = 25'b10011110_11000101_01100011_1;
      patterns[40648] = 25'b10011110_11000110_01100100_1;
      patterns[40649] = 25'b10011110_11000111_01100101_1;
      patterns[40650] = 25'b10011110_11001000_01100110_1;
      patterns[40651] = 25'b10011110_11001001_01100111_1;
      patterns[40652] = 25'b10011110_11001010_01101000_1;
      patterns[40653] = 25'b10011110_11001011_01101001_1;
      patterns[40654] = 25'b10011110_11001100_01101010_1;
      patterns[40655] = 25'b10011110_11001101_01101011_1;
      patterns[40656] = 25'b10011110_11001110_01101100_1;
      patterns[40657] = 25'b10011110_11001111_01101101_1;
      patterns[40658] = 25'b10011110_11010000_01101110_1;
      patterns[40659] = 25'b10011110_11010001_01101111_1;
      patterns[40660] = 25'b10011110_11010010_01110000_1;
      patterns[40661] = 25'b10011110_11010011_01110001_1;
      patterns[40662] = 25'b10011110_11010100_01110010_1;
      patterns[40663] = 25'b10011110_11010101_01110011_1;
      patterns[40664] = 25'b10011110_11010110_01110100_1;
      patterns[40665] = 25'b10011110_11010111_01110101_1;
      patterns[40666] = 25'b10011110_11011000_01110110_1;
      patterns[40667] = 25'b10011110_11011001_01110111_1;
      patterns[40668] = 25'b10011110_11011010_01111000_1;
      patterns[40669] = 25'b10011110_11011011_01111001_1;
      patterns[40670] = 25'b10011110_11011100_01111010_1;
      patterns[40671] = 25'b10011110_11011101_01111011_1;
      patterns[40672] = 25'b10011110_11011110_01111100_1;
      patterns[40673] = 25'b10011110_11011111_01111101_1;
      patterns[40674] = 25'b10011110_11100000_01111110_1;
      patterns[40675] = 25'b10011110_11100001_01111111_1;
      patterns[40676] = 25'b10011110_11100010_10000000_1;
      patterns[40677] = 25'b10011110_11100011_10000001_1;
      patterns[40678] = 25'b10011110_11100100_10000010_1;
      patterns[40679] = 25'b10011110_11100101_10000011_1;
      patterns[40680] = 25'b10011110_11100110_10000100_1;
      patterns[40681] = 25'b10011110_11100111_10000101_1;
      patterns[40682] = 25'b10011110_11101000_10000110_1;
      patterns[40683] = 25'b10011110_11101001_10000111_1;
      patterns[40684] = 25'b10011110_11101010_10001000_1;
      patterns[40685] = 25'b10011110_11101011_10001001_1;
      patterns[40686] = 25'b10011110_11101100_10001010_1;
      patterns[40687] = 25'b10011110_11101101_10001011_1;
      patterns[40688] = 25'b10011110_11101110_10001100_1;
      patterns[40689] = 25'b10011110_11101111_10001101_1;
      patterns[40690] = 25'b10011110_11110000_10001110_1;
      patterns[40691] = 25'b10011110_11110001_10001111_1;
      patterns[40692] = 25'b10011110_11110010_10010000_1;
      patterns[40693] = 25'b10011110_11110011_10010001_1;
      patterns[40694] = 25'b10011110_11110100_10010010_1;
      patterns[40695] = 25'b10011110_11110101_10010011_1;
      patterns[40696] = 25'b10011110_11110110_10010100_1;
      patterns[40697] = 25'b10011110_11110111_10010101_1;
      patterns[40698] = 25'b10011110_11111000_10010110_1;
      patterns[40699] = 25'b10011110_11111001_10010111_1;
      patterns[40700] = 25'b10011110_11111010_10011000_1;
      patterns[40701] = 25'b10011110_11111011_10011001_1;
      patterns[40702] = 25'b10011110_11111100_10011010_1;
      patterns[40703] = 25'b10011110_11111101_10011011_1;
      patterns[40704] = 25'b10011110_11111110_10011100_1;
      patterns[40705] = 25'b10011110_11111111_10011101_1;
      patterns[40706] = 25'b10011111_00000000_10011111_0;
      patterns[40707] = 25'b10011111_00000001_10100000_0;
      patterns[40708] = 25'b10011111_00000010_10100001_0;
      patterns[40709] = 25'b10011111_00000011_10100010_0;
      patterns[40710] = 25'b10011111_00000100_10100011_0;
      patterns[40711] = 25'b10011111_00000101_10100100_0;
      patterns[40712] = 25'b10011111_00000110_10100101_0;
      patterns[40713] = 25'b10011111_00000111_10100110_0;
      patterns[40714] = 25'b10011111_00001000_10100111_0;
      patterns[40715] = 25'b10011111_00001001_10101000_0;
      patterns[40716] = 25'b10011111_00001010_10101001_0;
      patterns[40717] = 25'b10011111_00001011_10101010_0;
      patterns[40718] = 25'b10011111_00001100_10101011_0;
      patterns[40719] = 25'b10011111_00001101_10101100_0;
      patterns[40720] = 25'b10011111_00001110_10101101_0;
      patterns[40721] = 25'b10011111_00001111_10101110_0;
      patterns[40722] = 25'b10011111_00010000_10101111_0;
      patterns[40723] = 25'b10011111_00010001_10110000_0;
      patterns[40724] = 25'b10011111_00010010_10110001_0;
      patterns[40725] = 25'b10011111_00010011_10110010_0;
      patterns[40726] = 25'b10011111_00010100_10110011_0;
      patterns[40727] = 25'b10011111_00010101_10110100_0;
      patterns[40728] = 25'b10011111_00010110_10110101_0;
      patterns[40729] = 25'b10011111_00010111_10110110_0;
      patterns[40730] = 25'b10011111_00011000_10110111_0;
      patterns[40731] = 25'b10011111_00011001_10111000_0;
      patterns[40732] = 25'b10011111_00011010_10111001_0;
      patterns[40733] = 25'b10011111_00011011_10111010_0;
      patterns[40734] = 25'b10011111_00011100_10111011_0;
      patterns[40735] = 25'b10011111_00011101_10111100_0;
      patterns[40736] = 25'b10011111_00011110_10111101_0;
      patterns[40737] = 25'b10011111_00011111_10111110_0;
      patterns[40738] = 25'b10011111_00100000_10111111_0;
      patterns[40739] = 25'b10011111_00100001_11000000_0;
      patterns[40740] = 25'b10011111_00100010_11000001_0;
      patterns[40741] = 25'b10011111_00100011_11000010_0;
      patterns[40742] = 25'b10011111_00100100_11000011_0;
      patterns[40743] = 25'b10011111_00100101_11000100_0;
      patterns[40744] = 25'b10011111_00100110_11000101_0;
      patterns[40745] = 25'b10011111_00100111_11000110_0;
      patterns[40746] = 25'b10011111_00101000_11000111_0;
      patterns[40747] = 25'b10011111_00101001_11001000_0;
      patterns[40748] = 25'b10011111_00101010_11001001_0;
      patterns[40749] = 25'b10011111_00101011_11001010_0;
      patterns[40750] = 25'b10011111_00101100_11001011_0;
      patterns[40751] = 25'b10011111_00101101_11001100_0;
      patterns[40752] = 25'b10011111_00101110_11001101_0;
      patterns[40753] = 25'b10011111_00101111_11001110_0;
      patterns[40754] = 25'b10011111_00110000_11001111_0;
      patterns[40755] = 25'b10011111_00110001_11010000_0;
      patterns[40756] = 25'b10011111_00110010_11010001_0;
      patterns[40757] = 25'b10011111_00110011_11010010_0;
      patterns[40758] = 25'b10011111_00110100_11010011_0;
      patterns[40759] = 25'b10011111_00110101_11010100_0;
      patterns[40760] = 25'b10011111_00110110_11010101_0;
      patterns[40761] = 25'b10011111_00110111_11010110_0;
      patterns[40762] = 25'b10011111_00111000_11010111_0;
      patterns[40763] = 25'b10011111_00111001_11011000_0;
      patterns[40764] = 25'b10011111_00111010_11011001_0;
      patterns[40765] = 25'b10011111_00111011_11011010_0;
      patterns[40766] = 25'b10011111_00111100_11011011_0;
      patterns[40767] = 25'b10011111_00111101_11011100_0;
      patterns[40768] = 25'b10011111_00111110_11011101_0;
      patterns[40769] = 25'b10011111_00111111_11011110_0;
      patterns[40770] = 25'b10011111_01000000_11011111_0;
      patterns[40771] = 25'b10011111_01000001_11100000_0;
      patterns[40772] = 25'b10011111_01000010_11100001_0;
      patterns[40773] = 25'b10011111_01000011_11100010_0;
      patterns[40774] = 25'b10011111_01000100_11100011_0;
      patterns[40775] = 25'b10011111_01000101_11100100_0;
      patterns[40776] = 25'b10011111_01000110_11100101_0;
      patterns[40777] = 25'b10011111_01000111_11100110_0;
      patterns[40778] = 25'b10011111_01001000_11100111_0;
      patterns[40779] = 25'b10011111_01001001_11101000_0;
      patterns[40780] = 25'b10011111_01001010_11101001_0;
      patterns[40781] = 25'b10011111_01001011_11101010_0;
      patterns[40782] = 25'b10011111_01001100_11101011_0;
      patterns[40783] = 25'b10011111_01001101_11101100_0;
      patterns[40784] = 25'b10011111_01001110_11101101_0;
      patterns[40785] = 25'b10011111_01001111_11101110_0;
      patterns[40786] = 25'b10011111_01010000_11101111_0;
      patterns[40787] = 25'b10011111_01010001_11110000_0;
      patterns[40788] = 25'b10011111_01010010_11110001_0;
      patterns[40789] = 25'b10011111_01010011_11110010_0;
      patterns[40790] = 25'b10011111_01010100_11110011_0;
      patterns[40791] = 25'b10011111_01010101_11110100_0;
      patterns[40792] = 25'b10011111_01010110_11110101_0;
      patterns[40793] = 25'b10011111_01010111_11110110_0;
      patterns[40794] = 25'b10011111_01011000_11110111_0;
      patterns[40795] = 25'b10011111_01011001_11111000_0;
      patterns[40796] = 25'b10011111_01011010_11111001_0;
      patterns[40797] = 25'b10011111_01011011_11111010_0;
      patterns[40798] = 25'b10011111_01011100_11111011_0;
      patterns[40799] = 25'b10011111_01011101_11111100_0;
      patterns[40800] = 25'b10011111_01011110_11111101_0;
      patterns[40801] = 25'b10011111_01011111_11111110_0;
      patterns[40802] = 25'b10011111_01100000_11111111_0;
      patterns[40803] = 25'b10011111_01100001_00000000_1;
      patterns[40804] = 25'b10011111_01100010_00000001_1;
      patterns[40805] = 25'b10011111_01100011_00000010_1;
      patterns[40806] = 25'b10011111_01100100_00000011_1;
      patterns[40807] = 25'b10011111_01100101_00000100_1;
      patterns[40808] = 25'b10011111_01100110_00000101_1;
      patterns[40809] = 25'b10011111_01100111_00000110_1;
      patterns[40810] = 25'b10011111_01101000_00000111_1;
      patterns[40811] = 25'b10011111_01101001_00001000_1;
      patterns[40812] = 25'b10011111_01101010_00001001_1;
      patterns[40813] = 25'b10011111_01101011_00001010_1;
      patterns[40814] = 25'b10011111_01101100_00001011_1;
      patterns[40815] = 25'b10011111_01101101_00001100_1;
      patterns[40816] = 25'b10011111_01101110_00001101_1;
      patterns[40817] = 25'b10011111_01101111_00001110_1;
      patterns[40818] = 25'b10011111_01110000_00001111_1;
      patterns[40819] = 25'b10011111_01110001_00010000_1;
      patterns[40820] = 25'b10011111_01110010_00010001_1;
      patterns[40821] = 25'b10011111_01110011_00010010_1;
      patterns[40822] = 25'b10011111_01110100_00010011_1;
      patterns[40823] = 25'b10011111_01110101_00010100_1;
      patterns[40824] = 25'b10011111_01110110_00010101_1;
      patterns[40825] = 25'b10011111_01110111_00010110_1;
      patterns[40826] = 25'b10011111_01111000_00010111_1;
      patterns[40827] = 25'b10011111_01111001_00011000_1;
      patterns[40828] = 25'b10011111_01111010_00011001_1;
      patterns[40829] = 25'b10011111_01111011_00011010_1;
      patterns[40830] = 25'b10011111_01111100_00011011_1;
      patterns[40831] = 25'b10011111_01111101_00011100_1;
      patterns[40832] = 25'b10011111_01111110_00011101_1;
      patterns[40833] = 25'b10011111_01111111_00011110_1;
      patterns[40834] = 25'b10011111_10000000_00011111_1;
      patterns[40835] = 25'b10011111_10000001_00100000_1;
      patterns[40836] = 25'b10011111_10000010_00100001_1;
      patterns[40837] = 25'b10011111_10000011_00100010_1;
      patterns[40838] = 25'b10011111_10000100_00100011_1;
      patterns[40839] = 25'b10011111_10000101_00100100_1;
      patterns[40840] = 25'b10011111_10000110_00100101_1;
      patterns[40841] = 25'b10011111_10000111_00100110_1;
      patterns[40842] = 25'b10011111_10001000_00100111_1;
      patterns[40843] = 25'b10011111_10001001_00101000_1;
      patterns[40844] = 25'b10011111_10001010_00101001_1;
      patterns[40845] = 25'b10011111_10001011_00101010_1;
      patterns[40846] = 25'b10011111_10001100_00101011_1;
      patterns[40847] = 25'b10011111_10001101_00101100_1;
      patterns[40848] = 25'b10011111_10001110_00101101_1;
      patterns[40849] = 25'b10011111_10001111_00101110_1;
      patterns[40850] = 25'b10011111_10010000_00101111_1;
      patterns[40851] = 25'b10011111_10010001_00110000_1;
      patterns[40852] = 25'b10011111_10010010_00110001_1;
      patterns[40853] = 25'b10011111_10010011_00110010_1;
      patterns[40854] = 25'b10011111_10010100_00110011_1;
      patterns[40855] = 25'b10011111_10010101_00110100_1;
      patterns[40856] = 25'b10011111_10010110_00110101_1;
      patterns[40857] = 25'b10011111_10010111_00110110_1;
      patterns[40858] = 25'b10011111_10011000_00110111_1;
      patterns[40859] = 25'b10011111_10011001_00111000_1;
      patterns[40860] = 25'b10011111_10011010_00111001_1;
      patterns[40861] = 25'b10011111_10011011_00111010_1;
      patterns[40862] = 25'b10011111_10011100_00111011_1;
      patterns[40863] = 25'b10011111_10011101_00111100_1;
      patterns[40864] = 25'b10011111_10011110_00111101_1;
      patterns[40865] = 25'b10011111_10011111_00111110_1;
      patterns[40866] = 25'b10011111_10100000_00111111_1;
      patterns[40867] = 25'b10011111_10100001_01000000_1;
      patterns[40868] = 25'b10011111_10100010_01000001_1;
      patterns[40869] = 25'b10011111_10100011_01000010_1;
      patterns[40870] = 25'b10011111_10100100_01000011_1;
      patterns[40871] = 25'b10011111_10100101_01000100_1;
      patterns[40872] = 25'b10011111_10100110_01000101_1;
      patterns[40873] = 25'b10011111_10100111_01000110_1;
      patterns[40874] = 25'b10011111_10101000_01000111_1;
      patterns[40875] = 25'b10011111_10101001_01001000_1;
      patterns[40876] = 25'b10011111_10101010_01001001_1;
      patterns[40877] = 25'b10011111_10101011_01001010_1;
      patterns[40878] = 25'b10011111_10101100_01001011_1;
      patterns[40879] = 25'b10011111_10101101_01001100_1;
      patterns[40880] = 25'b10011111_10101110_01001101_1;
      patterns[40881] = 25'b10011111_10101111_01001110_1;
      patterns[40882] = 25'b10011111_10110000_01001111_1;
      patterns[40883] = 25'b10011111_10110001_01010000_1;
      patterns[40884] = 25'b10011111_10110010_01010001_1;
      patterns[40885] = 25'b10011111_10110011_01010010_1;
      patterns[40886] = 25'b10011111_10110100_01010011_1;
      patterns[40887] = 25'b10011111_10110101_01010100_1;
      patterns[40888] = 25'b10011111_10110110_01010101_1;
      patterns[40889] = 25'b10011111_10110111_01010110_1;
      patterns[40890] = 25'b10011111_10111000_01010111_1;
      patterns[40891] = 25'b10011111_10111001_01011000_1;
      patterns[40892] = 25'b10011111_10111010_01011001_1;
      patterns[40893] = 25'b10011111_10111011_01011010_1;
      patterns[40894] = 25'b10011111_10111100_01011011_1;
      patterns[40895] = 25'b10011111_10111101_01011100_1;
      patterns[40896] = 25'b10011111_10111110_01011101_1;
      patterns[40897] = 25'b10011111_10111111_01011110_1;
      patterns[40898] = 25'b10011111_11000000_01011111_1;
      patterns[40899] = 25'b10011111_11000001_01100000_1;
      patterns[40900] = 25'b10011111_11000010_01100001_1;
      patterns[40901] = 25'b10011111_11000011_01100010_1;
      patterns[40902] = 25'b10011111_11000100_01100011_1;
      patterns[40903] = 25'b10011111_11000101_01100100_1;
      patterns[40904] = 25'b10011111_11000110_01100101_1;
      patterns[40905] = 25'b10011111_11000111_01100110_1;
      patterns[40906] = 25'b10011111_11001000_01100111_1;
      patterns[40907] = 25'b10011111_11001001_01101000_1;
      patterns[40908] = 25'b10011111_11001010_01101001_1;
      patterns[40909] = 25'b10011111_11001011_01101010_1;
      patterns[40910] = 25'b10011111_11001100_01101011_1;
      patterns[40911] = 25'b10011111_11001101_01101100_1;
      patterns[40912] = 25'b10011111_11001110_01101101_1;
      patterns[40913] = 25'b10011111_11001111_01101110_1;
      patterns[40914] = 25'b10011111_11010000_01101111_1;
      patterns[40915] = 25'b10011111_11010001_01110000_1;
      patterns[40916] = 25'b10011111_11010010_01110001_1;
      patterns[40917] = 25'b10011111_11010011_01110010_1;
      patterns[40918] = 25'b10011111_11010100_01110011_1;
      patterns[40919] = 25'b10011111_11010101_01110100_1;
      patterns[40920] = 25'b10011111_11010110_01110101_1;
      patterns[40921] = 25'b10011111_11010111_01110110_1;
      patterns[40922] = 25'b10011111_11011000_01110111_1;
      patterns[40923] = 25'b10011111_11011001_01111000_1;
      patterns[40924] = 25'b10011111_11011010_01111001_1;
      patterns[40925] = 25'b10011111_11011011_01111010_1;
      patterns[40926] = 25'b10011111_11011100_01111011_1;
      patterns[40927] = 25'b10011111_11011101_01111100_1;
      patterns[40928] = 25'b10011111_11011110_01111101_1;
      patterns[40929] = 25'b10011111_11011111_01111110_1;
      patterns[40930] = 25'b10011111_11100000_01111111_1;
      patterns[40931] = 25'b10011111_11100001_10000000_1;
      patterns[40932] = 25'b10011111_11100010_10000001_1;
      patterns[40933] = 25'b10011111_11100011_10000010_1;
      patterns[40934] = 25'b10011111_11100100_10000011_1;
      patterns[40935] = 25'b10011111_11100101_10000100_1;
      patterns[40936] = 25'b10011111_11100110_10000101_1;
      patterns[40937] = 25'b10011111_11100111_10000110_1;
      patterns[40938] = 25'b10011111_11101000_10000111_1;
      patterns[40939] = 25'b10011111_11101001_10001000_1;
      patterns[40940] = 25'b10011111_11101010_10001001_1;
      patterns[40941] = 25'b10011111_11101011_10001010_1;
      patterns[40942] = 25'b10011111_11101100_10001011_1;
      patterns[40943] = 25'b10011111_11101101_10001100_1;
      patterns[40944] = 25'b10011111_11101110_10001101_1;
      patterns[40945] = 25'b10011111_11101111_10001110_1;
      patterns[40946] = 25'b10011111_11110000_10001111_1;
      patterns[40947] = 25'b10011111_11110001_10010000_1;
      patterns[40948] = 25'b10011111_11110010_10010001_1;
      patterns[40949] = 25'b10011111_11110011_10010010_1;
      patterns[40950] = 25'b10011111_11110100_10010011_1;
      patterns[40951] = 25'b10011111_11110101_10010100_1;
      patterns[40952] = 25'b10011111_11110110_10010101_1;
      patterns[40953] = 25'b10011111_11110111_10010110_1;
      patterns[40954] = 25'b10011111_11111000_10010111_1;
      patterns[40955] = 25'b10011111_11111001_10011000_1;
      patterns[40956] = 25'b10011111_11111010_10011001_1;
      patterns[40957] = 25'b10011111_11111011_10011010_1;
      patterns[40958] = 25'b10011111_11111100_10011011_1;
      patterns[40959] = 25'b10011111_11111101_10011100_1;
      patterns[40960] = 25'b10011111_11111110_10011101_1;
      patterns[40961] = 25'b10011111_11111111_10011110_1;
      patterns[40962] = 25'b10100000_00000000_10100000_0;
      patterns[40963] = 25'b10100000_00000001_10100001_0;
      patterns[40964] = 25'b10100000_00000010_10100010_0;
      patterns[40965] = 25'b10100000_00000011_10100011_0;
      patterns[40966] = 25'b10100000_00000100_10100100_0;
      patterns[40967] = 25'b10100000_00000101_10100101_0;
      patterns[40968] = 25'b10100000_00000110_10100110_0;
      patterns[40969] = 25'b10100000_00000111_10100111_0;
      patterns[40970] = 25'b10100000_00001000_10101000_0;
      patterns[40971] = 25'b10100000_00001001_10101001_0;
      patterns[40972] = 25'b10100000_00001010_10101010_0;
      patterns[40973] = 25'b10100000_00001011_10101011_0;
      patterns[40974] = 25'b10100000_00001100_10101100_0;
      patterns[40975] = 25'b10100000_00001101_10101101_0;
      patterns[40976] = 25'b10100000_00001110_10101110_0;
      patterns[40977] = 25'b10100000_00001111_10101111_0;
      patterns[40978] = 25'b10100000_00010000_10110000_0;
      patterns[40979] = 25'b10100000_00010001_10110001_0;
      patterns[40980] = 25'b10100000_00010010_10110010_0;
      patterns[40981] = 25'b10100000_00010011_10110011_0;
      patterns[40982] = 25'b10100000_00010100_10110100_0;
      patterns[40983] = 25'b10100000_00010101_10110101_0;
      patterns[40984] = 25'b10100000_00010110_10110110_0;
      patterns[40985] = 25'b10100000_00010111_10110111_0;
      patterns[40986] = 25'b10100000_00011000_10111000_0;
      patterns[40987] = 25'b10100000_00011001_10111001_0;
      patterns[40988] = 25'b10100000_00011010_10111010_0;
      patterns[40989] = 25'b10100000_00011011_10111011_0;
      patterns[40990] = 25'b10100000_00011100_10111100_0;
      patterns[40991] = 25'b10100000_00011101_10111101_0;
      patterns[40992] = 25'b10100000_00011110_10111110_0;
      patterns[40993] = 25'b10100000_00011111_10111111_0;
      patterns[40994] = 25'b10100000_00100000_11000000_0;
      patterns[40995] = 25'b10100000_00100001_11000001_0;
      patterns[40996] = 25'b10100000_00100010_11000010_0;
      patterns[40997] = 25'b10100000_00100011_11000011_0;
      patterns[40998] = 25'b10100000_00100100_11000100_0;
      patterns[40999] = 25'b10100000_00100101_11000101_0;
      patterns[41000] = 25'b10100000_00100110_11000110_0;
      patterns[41001] = 25'b10100000_00100111_11000111_0;
      patterns[41002] = 25'b10100000_00101000_11001000_0;
      patterns[41003] = 25'b10100000_00101001_11001001_0;
      patterns[41004] = 25'b10100000_00101010_11001010_0;
      patterns[41005] = 25'b10100000_00101011_11001011_0;
      patterns[41006] = 25'b10100000_00101100_11001100_0;
      patterns[41007] = 25'b10100000_00101101_11001101_0;
      patterns[41008] = 25'b10100000_00101110_11001110_0;
      patterns[41009] = 25'b10100000_00101111_11001111_0;
      patterns[41010] = 25'b10100000_00110000_11010000_0;
      patterns[41011] = 25'b10100000_00110001_11010001_0;
      patterns[41012] = 25'b10100000_00110010_11010010_0;
      patterns[41013] = 25'b10100000_00110011_11010011_0;
      patterns[41014] = 25'b10100000_00110100_11010100_0;
      patterns[41015] = 25'b10100000_00110101_11010101_0;
      patterns[41016] = 25'b10100000_00110110_11010110_0;
      patterns[41017] = 25'b10100000_00110111_11010111_0;
      patterns[41018] = 25'b10100000_00111000_11011000_0;
      patterns[41019] = 25'b10100000_00111001_11011001_0;
      patterns[41020] = 25'b10100000_00111010_11011010_0;
      patterns[41021] = 25'b10100000_00111011_11011011_0;
      patterns[41022] = 25'b10100000_00111100_11011100_0;
      patterns[41023] = 25'b10100000_00111101_11011101_0;
      patterns[41024] = 25'b10100000_00111110_11011110_0;
      patterns[41025] = 25'b10100000_00111111_11011111_0;
      patterns[41026] = 25'b10100000_01000000_11100000_0;
      patterns[41027] = 25'b10100000_01000001_11100001_0;
      patterns[41028] = 25'b10100000_01000010_11100010_0;
      patterns[41029] = 25'b10100000_01000011_11100011_0;
      patterns[41030] = 25'b10100000_01000100_11100100_0;
      patterns[41031] = 25'b10100000_01000101_11100101_0;
      patterns[41032] = 25'b10100000_01000110_11100110_0;
      patterns[41033] = 25'b10100000_01000111_11100111_0;
      patterns[41034] = 25'b10100000_01001000_11101000_0;
      patterns[41035] = 25'b10100000_01001001_11101001_0;
      patterns[41036] = 25'b10100000_01001010_11101010_0;
      patterns[41037] = 25'b10100000_01001011_11101011_0;
      patterns[41038] = 25'b10100000_01001100_11101100_0;
      patterns[41039] = 25'b10100000_01001101_11101101_0;
      patterns[41040] = 25'b10100000_01001110_11101110_0;
      patterns[41041] = 25'b10100000_01001111_11101111_0;
      patterns[41042] = 25'b10100000_01010000_11110000_0;
      patterns[41043] = 25'b10100000_01010001_11110001_0;
      patterns[41044] = 25'b10100000_01010010_11110010_0;
      patterns[41045] = 25'b10100000_01010011_11110011_0;
      patterns[41046] = 25'b10100000_01010100_11110100_0;
      patterns[41047] = 25'b10100000_01010101_11110101_0;
      patterns[41048] = 25'b10100000_01010110_11110110_0;
      patterns[41049] = 25'b10100000_01010111_11110111_0;
      patterns[41050] = 25'b10100000_01011000_11111000_0;
      patterns[41051] = 25'b10100000_01011001_11111001_0;
      patterns[41052] = 25'b10100000_01011010_11111010_0;
      patterns[41053] = 25'b10100000_01011011_11111011_0;
      patterns[41054] = 25'b10100000_01011100_11111100_0;
      patterns[41055] = 25'b10100000_01011101_11111101_0;
      patterns[41056] = 25'b10100000_01011110_11111110_0;
      patterns[41057] = 25'b10100000_01011111_11111111_0;
      patterns[41058] = 25'b10100000_01100000_00000000_1;
      patterns[41059] = 25'b10100000_01100001_00000001_1;
      patterns[41060] = 25'b10100000_01100010_00000010_1;
      patterns[41061] = 25'b10100000_01100011_00000011_1;
      patterns[41062] = 25'b10100000_01100100_00000100_1;
      patterns[41063] = 25'b10100000_01100101_00000101_1;
      patterns[41064] = 25'b10100000_01100110_00000110_1;
      patterns[41065] = 25'b10100000_01100111_00000111_1;
      patterns[41066] = 25'b10100000_01101000_00001000_1;
      patterns[41067] = 25'b10100000_01101001_00001001_1;
      patterns[41068] = 25'b10100000_01101010_00001010_1;
      patterns[41069] = 25'b10100000_01101011_00001011_1;
      patterns[41070] = 25'b10100000_01101100_00001100_1;
      patterns[41071] = 25'b10100000_01101101_00001101_1;
      patterns[41072] = 25'b10100000_01101110_00001110_1;
      patterns[41073] = 25'b10100000_01101111_00001111_1;
      patterns[41074] = 25'b10100000_01110000_00010000_1;
      patterns[41075] = 25'b10100000_01110001_00010001_1;
      patterns[41076] = 25'b10100000_01110010_00010010_1;
      patterns[41077] = 25'b10100000_01110011_00010011_1;
      patterns[41078] = 25'b10100000_01110100_00010100_1;
      patterns[41079] = 25'b10100000_01110101_00010101_1;
      patterns[41080] = 25'b10100000_01110110_00010110_1;
      patterns[41081] = 25'b10100000_01110111_00010111_1;
      patterns[41082] = 25'b10100000_01111000_00011000_1;
      patterns[41083] = 25'b10100000_01111001_00011001_1;
      patterns[41084] = 25'b10100000_01111010_00011010_1;
      patterns[41085] = 25'b10100000_01111011_00011011_1;
      patterns[41086] = 25'b10100000_01111100_00011100_1;
      patterns[41087] = 25'b10100000_01111101_00011101_1;
      patterns[41088] = 25'b10100000_01111110_00011110_1;
      patterns[41089] = 25'b10100000_01111111_00011111_1;
      patterns[41090] = 25'b10100000_10000000_00100000_1;
      patterns[41091] = 25'b10100000_10000001_00100001_1;
      patterns[41092] = 25'b10100000_10000010_00100010_1;
      patterns[41093] = 25'b10100000_10000011_00100011_1;
      patterns[41094] = 25'b10100000_10000100_00100100_1;
      patterns[41095] = 25'b10100000_10000101_00100101_1;
      patterns[41096] = 25'b10100000_10000110_00100110_1;
      patterns[41097] = 25'b10100000_10000111_00100111_1;
      patterns[41098] = 25'b10100000_10001000_00101000_1;
      patterns[41099] = 25'b10100000_10001001_00101001_1;
      patterns[41100] = 25'b10100000_10001010_00101010_1;
      patterns[41101] = 25'b10100000_10001011_00101011_1;
      patterns[41102] = 25'b10100000_10001100_00101100_1;
      patterns[41103] = 25'b10100000_10001101_00101101_1;
      patterns[41104] = 25'b10100000_10001110_00101110_1;
      patterns[41105] = 25'b10100000_10001111_00101111_1;
      patterns[41106] = 25'b10100000_10010000_00110000_1;
      patterns[41107] = 25'b10100000_10010001_00110001_1;
      patterns[41108] = 25'b10100000_10010010_00110010_1;
      patterns[41109] = 25'b10100000_10010011_00110011_1;
      patterns[41110] = 25'b10100000_10010100_00110100_1;
      patterns[41111] = 25'b10100000_10010101_00110101_1;
      patterns[41112] = 25'b10100000_10010110_00110110_1;
      patterns[41113] = 25'b10100000_10010111_00110111_1;
      patterns[41114] = 25'b10100000_10011000_00111000_1;
      patterns[41115] = 25'b10100000_10011001_00111001_1;
      patterns[41116] = 25'b10100000_10011010_00111010_1;
      patterns[41117] = 25'b10100000_10011011_00111011_1;
      patterns[41118] = 25'b10100000_10011100_00111100_1;
      patterns[41119] = 25'b10100000_10011101_00111101_1;
      patterns[41120] = 25'b10100000_10011110_00111110_1;
      patterns[41121] = 25'b10100000_10011111_00111111_1;
      patterns[41122] = 25'b10100000_10100000_01000000_1;
      patterns[41123] = 25'b10100000_10100001_01000001_1;
      patterns[41124] = 25'b10100000_10100010_01000010_1;
      patterns[41125] = 25'b10100000_10100011_01000011_1;
      patterns[41126] = 25'b10100000_10100100_01000100_1;
      patterns[41127] = 25'b10100000_10100101_01000101_1;
      patterns[41128] = 25'b10100000_10100110_01000110_1;
      patterns[41129] = 25'b10100000_10100111_01000111_1;
      patterns[41130] = 25'b10100000_10101000_01001000_1;
      patterns[41131] = 25'b10100000_10101001_01001001_1;
      patterns[41132] = 25'b10100000_10101010_01001010_1;
      patterns[41133] = 25'b10100000_10101011_01001011_1;
      patterns[41134] = 25'b10100000_10101100_01001100_1;
      patterns[41135] = 25'b10100000_10101101_01001101_1;
      patterns[41136] = 25'b10100000_10101110_01001110_1;
      patterns[41137] = 25'b10100000_10101111_01001111_1;
      patterns[41138] = 25'b10100000_10110000_01010000_1;
      patterns[41139] = 25'b10100000_10110001_01010001_1;
      patterns[41140] = 25'b10100000_10110010_01010010_1;
      patterns[41141] = 25'b10100000_10110011_01010011_1;
      patterns[41142] = 25'b10100000_10110100_01010100_1;
      patterns[41143] = 25'b10100000_10110101_01010101_1;
      patterns[41144] = 25'b10100000_10110110_01010110_1;
      patterns[41145] = 25'b10100000_10110111_01010111_1;
      patterns[41146] = 25'b10100000_10111000_01011000_1;
      patterns[41147] = 25'b10100000_10111001_01011001_1;
      patterns[41148] = 25'b10100000_10111010_01011010_1;
      patterns[41149] = 25'b10100000_10111011_01011011_1;
      patterns[41150] = 25'b10100000_10111100_01011100_1;
      patterns[41151] = 25'b10100000_10111101_01011101_1;
      patterns[41152] = 25'b10100000_10111110_01011110_1;
      patterns[41153] = 25'b10100000_10111111_01011111_1;
      patterns[41154] = 25'b10100000_11000000_01100000_1;
      patterns[41155] = 25'b10100000_11000001_01100001_1;
      patterns[41156] = 25'b10100000_11000010_01100010_1;
      patterns[41157] = 25'b10100000_11000011_01100011_1;
      patterns[41158] = 25'b10100000_11000100_01100100_1;
      patterns[41159] = 25'b10100000_11000101_01100101_1;
      patterns[41160] = 25'b10100000_11000110_01100110_1;
      patterns[41161] = 25'b10100000_11000111_01100111_1;
      patterns[41162] = 25'b10100000_11001000_01101000_1;
      patterns[41163] = 25'b10100000_11001001_01101001_1;
      patterns[41164] = 25'b10100000_11001010_01101010_1;
      patterns[41165] = 25'b10100000_11001011_01101011_1;
      patterns[41166] = 25'b10100000_11001100_01101100_1;
      patterns[41167] = 25'b10100000_11001101_01101101_1;
      patterns[41168] = 25'b10100000_11001110_01101110_1;
      patterns[41169] = 25'b10100000_11001111_01101111_1;
      patterns[41170] = 25'b10100000_11010000_01110000_1;
      patterns[41171] = 25'b10100000_11010001_01110001_1;
      patterns[41172] = 25'b10100000_11010010_01110010_1;
      patterns[41173] = 25'b10100000_11010011_01110011_1;
      patterns[41174] = 25'b10100000_11010100_01110100_1;
      patterns[41175] = 25'b10100000_11010101_01110101_1;
      patterns[41176] = 25'b10100000_11010110_01110110_1;
      patterns[41177] = 25'b10100000_11010111_01110111_1;
      patterns[41178] = 25'b10100000_11011000_01111000_1;
      patterns[41179] = 25'b10100000_11011001_01111001_1;
      patterns[41180] = 25'b10100000_11011010_01111010_1;
      patterns[41181] = 25'b10100000_11011011_01111011_1;
      patterns[41182] = 25'b10100000_11011100_01111100_1;
      patterns[41183] = 25'b10100000_11011101_01111101_1;
      patterns[41184] = 25'b10100000_11011110_01111110_1;
      patterns[41185] = 25'b10100000_11011111_01111111_1;
      patterns[41186] = 25'b10100000_11100000_10000000_1;
      patterns[41187] = 25'b10100000_11100001_10000001_1;
      patterns[41188] = 25'b10100000_11100010_10000010_1;
      patterns[41189] = 25'b10100000_11100011_10000011_1;
      patterns[41190] = 25'b10100000_11100100_10000100_1;
      patterns[41191] = 25'b10100000_11100101_10000101_1;
      patterns[41192] = 25'b10100000_11100110_10000110_1;
      patterns[41193] = 25'b10100000_11100111_10000111_1;
      patterns[41194] = 25'b10100000_11101000_10001000_1;
      patterns[41195] = 25'b10100000_11101001_10001001_1;
      patterns[41196] = 25'b10100000_11101010_10001010_1;
      patterns[41197] = 25'b10100000_11101011_10001011_1;
      patterns[41198] = 25'b10100000_11101100_10001100_1;
      patterns[41199] = 25'b10100000_11101101_10001101_1;
      patterns[41200] = 25'b10100000_11101110_10001110_1;
      patterns[41201] = 25'b10100000_11101111_10001111_1;
      patterns[41202] = 25'b10100000_11110000_10010000_1;
      patterns[41203] = 25'b10100000_11110001_10010001_1;
      patterns[41204] = 25'b10100000_11110010_10010010_1;
      patterns[41205] = 25'b10100000_11110011_10010011_1;
      patterns[41206] = 25'b10100000_11110100_10010100_1;
      patterns[41207] = 25'b10100000_11110101_10010101_1;
      patterns[41208] = 25'b10100000_11110110_10010110_1;
      patterns[41209] = 25'b10100000_11110111_10010111_1;
      patterns[41210] = 25'b10100000_11111000_10011000_1;
      patterns[41211] = 25'b10100000_11111001_10011001_1;
      patterns[41212] = 25'b10100000_11111010_10011010_1;
      patterns[41213] = 25'b10100000_11111011_10011011_1;
      patterns[41214] = 25'b10100000_11111100_10011100_1;
      patterns[41215] = 25'b10100000_11111101_10011101_1;
      patterns[41216] = 25'b10100000_11111110_10011110_1;
      patterns[41217] = 25'b10100000_11111111_10011111_1;
      patterns[41218] = 25'b10100001_00000000_10100001_0;
      patterns[41219] = 25'b10100001_00000001_10100010_0;
      patterns[41220] = 25'b10100001_00000010_10100011_0;
      patterns[41221] = 25'b10100001_00000011_10100100_0;
      patterns[41222] = 25'b10100001_00000100_10100101_0;
      patterns[41223] = 25'b10100001_00000101_10100110_0;
      patterns[41224] = 25'b10100001_00000110_10100111_0;
      patterns[41225] = 25'b10100001_00000111_10101000_0;
      patterns[41226] = 25'b10100001_00001000_10101001_0;
      patterns[41227] = 25'b10100001_00001001_10101010_0;
      patterns[41228] = 25'b10100001_00001010_10101011_0;
      patterns[41229] = 25'b10100001_00001011_10101100_0;
      patterns[41230] = 25'b10100001_00001100_10101101_0;
      patterns[41231] = 25'b10100001_00001101_10101110_0;
      patterns[41232] = 25'b10100001_00001110_10101111_0;
      patterns[41233] = 25'b10100001_00001111_10110000_0;
      patterns[41234] = 25'b10100001_00010000_10110001_0;
      patterns[41235] = 25'b10100001_00010001_10110010_0;
      patterns[41236] = 25'b10100001_00010010_10110011_0;
      patterns[41237] = 25'b10100001_00010011_10110100_0;
      patterns[41238] = 25'b10100001_00010100_10110101_0;
      patterns[41239] = 25'b10100001_00010101_10110110_0;
      patterns[41240] = 25'b10100001_00010110_10110111_0;
      patterns[41241] = 25'b10100001_00010111_10111000_0;
      patterns[41242] = 25'b10100001_00011000_10111001_0;
      patterns[41243] = 25'b10100001_00011001_10111010_0;
      patterns[41244] = 25'b10100001_00011010_10111011_0;
      patterns[41245] = 25'b10100001_00011011_10111100_0;
      patterns[41246] = 25'b10100001_00011100_10111101_0;
      patterns[41247] = 25'b10100001_00011101_10111110_0;
      patterns[41248] = 25'b10100001_00011110_10111111_0;
      patterns[41249] = 25'b10100001_00011111_11000000_0;
      patterns[41250] = 25'b10100001_00100000_11000001_0;
      patterns[41251] = 25'b10100001_00100001_11000010_0;
      patterns[41252] = 25'b10100001_00100010_11000011_0;
      patterns[41253] = 25'b10100001_00100011_11000100_0;
      patterns[41254] = 25'b10100001_00100100_11000101_0;
      patterns[41255] = 25'b10100001_00100101_11000110_0;
      patterns[41256] = 25'b10100001_00100110_11000111_0;
      patterns[41257] = 25'b10100001_00100111_11001000_0;
      patterns[41258] = 25'b10100001_00101000_11001001_0;
      patterns[41259] = 25'b10100001_00101001_11001010_0;
      patterns[41260] = 25'b10100001_00101010_11001011_0;
      patterns[41261] = 25'b10100001_00101011_11001100_0;
      patterns[41262] = 25'b10100001_00101100_11001101_0;
      patterns[41263] = 25'b10100001_00101101_11001110_0;
      patterns[41264] = 25'b10100001_00101110_11001111_0;
      patterns[41265] = 25'b10100001_00101111_11010000_0;
      patterns[41266] = 25'b10100001_00110000_11010001_0;
      patterns[41267] = 25'b10100001_00110001_11010010_0;
      patterns[41268] = 25'b10100001_00110010_11010011_0;
      patterns[41269] = 25'b10100001_00110011_11010100_0;
      patterns[41270] = 25'b10100001_00110100_11010101_0;
      patterns[41271] = 25'b10100001_00110101_11010110_0;
      patterns[41272] = 25'b10100001_00110110_11010111_0;
      patterns[41273] = 25'b10100001_00110111_11011000_0;
      patterns[41274] = 25'b10100001_00111000_11011001_0;
      patterns[41275] = 25'b10100001_00111001_11011010_0;
      patterns[41276] = 25'b10100001_00111010_11011011_0;
      patterns[41277] = 25'b10100001_00111011_11011100_0;
      patterns[41278] = 25'b10100001_00111100_11011101_0;
      patterns[41279] = 25'b10100001_00111101_11011110_0;
      patterns[41280] = 25'b10100001_00111110_11011111_0;
      patterns[41281] = 25'b10100001_00111111_11100000_0;
      patterns[41282] = 25'b10100001_01000000_11100001_0;
      patterns[41283] = 25'b10100001_01000001_11100010_0;
      patterns[41284] = 25'b10100001_01000010_11100011_0;
      patterns[41285] = 25'b10100001_01000011_11100100_0;
      patterns[41286] = 25'b10100001_01000100_11100101_0;
      patterns[41287] = 25'b10100001_01000101_11100110_0;
      patterns[41288] = 25'b10100001_01000110_11100111_0;
      patterns[41289] = 25'b10100001_01000111_11101000_0;
      patterns[41290] = 25'b10100001_01001000_11101001_0;
      patterns[41291] = 25'b10100001_01001001_11101010_0;
      patterns[41292] = 25'b10100001_01001010_11101011_0;
      patterns[41293] = 25'b10100001_01001011_11101100_0;
      patterns[41294] = 25'b10100001_01001100_11101101_0;
      patterns[41295] = 25'b10100001_01001101_11101110_0;
      patterns[41296] = 25'b10100001_01001110_11101111_0;
      patterns[41297] = 25'b10100001_01001111_11110000_0;
      patterns[41298] = 25'b10100001_01010000_11110001_0;
      patterns[41299] = 25'b10100001_01010001_11110010_0;
      patterns[41300] = 25'b10100001_01010010_11110011_0;
      patterns[41301] = 25'b10100001_01010011_11110100_0;
      patterns[41302] = 25'b10100001_01010100_11110101_0;
      patterns[41303] = 25'b10100001_01010101_11110110_0;
      patterns[41304] = 25'b10100001_01010110_11110111_0;
      patterns[41305] = 25'b10100001_01010111_11111000_0;
      patterns[41306] = 25'b10100001_01011000_11111001_0;
      patterns[41307] = 25'b10100001_01011001_11111010_0;
      patterns[41308] = 25'b10100001_01011010_11111011_0;
      patterns[41309] = 25'b10100001_01011011_11111100_0;
      patterns[41310] = 25'b10100001_01011100_11111101_0;
      patterns[41311] = 25'b10100001_01011101_11111110_0;
      patterns[41312] = 25'b10100001_01011110_11111111_0;
      patterns[41313] = 25'b10100001_01011111_00000000_1;
      patterns[41314] = 25'b10100001_01100000_00000001_1;
      patterns[41315] = 25'b10100001_01100001_00000010_1;
      patterns[41316] = 25'b10100001_01100010_00000011_1;
      patterns[41317] = 25'b10100001_01100011_00000100_1;
      patterns[41318] = 25'b10100001_01100100_00000101_1;
      patterns[41319] = 25'b10100001_01100101_00000110_1;
      patterns[41320] = 25'b10100001_01100110_00000111_1;
      patterns[41321] = 25'b10100001_01100111_00001000_1;
      patterns[41322] = 25'b10100001_01101000_00001001_1;
      patterns[41323] = 25'b10100001_01101001_00001010_1;
      patterns[41324] = 25'b10100001_01101010_00001011_1;
      patterns[41325] = 25'b10100001_01101011_00001100_1;
      patterns[41326] = 25'b10100001_01101100_00001101_1;
      patterns[41327] = 25'b10100001_01101101_00001110_1;
      patterns[41328] = 25'b10100001_01101110_00001111_1;
      patterns[41329] = 25'b10100001_01101111_00010000_1;
      patterns[41330] = 25'b10100001_01110000_00010001_1;
      patterns[41331] = 25'b10100001_01110001_00010010_1;
      patterns[41332] = 25'b10100001_01110010_00010011_1;
      patterns[41333] = 25'b10100001_01110011_00010100_1;
      patterns[41334] = 25'b10100001_01110100_00010101_1;
      patterns[41335] = 25'b10100001_01110101_00010110_1;
      patterns[41336] = 25'b10100001_01110110_00010111_1;
      patterns[41337] = 25'b10100001_01110111_00011000_1;
      patterns[41338] = 25'b10100001_01111000_00011001_1;
      patterns[41339] = 25'b10100001_01111001_00011010_1;
      patterns[41340] = 25'b10100001_01111010_00011011_1;
      patterns[41341] = 25'b10100001_01111011_00011100_1;
      patterns[41342] = 25'b10100001_01111100_00011101_1;
      patterns[41343] = 25'b10100001_01111101_00011110_1;
      patterns[41344] = 25'b10100001_01111110_00011111_1;
      patterns[41345] = 25'b10100001_01111111_00100000_1;
      patterns[41346] = 25'b10100001_10000000_00100001_1;
      patterns[41347] = 25'b10100001_10000001_00100010_1;
      patterns[41348] = 25'b10100001_10000010_00100011_1;
      patterns[41349] = 25'b10100001_10000011_00100100_1;
      patterns[41350] = 25'b10100001_10000100_00100101_1;
      patterns[41351] = 25'b10100001_10000101_00100110_1;
      patterns[41352] = 25'b10100001_10000110_00100111_1;
      patterns[41353] = 25'b10100001_10000111_00101000_1;
      patterns[41354] = 25'b10100001_10001000_00101001_1;
      patterns[41355] = 25'b10100001_10001001_00101010_1;
      patterns[41356] = 25'b10100001_10001010_00101011_1;
      patterns[41357] = 25'b10100001_10001011_00101100_1;
      patterns[41358] = 25'b10100001_10001100_00101101_1;
      patterns[41359] = 25'b10100001_10001101_00101110_1;
      patterns[41360] = 25'b10100001_10001110_00101111_1;
      patterns[41361] = 25'b10100001_10001111_00110000_1;
      patterns[41362] = 25'b10100001_10010000_00110001_1;
      patterns[41363] = 25'b10100001_10010001_00110010_1;
      patterns[41364] = 25'b10100001_10010010_00110011_1;
      patterns[41365] = 25'b10100001_10010011_00110100_1;
      patterns[41366] = 25'b10100001_10010100_00110101_1;
      patterns[41367] = 25'b10100001_10010101_00110110_1;
      patterns[41368] = 25'b10100001_10010110_00110111_1;
      patterns[41369] = 25'b10100001_10010111_00111000_1;
      patterns[41370] = 25'b10100001_10011000_00111001_1;
      patterns[41371] = 25'b10100001_10011001_00111010_1;
      patterns[41372] = 25'b10100001_10011010_00111011_1;
      patterns[41373] = 25'b10100001_10011011_00111100_1;
      patterns[41374] = 25'b10100001_10011100_00111101_1;
      patterns[41375] = 25'b10100001_10011101_00111110_1;
      patterns[41376] = 25'b10100001_10011110_00111111_1;
      patterns[41377] = 25'b10100001_10011111_01000000_1;
      patterns[41378] = 25'b10100001_10100000_01000001_1;
      patterns[41379] = 25'b10100001_10100001_01000010_1;
      patterns[41380] = 25'b10100001_10100010_01000011_1;
      patterns[41381] = 25'b10100001_10100011_01000100_1;
      patterns[41382] = 25'b10100001_10100100_01000101_1;
      patterns[41383] = 25'b10100001_10100101_01000110_1;
      patterns[41384] = 25'b10100001_10100110_01000111_1;
      patterns[41385] = 25'b10100001_10100111_01001000_1;
      patterns[41386] = 25'b10100001_10101000_01001001_1;
      patterns[41387] = 25'b10100001_10101001_01001010_1;
      patterns[41388] = 25'b10100001_10101010_01001011_1;
      patterns[41389] = 25'b10100001_10101011_01001100_1;
      patterns[41390] = 25'b10100001_10101100_01001101_1;
      patterns[41391] = 25'b10100001_10101101_01001110_1;
      patterns[41392] = 25'b10100001_10101110_01001111_1;
      patterns[41393] = 25'b10100001_10101111_01010000_1;
      patterns[41394] = 25'b10100001_10110000_01010001_1;
      patterns[41395] = 25'b10100001_10110001_01010010_1;
      patterns[41396] = 25'b10100001_10110010_01010011_1;
      patterns[41397] = 25'b10100001_10110011_01010100_1;
      patterns[41398] = 25'b10100001_10110100_01010101_1;
      patterns[41399] = 25'b10100001_10110101_01010110_1;
      patterns[41400] = 25'b10100001_10110110_01010111_1;
      patterns[41401] = 25'b10100001_10110111_01011000_1;
      patterns[41402] = 25'b10100001_10111000_01011001_1;
      patterns[41403] = 25'b10100001_10111001_01011010_1;
      patterns[41404] = 25'b10100001_10111010_01011011_1;
      patterns[41405] = 25'b10100001_10111011_01011100_1;
      patterns[41406] = 25'b10100001_10111100_01011101_1;
      patterns[41407] = 25'b10100001_10111101_01011110_1;
      patterns[41408] = 25'b10100001_10111110_01011111_1;
      patterns[41409] = 25'b10100001_10111111_01100000_1;
      patterns[41410] = 25'b10100001_11000000_01100001_1;
      patterns[41411] = 25'b10100001_11000001_01100010_1;
      patterns[41412] = 25'b10100001_11000010_01100011_1;
      patterns[41413] = 25'b10100001_11000011_01100100_1;
      patterns[41414] = 25'b10100001_11000100_01100101_1;
      patterns[41415] = 25'b10100001_11000101_01100110_1;
      patterns[41416] = 25'b10100001_11000110_01100111_1;
      patterns[41417] = 25'b10100001_11000111_01101000_1;
      patterns[41418] = 25'b10100001_11001000_01101001_1;
      patterns[41419] = 25'b10100001_11001001_01101010_1;
      patterns[41420] = 25'b10100001_11001010_01101011_1;
      patterns[41421] = 25'b10100001_11001011_01101100_1;
      patterns[41422] = 25'b10100001_11001100_01101101_1;
      patterns[41423] = 25'b10100001_11001101_01101110_1;
      patterns[41424] = 25'b10100001_11001110_01101111_1;
      patterns[41425] = 25'b10100001_11001111_01110000_1;
      patterns[41426] = 25'b10100001_11010000_01110001_1;
      patterns[41427] = 25'b10100001_11010001_01110010_1;
      patterns[41428] = 25'b10100001_11010010_01110011_1;
      patterns[41429] = 25'b10100001_11010011_01110100_1;
      patterns[41430] = 25'b10100001_11010100_01110101_1;
      patterns[41431] = 25'b10100001_11010101_01110110_1;
      patterns[41432] = 25'b10100001_11010110_01110111_1;
      patterns[41433] = 25'b10100001_11010111_01111000_1;
      patterns[41434] = 25'b10100001_11011000_01111001_1;
      patterns[41435] = 25'b10100001_11011001_01111010_1;
      patterns[41436] = 25'b10100001_11011010_01111011_1;
      patterns[41437] = 25'b10100001_11011011_01111100_1;
      patterns[41438] = 25'b10100001_11011100_01111101_1;
      patterns[41439] = 25'b10100001_11011101_01111110_1;
      patterns[41440] = 25'b10100001_11011110_01111111_1;
      patterns[41441] = 25'b10100001_11011111_10000000_1;
      patterns[41442] = 25'b10100001_11100000_10000001_1;
      patterns[41443] = 25'b10100001_11100001_10000010_1;
      patterns[41444] = 25'b10100001_11100010_10000011_1;
      patterns[41445] = 25'b10100001_11100011_10000100_1;
      patterns[41446] = 25'b10100001_11100100_10000101_1;
      patterns[41447] = 25'b10100001_11100101_10000110_1;
      patterns[41448] = 25'b10100001_11100110_10000111_1;
      patterns[41449] = 25'b10100001_11100111_10001000_1;
      patterns[41450] = 25'b10100001_11101000_10001001_1;
      patterns[41451] = 25'b10100001_11101001_10001010_1;
      patterns[41452] = 25'b10100001_11101010_10001011_1;
      patterns[41453] = 25'b10100001_11101011_10001100_1;
      patterns[41454] = 25'b10100001_11101100_10001101_1;
      patterns[41455] = 25'b10100001_11101101_10001110_1;
      patterns[41456] = 25'b10100001_11101110_10001111_1;
      patterns[41457] = 25'b10100001_11101111_10010000_1;
      patterns[41458] = 25'b10100001_11110000_10010001_1;
      patterns[41459] = 25'b10100001_11110001_10010010_1;
      patterns[41460] = 25'b10100001_11110010_10010011_1;
      patterns[41461] = 25'b10100001_11110011_10010100_1;
      patterns[41462] = 25'b10100001_11110100_10010101_1;
      patterns[41463] = 25'b10100001_11110101_10010110_1;
      patterns[41464] = 25'b10100001_11110110_10010111_1;
      patterns[41465] = 25'b10100001_11110111_10011000_1;
      patterns[41466] = 25'b10100001_11111000_10011001_1;
      patterns[41467] = 25'b10100001_11111001_10011010_1;
      patterns[41468] = 25'b10100001_11111010_10011011_1;
      patterns[41469] = 25'b10100001_11111011_10011100_1;
      patterns[41470] = 25'b10100001_11111100_10011101_1;
      patterns[41471] = 25'b10100001_11111101_10011110_1;
      patterns[41472] = 25'b10100001_11111110_10011111_1;
      patterns[41473] = 25'b10100001_11111111_10100000_1;
      patterns[41474] = 25'b10100010_00000000_10100010_0;
      patterns[41475] = 25'b10100010_00000001_10100011_0;
      patterns[41476] = 25'b10100010_00000010_10100100_0;
      patterns[41477] = 25'b10100010_00000011_10100101_0;
      patterns[41478] = 25'b10100010_00000100_10100110_0;
      patterns[41479] = 25'b10100010_00000101_10100111_0;
      patterns[41480] = 25'b10100010_00000110_10101000_0;
      patterns[41481] = 25'b10100010_00000111_10101001_0;
      patterns[41482] = 25'b10100010_00001000_10101010_0;
      patterns[41483] = 25'b10100010_00001001_10101011_0;
      patterns[41484] = 25'b10100010_00001010_10101100_0;
      patterns[41485] = 25'b10100010_00001011_10101101_0;
      patterns[41486] = 25'b10100010_00001100_10101110_0;
      patterns[41487] = 25'b10100010_00001101_10101111_0;
      patterns[41488] = 25'b10100010_00001110_10110000_0;
      patterns[41489] = 25'b10100010_00001111_10110001_0;
      patterns[41490] = 25'b10100010_00010000_10110010_0;
      patterns[41491] = 25'b10100010_00010001_10110011_0;
      patterns[41492] = 25'b10100010_00010010_10110100_0;
      patterns[41493] = 25'b10100010_00010011_10110101_0;
      patterns[41494] = 25'b10100010_00010100_10110110_0;
      patterns[41495] = 25'b10100010_00010101_10110111_0;
      patterns[41496] = 25'b10100010_00010110_10111000_0;
      patterns[41497] = 25'b10100010_00010111_10111001_0;
      patterns[41498] = 25'b10100010_00011000_10111010_0;
      patterns[41499] = 25'b10100010_00011001_10111011_0;
      patterns[41500] = 25'b10100010_00011010_10111100_0;
      patterns[41501] = 25'b10100010_00011011_10111101_0;
      patterns[41502] = 25'b10100010_00011100_10111110_0;
      patterns[41503] = 25'b10100010_00011101_10111111_0;
      patterns[41504] = 25'b10100010_00011110_11000000_0;
      patterns[41505] = 25'b10100010_00011111_11000001_0;
      patterns[41506] = 25'b10100010_00100000_11000010_0;
      patterns[41507] = 25'b10100010_00100001_11000011_0;
      patterns[41508] = 25'b10100010_00100010_11000100_0;
      patterns[41509] = 25'b10100010_00100011_11000101_0;
      patterns[41510] = 25'b10100010_00100100_11000110_0;
      patterns[41511] = 25'b10100010_00100101_11000111_0;
      patterns[41512] = 25'b10100010_00100110_11001000_0;
      patterns[41513] = 25'b10100010_00100111_11001001_0;
      patterns[41514] = 25'b10100010_00101000_11001010_0;
      patterns[41515] = 25'b10100010_00101001_11001011_0;
      patterns[41516] = 25'b10100010_00101010_11001100_0;
      patterns[41517] = 25'b10100010_00101011_11001101_0;
      patterns[41518] = 25'b10100010_00101100_11001110_0;
      patterns[41519] = 25'b10100010_00101101_11001111_0;
      patterns[41520] = 25'b10100010_00101110_11010000_0;
      patterns[41521] = 25'b10100010_00101111_11010001_0;
      patterns[41522] = 25'b10100010_00110000_11010010_0;
      patterns[41523] = 25'b10100010_00110001_11010011_0;
      patterns[41524] = 25'b10100010_00110010_11010100_0;
      patterns[41525] = 25'b10100010_00110011_11010101_0;
      patterns[41526] = 25'b10100010_00110100_11010110_0;
      patterns[41527] = 25'b10100010_00110101_11010111_0;
      patterns[41528] = 25'b10100010_00110110_11011000_0;
      patterns[41529] = 25'b10100010_00110111_11011001_0;
      patterns[41530] = 25'b10100010_00111000_11011010_0;
      patterns[41531] = 25'b10100010_00111001_11011011_0;
      patterns[41532] = 25'b10100010_00111010_11011100_0;
      patterns[41533] = 25'b10100010_00111011_11011101_0;
      patterns[41534] = 25'b10100010_00111100_11011110_0;
      patterns[41535] = 25'b10100010_00111101_11011111_0;
      patterns[41536] = 25'b10100010_00111110_11100000_0;
      patterns[41537] = 25'b10100010_00111111_11100001_0;
      patterns[41538] = 25'b10100010_01000000_11100010_0;
      patterns[41539] = 25'b10100010_01000001_11100011_0;
      patterns[41540] = 25'b10100010_01000010_11100100_0;
      patterns[41541] = 25'b10100010_01000011_11100101_0;
      patterns[41542] = 25'b10100010_01000100_11100110_0;
      patterns[41543] = 25'b10100010_01000101_11100111_0;
      patterns[41544] = 25'b10100010_01000110_11101000_0;
      patterns[41545] = 25'b10100010_01000111_11101001_0;
      patterns[41546] = 25'b10100010_01001000_11101010_0;
      patterns[41547] = 25'b10100010_01001001_11101011_0;
      patterns[41548] = 25'b10100010_01001010_11101100_0;
      patterns[41549] = 25'b10100010_01001011_11101101_0;
      patterns[41550] = 25'b10100010_01001100_11101110_0;
      patterns[41551] = 25'b10100010_01001101_11101111_0;
      patterns[41552] = 25'b10100010_01001110_11110000_0;
      patterns[41553] = 25'b10100010_01001111_11110001_0;
      patterns[41554] = 25'b10100010_01010000_11110010_0;
      patterns[41555] = 25'b10100010_01010001_11110011_0;
      patterns[41556] = 25'b10100010_01010010_11110100_0;
      patterns[41557] = 25'b10100010_01010011_11110101_0;
      patterns[41558] = 25'b10100010_01010100_11110110_0;
      patterns[41559] = 25'b10100010_01010101_11110111_0;
      patterns[41560] = 25'b10100010_01010110_11111000_0;
      patterns[41561] = 25'b10100010_01010111_11111001_0;
      patterns[41562] = 25'b10100010_01011000_11111010_0;
      patterns[41563] = 25'b10100010_01011001_11111011_0;
      patterns[41564] = 25'b10100010_01011010_11111100_0;
      patterns[41565] = 25'b10100010_01011011_11111101_0;
      patterns[41566] = 25'b10100010_01011100_11111110_0;
      patterns[41567] = 25'b10100010_01011101_11111111_0;
      patterns[41568] = 25'b10100010_01011110_00000000_1;
      patterns[41569] = 25'b10100010_01011111_00000001_1;
      patterns[41570] = 25'b10100010_01100000_00000010_1;
      patterns[41571] = 25'b10100010_01100001_00000011_1;
      patterns[41572] = 25'b10100010_01100010_00000100_1;
      patterns[41573] = 25'b10100010_01100011_00000101_1;
      patterns[41574] = 25'b10100010_01100100_00000110_1;
      patterns[41575] = 25'b10100010_01100101_00000111_1;
      patterns[41576] = 25'b10100010_01100110_00001000_1;
      patterns[41577] = 25'b10100010_01100111_00001001_1;
      patterns[41578] = 25'b10100010_01101000_00001010_1;
      patterns[41579] = 25'b10100010_01101001_00001011_1;
      patterns[41580] = 25'b10100010_01101010_00001100_1;
      patterns[41581] = 25'b10100010_01101011_00001101_1;
      patterns[41582] = 25'b10100010_01101100_00001110_1;
      patterns[41583] = 25'b10100010_01101101_00001111_1;
      patterns[41584] = 25'b10100010_01101110_00010000_1;
      patterns[41585] = 25'b10100010_01101111_00010001_1;
      patterns[41586] = 25'b10100010_01110000_00010010_1;
      patterns[41587] = 25'b10100010_01110001_00010011_1;
      patterns[41588] = 25'b10100010_01110010_00010100_1;
      patterns[41589] = 25'b10100010_01110011_00010101_1;
      patterns[41590] = 25'b10100010_01110100_00010110_1;
      patterns[41591] = 25'b10100010_01110101_00010111_1;
      patterns[41592] = 25'b10100010_01110110_00011000_1;
      patterns[41593] = 25'b10100010_01110111_00011001_1;
      patterns[41594] = 25'b10100010_01111000_00011010_1;
      patterns[41595] = 25'b10100010_01111001_00011011_1;
      patterns[41596] = 25'b10100010_01111010_00011100_1;
      patterns[41597] = 25'b10100010_01111011_00011101_1;
      patterns[41598] = 25'b10100010_01111100_00011110_1;
      patterns[41599] = 25'b10100010_01111101_00011111_1;
      patterns[41600] = 25'b10100010_01111110_00100000_1;
      patterns[41601] = 25'b10100010_01111111_00100001_1;
      patterns[41602] = 25'b10100010_10000000_00100010_1;
      patterns[41603] = 25'b10100010_10000001_00100011_1;
      patterns[41604] = 25'b10100010_10000010_00100100_1;
      patterns[41605] = 25'b10100010_10000011_00100101_1;
      patterns[41606] = 25'b10100010_10000100_00100110_1;
      patterns[41607] = 25'b10100010_10000101_00100111_1;
      patterns[41608] = 25'b10100010_10000110_00101000_1;
      patterns[41609] = 25'b10100010_10000111_00101001_1;
      patterns[41610] = 25'b10100010_10001000_00101010_1;
      patterns[41611] = 25'b10100010_10001001_00101011_1;
      patterns[41612] = 25'b10100010_10001010_00101100_1;
      patterns[41613] = 25'b10100010_10001011_00101101_1;
      patterns[41614] = 25'b10100010_10001100_00101110_1;
      patterns[41615] = 25'b10100010_10001101_00101111_1;
      patterns[41616] = 25'b10100010_10001110_00110000_1;
      patterns[41617] = 25'b10100010_10001111_00110001_1;
      patterns[41618] = 25'b10100010_10010000_00110010_1;
      patterns[41619] = 25'b10100010_10010001_00110011_1;
      patterns[41620] = 25'b10100010_10010010_00110100_1;
      patterns[41621] = 25'b10100010_10010011_00110101_1;
      patterns[41622] = 25'b10100010_10010100_00110110_1;
      patterns[41623] = 25'b10100010_10010101_00110111_1;
      patterns[41624] = 25'b10100010_10010110_00111000_1;
      patterns[41625] = 25'b10100010_10010111_00111001_1;
      patterns[41626] = 25'b10100010_10011000_00111010_1;
      patterns[41627] = 25'b10100010_10011001_00111011_1;
      patterns[41628] = 25'b10100010_10011010_00111100_1;
      patterns[41629] = 25'b10100010_10011011_00111101_1;
      patterns[41630] = 25'b10100010_10011100_00111110_1;
      patterns[41631] = 25'b10100010_10011101_00111111_1;
      patterns[41632] = 25'b10100010_10011110_01000000_1;
      patterns[41633] = 25'b10100010_10011111_01000001_1;
      patterns[41634] = 25'b10100010_10100000_01000010_1;
      patterns[41635] = 25'b10100010_10100001_01000011_1;
      patterns[41636] = 25'b10100010_10100010_01000100_1;
      patterns[41637] = 25'b10100010_10100011_01000101_1;
      patterns[41638] = 25'b10100010_10100100_01000110_1;
      patterns[41639] = 25'b10100010_10100101_01000111_1;
      patterns[41640] = 25'b10100010_10100110_01001000_1;
      patterns[41641] = 25'b10100010_10100111_01001001_1;
      patterns[41642] = 25'b10100010_10101000_01001010_1;
      patterns[41643] = 25'b10100010_10101001_01001011_1;
      patterns[41644] = 25'b10100010_10101010_01001100_1;
      patterns[41645] = 25'b10100010_10101011_01001101_1;
      patterns[41646] = 25'b10100010_10101100_01001110_1;
      patterns[41647] = 25'b10100010_10101101_01001111_1;
      patterns[41648] = 25'b10100010_10101110_01010000_1;
      patterns[41649] = 25'b10100010_10101111_01010001_1;
      patterns[41650] = 25'b10100010_10110000_01010010_1;
      patterns[41651] = 25'b10100010_10110001_01010011_1;
      patterns[41652] = 25'b10100010_10110010_01010100_1;
      patterns[41653] = 25'b10100010_10110011_01010101_1;
      patterns[41654] = 25'b10100010_10110100_01010110_1;
      patterns[41655] = 25'b10100010_10110101_01010111_1;
      patterns[41656] = 25'b10100010_10110110_01011000_1;
      patterns[41657] = 25'b10100010_10110111_01011001_1;
      patterns[41658] = 25'b10100010_10111000_01011010_1;
      patterns[41659] = 25'b10100010_10111001_01011011_1;
      patterns[41660] = 25'b10100010_10111010_01011100_1;
      patterns[41661] = 25'b10100010_10111011_01011101_1;
      patterns[41662] = 25'b10100010_10111100_01011110_1;
      patterns[41663] = 25'b10100010_10111101_01011111_1;
      patterns[41664] = 25'b10100010_10111110_01100000_1;
      patterns[41665] = 25'b10100010_10111111_01100001_1;
      patterns[41666] = 25'b10100010_11000000_01100010_1;
      patterns[41667] = 25'b10100010_11000001_01100011_1;
      patterns[41668] = 25'b10100010_11000010_01100100_1;
      patterns[41669] = 25'b10100010_11000011_01100101_1;
      patterns[41670] = 25'b10100010_11000100_01100110_1;
      patterns[41671] = 25'b10100010_11000101_01100111_1;
      patterns[41672] = 25'b10100010_11000110_01101000_1;
      patterns[41673] = 25'b10100010_11000111_01101001_1;
      patterns[41674] = 25'b10100010_11001000_01101010_1;
      patterns[41675] = 25'b10100010_11001001_01101011_1;
      patterns[41676] = 25'b10100010_11001010_01101100_1;
      patterns[41677] = 25'b10100010_11001011_01101101_1;
      patterns[41678] = 25'b10100010_11001100_01101110_1;
      patterns[41679] = 25'b10100010_11001101_01101111_1;
      patterns[41680] = 25'b10100010_11001110_01110000_1;
      patterns[41681] = 25'b10100010_11001111_01110001_1;
      patterns[41682] = 25'b10100010_11010000_01110010_1;
      patterns[41683] = 25'b10100010_11010001_01110011_1;
      patterns[41684] = 25'b10100010_11010010_01110100_1;
      patterns[41685] = 25'b10100010_11010011_01110101_1;
      patterns[41686] = 25'b10100010_11010100_01110110_1;
      patterns[41687] = 25'b10100010_11010101_01110111_1;
      patterns[41688] = 25'b10100010_11010110_01111000_1;
      patterns[41689] = 25'b10100010_11010111_01111001_1;
      patterns[41690] = 25'b10100010_11011000_01111010_1;
      patterns[41691] = 25'b10100010_11011001_01111011_1;
      patterns[41692] = 25'b10100010_11011010_01111100_1;
      patterns[41693] = 25'b10100010_11011011_01111101_1;
      patterns[41694] = 25'b10100010_11011100_01111110_1;
      patterns[41695] = 25'b10100010_11011101_01111111_1;
      patterns[41696] = 25'b10100010_11011110_10000000_1;
      patterns[41697] = 25'b10100010_11011111_10000001_1;
      patterns[41698] = 25'b10100010_11100000_10000010_1;
      patterns[41699] = 25'b10100010_11100001_10000011_1;
      patterns[41700] = 25'b10100010_11100010_10000100_1;
      patterns[41701] = 25'b10100010_11100011_10000101_1;
      patterns[41702] = 25'b10100010_11100100_10000110_1;
      patterns[41703] = 25'b10100010_11100101_10000111_1;
      patterns[41704] = 25'b10100010_11100110_10001000_1;
      patterns[41705] = 25'b10100010_11100111_10001001_1;
      patterns[41706] = 25'b10100010_11101000_10001010_1;
      patterns[41707] = 25'b10100010_11101001_10001011_1;
      patterns[41708] = 25'b10100010_11101010_10001100_1;
      patterns[41709] = 25'b10100010_11101011_10001101_1;
      patterns[41710] = 25'b10100010_11101100_10001110_1;
      patterns[41711] = 25'b10100010_11101101_10001111_1;
      patterns[41712] = 25'b10100010_11101110_10010000_1;
      patterns[41713] = 25'b10100010_11101111_10010001_1;
      patterns[41714] = 25'b10100010_11110000_10010010_1;
      patterns[41715] = 25'b10100010_11110001_10010011_1;
      patterns[41716] = 25'b10100010_11110010_10010100_1;
      patterns[41717] = 25'b10100010_11110011_10010101_1;
      patterns[41718] = 25'b10100010_11110100_10010110_1;
      patterns[41719] = 25'b10100010_11110101_10010111_1;
      patterns[41720] = 25'b10100010_11110110_10011000_1;
      patterns[41721] = 25'b10100010_11110111_10011001_1;
      patterns[41722] = 25'b10100010_11111000_10011010_1;
      patterns[41723] = 25'b10100010_11111001_10011011_1;
      patterns[41724] = 25'b10100010_11111010_10011100_1;
      patterns[41725] = 25'b10100010_11111011_10011101_1;
      patterns[41726] = 25'b10100010_11111100_10011110_1;
      patterns[41727] = 25'b10100010_11111101_10011111_1;
      patterns[41728] = 25'b10100010_11111110_10100000_1;
      patterns[41729] = 25'b10100010_11111111_10100001_1;
      patterns[41730] = 25'b10100011_00000000_10100011_0;
      patterns[41731] = 25'b10100011_00000001_10100100_0;
      patterns[41732] = 25'b10100011_00000010_10100101_0;
      patterns[41733] = 25'b10100011_00000011_10100110_0;
      patterns[41734] = 25'b10100011_00000100_10100111_0;
      patterns[41735] = 25'b10100011_00000101_10101000_0;
      patterns[41736] = 25'b10100011_00000110_10101001_0;
      patterns[41737] = 25'b10100011_00000111_10101010_0;
      patterns[41738] = 25'b10100011_00001000_10101011_0;
      patterns[41739] = 25'b10100011_00001001_10101100_0;
      patterns[41740] = 25'b10100011_00001010_10101101_0;
      patterns[41741] = 25'b10100011_00001011_10101110_0;
      patterns[41742] = 25'b10100011_00001100_10101111_0;
      patterns[41743] = 25'b10100011_00001101_10110000_0;
      patterns[41744] = 25'b10100011_00001110_10110001_0;
      patterns[41745] = 25'b10100011_00001111_10110010_0;
      patterns[41746] = 25'b10100011_00010000_10110011_0;
      patterns[41747] = 25'b10100011_00010001_10110100_0;
      patterns[41748] = 25'b10100011_00010010_10110101_0;
      patterns[41749] = 25'b10100011_00010011_10110110_0;
      patterns[41750] = 25'b10100011_00010100_10110111_0;
      patterns[41751] = 25'b10100011_00010101_10111000_0;
      patterns[41752] = 25'b10100011_00010110_10111001_0;
      patterns[41753] = 25'b10100011_00010111_10111010_0;
      patterns[41754] = 25'b10100011_00011000_10111011_0;
      patterns[41755] = 25'b10100011_00011001_10111100_0;
      patterns[41756] = 25'b10100011_00011010_10111101_0;
      patterns[41757] = 25'b10100011_00011011_10111110_0;
      patterns[41758] = 25'b10100011_00011100_10111111_0;
      patterns[41759] = 25'b10100011_00011101_11000000_0;
      patterns[41760] = 25'b10100011_00011110_11000001_0;
      patterns[41761] = 25'b10100011_00011111_11000010_0;
      patterns[41762] = 25'b10100011_00100000_11000011_0;
      patterns[41763] = 25'b10100011_00100001_11000100_0;
      patterns[41764] = 25'b10100011_00100010_11000101_0;
      patterns[41765] = 25'b10100011_00100011_11000110_0;
      patterns[41766] = 25'b10100011_00100100_11000111_0;
      patterns[41767] = 25'b10100011_00100101_11001000_0;
      patterns[41768] = 25'b10100011_00100110_11001001_0;
      patterns[41769] = 25'b10100011_00100111_11001010_0;
      patterns[41770] = 25'b10100011_00101000_11001011_0;
      patterns[41771] = 25'b10100011_00101001_11001100_0;
      patterns[41772] = 25'b10100011_00101010_11001101_0;
      patterns[41773] = 25'b10100011_00101011_11001110_0;
      patterns[41774] = 25'b10100011_00101100_11001111_0;
      patterns[41775] = 25'b10100011_00101101_11010000_0;
      patterns[41776] = 25'b10100011_00101110_11010001_0;
      patterns[41777] = 25'b10100011_00101111_11010010_0;
      patterns[41778] = 25'b10100011_00110000_11010011_0;
      patterns[41779] = 25'b10100011_00110001_11010100_0;
      patterns[41780] = 25'b10100011_00110010_11010101_0;
      patterns[41781] = 25'b10100011_00110011_11010110_0;
      patterns[41782] = 25'b10100011_00110100_11010111_0;
      patterns[41783] = 25'b10100011_00110101_11011000_0;
      patterns[41784] = 25'b10100011_00110110_11011001_0;
      patterns[41785] = 25'b10100011_00110111_11011010_0;
      patterns[41786] = 25'b10100011_00111000_11011011_0;
      patterns[41787] = 25'b10100011_00111001_11011100_0;
      patterns[41788] = 25'b10100011_00111010_11011101_0;
      patterns[41789] = 25'b10100011_00111011_11011110_0;
      patterns[41790] = 25'b10100011_00111100_11011111_0;
      patterns[41791] = 25'b10100011_00111101_11100000_0;
      patterns[41792] = 25'b10100011_00111110_11100001_0;
      patterns[41793] = 25'b10100011_00111111_11100010_0;
      patterns[41794] = 25'b10100011_01000000_11100011_0;
      patterns[41795] = 25'b10100011_01000001_11100100_0;
      patterns[41796] = 25'b10100011_01000010_11100101_0;
      patterns[41797] = 25'b10100011_01000011_11100110_0;
      patterns[41798] = 25'b10100011_01000100_11100111_0;
      patterns[41799] = 25'b10100011_01000101_11101000_0;
      patterns[41800] = 25'b10100011_01000110_11101001_0;
      patterns[41801] = 25'b10100011_01000111_11101010_0;
      patterns[41802] = 25'b10100011_01001000_11101011_0;
      patterns[41803] = 25'b10100011_01001001_11101100_0;
      patterns[41804] = 25'b10100011_01001010_11101101_0;
      patterns[41805] = 25'b10100011_01001011_11101110_0;
      patterns[41806] = 25'b10100011_01001100_11101111_0;
      patterns[41807] = 25'b10100011_01001101_11110000_0;
      patterns[41808] = 25'b10100011_01001110_11110001_0;
      patterns[41809] = 25'b10100011_01001111_11110010_0;
      patterns[41810] = 25'b10100011_01010000_11110011_0;
      patterns[41811] = 25'b10100011_01010001_11110100_0;
      patterns[41812] = 25'b10100011_01010010_11110101_0;
      patterns[41813] = 25'b10100011_01010011_11110110_0;
      patterns[41814] = 25'b10100011_01010100_11110111_0;
      patterns[41815] = 25'b10100011_01010101_11111000_0;
      patterns[41816] = 25'b10100011_01010110_11111001_0;
      patterns[41817] = 25'b10100011_01010111_11111010_0;
      patterns[41818] = 25'b10100011_01011000_11111011_0;
      patterns[41819] = 25'b10100011_01011001_11111100_0;
      patterns[41820] = 25'b10100011_01011010_11111101_0;
      patterns[41821] = 25'b10100011_01011011_11111110_0;
      patterns[41822] = 25'b10100011_01011100_11111111_0;
      patterns[41823] = 25'b10100011_01011101_00000000_1;
      patterns[41824] = 25'b10100011_01011110_00000001_1;
      patterns[41825] = 25'b10100011_01011111_00000010_1;
      patterns[41826] = 25'b10100011_01100000_00000011_1;
      patterns[41827] = 25'b10100011_01100001_00000100_1;
      patterns[41828] = 25'b10100011_01100010_00000101_1;
      patterns[41829] = 25'b10100011_01100011_00000110_1;
      patterns[41830] = 25'b10100011_01100100_00000111_1;
      patterns[41831] = 25'b10100011_01100101_00001000_1;
      patterns[41832] = 25'b10100011_01100110_00001001_1;
      patterns[41833] = 25'b10100011_01100111_00001010_1;
      patterns[41834] = 25'b10100011_01101000_00001011_1;
      patterns[41835] = 25'b10100011_01101001_00001100_1;
      patterns[41836] = 25'b10100011_01101010_00001101_1;
      patterns[41837] = 25'b10100011_01101011_00001110_1;
      patterns[41838] = 25'b10100011_01101100_00001111_1;
      patterns[41839] = 25'b10100011_01101101_00010000_1;
      patterns[41840] = 25'b10100011_01101110_00010001_1;
      patterns[41841] = 25'b10100011_01101111_00010010_1;
      patterns[41842] = 25'b10100011_01110000_00010011_1;
      patterns[41843] = 25'b10100011_01110001_00010100_1;
      patterns[41844] = 25'b10100011_01110010_00010101_1;
      patterns[41845] = 25'b10100011_01110011_00010110_1;
      patterns[41846] = 25'b10100011_01110100_00010111_1;
      patterns[41847] = 25'b10100011_01110101_00011000_1;
      patterns[41848] = 25'b10100011_01110110_00011001_1;
      patterns[41849] = 25'b10100011_01110111_00011010_1;
      patterns[41850] = 25'b10100011_01111000_00011011_1;
      patterns[41851] = 25'b10100011_01111001_00011100_1;
      patterns[41852] = 25'b10100011_01111010_00011101_1;
      patterns[41853] = 25'b10100011_01111011_00011110_1;
      patterns[41854] = 25'b10100011_01111100_00011111_1;
      patterns[41855] = 25'b10100011_01111101_00100000_1;
      patterns[41856] = 25'b10100011_01111110_00100001_1;
      patterns[41857] = 25'b10100011_01111111_00100010_1;
      patterns[41858] = 25'b10100011_10000000_00100011_1;
      patterns[41859] = 25'b10100011_10000001_00100100_1;
      patterns[41860] = 25'b10100011_10000010_00100101_1;
      patterns[41861] = 25'b10100011_10000011_00100110_1;
      patterns[41862] = 25'b10100011_10000100_00100111_1;
      patterns[41863] = 25'b10100011_10000101_00101000_1;
      patterns[41864] = 25'b10100011_10000110_00101001_1;
      patterns[41865] = 25'b10100011_10000111_00101010_1;
      patterns[41866] = 25'b10100011_10001000_00101011_1;
      patterns[41867] = 25'b10100011_10001001_00101100_1;
      patterns[41868] = 25'b10100011_10001010_00101101_1;
      patterns[41869] = 25'b10100011_10001011_00101110_1;
      patterns[41870] = 25'b10100011_10001100_00101111_1;
      patterns[41871] = 25'b10100011_10001101_00110000_1;
      patterns[41872] = 25'b10100011_10001110_00110001_1;
      patterns[41873] = 25'b10100011_10001111_00110010_1;
      patterns[41874] = 25'b10100011_10010000_00110011_1;
      patterns[41875] = 25'b10100011_10010001_00110100_1;
      patterns[41876] = 25'b10100011_10010010_00110101_1;
      patterns[41877] = 25'b10100011_10010011_00110110_1;
      patterns[41878] = 25'b10100011_10010100_00110111_1;
      patterns[41879] = 25'b10100011_10010101_00111000_1;
      patterns[41880] = 25'b10100011_10010110_00111001_1;
      patterns[41881] = 25'b10100011_10010111_00111010_1;
      patterns[41882] = 25'b10100011_10011000_00111011_1;
      patterns[41883] = 25'b10100011_10011001_00111100_1;
      patterns[41884] = 25'b10100011_10011010_00111101_1;
      patterns[41885] = 25'b10100011_10011011_00111110_1;
      patterns[41886] = 25'b10100011_10011100_00111111_1;
      patterns[41887] = 25'b10100011_10011101_01000000_1;
      patterns[41888] = 25'b10100011_10011110_01000001_1;
      patterns[41889] = 25'b10100011_10011111_01000010_1;
      patterns[41890] = 25'b10100011_10100000_01000011_1;
      patterns[41891] = 25'b10100011_10100001_01000100_1;
      patterns[41892] = 25'b10100011_10100010_01000101_1;
      patterns[41893] = 25'b10100011_10100011_01000110_1;
      patterns[41894] = 25'b10100011_10100100_01000111_1;
      patterns[41895] = 25'b10100011_10100101_01001000_1;
      patterns[41896] = 25'b10100011_10100110_01001001_1;
      patterns[41897] = 25'b10100011_10100111_01001010_1;
      patterns[41898] = 25'b10100011_10101000_01001011_1;
      patterns[41899] = 25'b10100011_10101001_01001100_1;
      patterns[41900] = 25'b10100011_10101010_01001101_1;
      patterns[41901] = 25'b10100011_10101011_01001110_1;
      patterns[41902] = 25'b10100011_10101100_01001111_1;
      patterns[41903] = 25'b10100011_10101101_01010000_1;
      patterns[41904] = 25'b10100011_10101110_01010001_1;
      patterns[41905] = 25'b10100011_10101111_01010010_1;
      patterns[41906] = 25'b10100011_10110000_01010011_1;
      patterns[41907] = 25'b10100011_10110001_01010100_1;
      patterns[41908] = 25'b10100011_10110010_01010101_1;
      patterns[41909] = 25'b10100011_10110011_01010110_1;
      patterns[41910] = 25'b10100011_10110100_01010111_1;
      patterns[41911] = 25'b10100011_10110101_01011000_1;
      patterns[41912] = 25'b10100011_10110110_01011001_1;
      patterns[41913] = 25'b10100011_10110111_01011010_1;
      patterns[41914] = 25'b10100011_10111000_01011011_1;
      patterns[41915] = 25'b10100011_10111001_01011100_1;
      patterns[41916] = 25'b10100011_10111010_01011101_1;
      patterns[41917] = 25'b10100011_10111011_01011110_1;
      patterns[41918] = 25'b10100011_10111100_01011111_1;
      patterns[41919] = 25'b10100011_10111101_01100000_1;
      patterns[41920] = 25'b10100011_10111110_01100001_1;
      patterns[41921] = 25'b10100011_10111111_01100010_1;
      patterns[41922] = 25'b10100011_11000000_01100011_1;
      patterns[41923] = 25'b10100011_11000001_01100100_1;
      patterns[41924] = 25'b10100011_11000010_01100101_1;
      patterns[41925] = 25'b10100011_11000011_01100110_1;
      patterns[41926] = 25'b10100011_11000100_01100111_1;
      patterns[41927] = 25'b10100011_11000101_01101000_1;
      patterns[41928] = 25'b10100011_11000110_01101001_1;
      patterns[41929] = 25'b10100011_11000111_01101010_1;
      patterns[41930] = 25'b10100011_11001000_01101011_1;
      patterns[41931] = 25'b10100011_11001001_01101100_1;
      patterns[41932] = 25'b10100011_11001010_01101101_1;
      patterns[41933] = 25'b10100011_11001011_01101110_1;
      patterns[41934] = 25'b10100011_11001100_01101111_1;
      patterns[41935] = 25'b10100011_11001101_01110000_1;
      patterns[41936] = 25'b10100011_11001110_01110001_1;
      patterns[41937] = 25'b10100011_11001111_01110010_1;
      patterns[41938] = 25'b10100011_11010000_01110011_1;
      patterns[41939] = 25'b10100011_11010001_01110100_1;
      patterns[41940] = 25'b10100011_11010010_01110101_1;
      patterns[41941] = 25'b10100011_11010011_01110110_1;
      patterns[41942] = 25'b10100011_11010100_01110111_1;
      patterns[41943] = 25'b10100011_11010101_01111000_1;
      patterns[41944] = 25'b10100011_11010110_01111001_1;
      patterns[41945] = 25'b10100011_11010111_01111010_1;
      patterns[41946] = 25'b10100011_11011000_01111011_1;
      patterns[41947] = 25'b10100011_11011001_01111100_1;
      patterns[41948] = 25'b10100011_11011010_01111101_1;
      patterns[41949] = 25'b10100011_11011011_01111110_1;
      patterns[41950] = 25'b10100011_11011100_01111111_1;
      patterns[41951] = 25'b10100011_11011101_10000000_1;
      patterns[41952] = 25'b10100011_11011110_10000001_1;
      patterns[41953] = 25'b10100011_11011111_10000010_1;
      patterns[41954] = 25'b10100011_11100000_10000011_1;
      patterns[41955] = 25'b10100011_11100001_10000100_1;
      patterns[41956] = 25'b10100011_11100010_10000101_1;
      patterns[41957] = 25'b10100011_11100011_10000110_1;
      patterns[41958] = 25'b10100011_11100100_10000111_1;
      patterns[41959] = 25'b10100011_11100101_10001000_1;
      patterns[41960] = 25'b10100011_11100110_10001001_1;
      patterns[41961] = 25'b10100011_11100111_10001010_1;
      patterns[41962] = 25'b10100011_11101000_10001011_1;
      patterns[41963] = 25'b10100011_11101001_10001100_1;
      patterns[41964] = 25'b10100011_11101010_10001101_1;
      patterns[41965] = 25'b10100011_11101011_10001110_1;
      patterns[41966] = 25'b10100011_11101100_10001111_1;
      patterns[41967] = 25'b10100011_11101101_10010000_1;
      patterns[41968] = 25'b10100011_11101110_10010001_1;
      patterns[41969] = 25'b10100011_11101111_10010010_1;
      patterns[41970] = 25'b10100011_11110000_10010011_1;
      patterns[41971] = 25'b10100011_11110001_10010100_1;
      patterns[41972] = 25'b10100011_11110010_10010101_1;
      patterns[41973] = 25'b10100011_11110011_10010110_1;
      patterns[41974] = 25'b10100011_11110100_10010111_1;
      patterns[41975] = 25'b10100011_11110101_10011000_1;
      patterns[41976] = 25'b10100011_11110110_10011001_1;
      patterns[41977] = 25'b10100011_11110111_10011010_1;
      patterns[41978] = 25'b10100011_11111000_10011011_1;
      patterns[41979] = 25'b10100011_11111001_10011100_1;
      patterns[41980] = 25'b10100011_11111010_10011101_1;
      patterns[41981] = 25'b10100011_11111011_10011110_1;
      patterns[41982] = 25'b10100011_11111100_10011111_1;
      patterns[41983] = 25'b10100011_11111101_10100000_1;
      patterns[41984] = 25'b10100011_11111110_10100001_1;
      patterns[41985] = 25'b10100011_11111111_10100010_1;
      patterns[41986] = 25'b10100100_00000000_10100100_0;
      patterns[41987] = 25'b10100100_00000001_10100101_0;
      patterns[41988] = 25'b10100100_00000010_10100110_0;
      patterns[41989] = 25'b10100100_00000011_10100111_0;
      patterns[41990] = 25'b10100100_00000100_10101000_0;
      patterns[41991] = 25'b10100100_00000101_10101001_0;
      patterns[41992] = 25'b10100100_00000110_10101010_0;
      patterns[41993] = 25'b10100100_00000111_10101011_0;
      patterns[41994] = 25'b10100100_00001000_10101100_0;
      patterns[41995] = 25'b10100100_00001001_10101101_0;
      patterns[41996] = 25'b10100100_00001010_10101110_0;
      patterns[41997] = 25'b10100100_00001011_10101111_0;
      patterns[41998] = 25'b10100100_00001100_10110000_0;
      patterns[41999] = 25'b10100100_00001101_10110001_0;
      patterns[42000] = 25'b10100100_00001110_10110010_0;
      patterns[42001] = 25'b10100100_00001111_10110011_0;
      patterns[42002] = 25'b10100100_00010000_10110100_0;
      patterns[42003] = 25'b10100100_00010001_10110101_0;
      patterns[42004] = 25'b10100100_00010010_10110110_0;
      patterns[42005] = 25'b10100100_00010011_10110111_0;
      patterns[42006] = 25'b10100100_00010100_10111000_0;
      patterns[42007] = 25'b10100100_00010101_10111001_0;
      patterns[42008] = 25'b10100100_00010110_10111010_0;
      patterns[42009] = 25'b10100100_00010111_10111011_0;
      patterns[42010] = 25'b10100100_00011000_10111100_0;
      patterns[42011] = 25'b10100100_00011001_10111101_0;
      patterns[42012] = 25'b10100100_00011010_10111110_0;
      patterns[42013] = 25'b10100100_00011011_10111111_0;
      patterns[42014] = 25'b10100100_00011100_11000000_0;
      patterns[42015] = 25'b10100100_00011101_11000001_0;
      patterns[42016] = 25'b10100100_00011110_11000010_0;
      patterns[42017] = 25'b10100100_00011111_11000011_0;
      patterns[42018] = 25'b10100100_00100000_11000100_0;
      patterns[42019] = 25'b10100100_00100001_11000101_0;
      patterns[42020] = 25'b10100100_00100010_11000110_0;
      patterns[42021] = 25'b10100100_00100011_11000111_0;
      patterns[42022] = 25'b10100100_00100100_11001000_0;
      patterns[42023] = 25'b10100100_00100101_11001001_0;
      patterns[42024] = 25'b10100100_00100110_11001010_0;
      patterns[42025] = 25'b10100100_00100111_11001011_0;
      patterns[42026] = 25'b10100100_00101000_11001100_0;
      patterns[42027] = 25'b10100100_00101001_11001101_0;
      patterns[42028] = 25'b10100100_00101010_11001110_0;
      patterns[42029] = 25'b10100100_00101011_11001111_0;
      patterns[42030] = 25'b10100100_00101100_11010000_0;
      patterns[42031] = 25'b10100100_00101101_11010001_0;
      patterns[42032] = 25'b10100100_00101110_11010010_0;
      patterns[42033] = 25'b10100100_00101111_11010011_0;
      patterns[42034] = 25'b10100100_00110000_11010100_0;
      patterns[42035] = 25'b10100100_00110001_11010101_0;
      patterns[42036] = 25'b10100100_00110010_11010110_0;
      patterns[42037] = 25'b10100100_00110011_11010111_0;
      patterns[42038] = 25'b10100100_00110100_11011000_0;
      patterns[42039] = 25'b10100100_00110101_11011001_0;
      patterns[42040] = 25'b10100100_00110110_11011010_0;
      patterns[42041] = 25'b10100100_00110111_11011011_0;
      patterns[42042] = 25'b10100100_00111000_11011100_0;
      patterns[42043] = 25'b10100100_00111001_11011101_0;
      patterns[42044] = 25'b10100100_00111010_11011110_0;
      patterns[42045] = 25'b10100100_00111011_11011111_0;
      patterns[42046] = 25'b10100100_00111100_11100000_0;
      patterns[42047] = 25'b10100100_00111101_11100001_0;
      patterns[42048] = 25'b10100100_00111110_11100010_0;
      patterns[42049] = 25'b10100100_00111111_11100011_0;
      patterns[42050] = 25'b10100100_01000000_11100100_0;
      patterns[42051] = 25'b10100100_01000001_11100101_0;
      patterns[42052] = 25'b10100100_01000010_11100110_0;
      patterns[42053] = 25'b10100100_01000011_11100111_0;
      patterns[42054] = 25'b10100100_01000100_11101000_0;
      patterns[42055] = 25'b10100100_01000101_11101001_0;
      patterns[42056] = 25'b10100100_01000110_11101010_0;
      patterns[42057] = 25'b10100100_01000111_11101011_0;
      patterns[42058] = 25'b10100100_01001000_11101100_0;
      patterns[42059] = 25'b10100100_01001001_11101101_0;
      patterns[42060] = 25'b10100100_01001010_11101110_0;
      patterns[42061] = 25'b10100100_01001011_11101111_0;
      patterns[42062] = 25'b10100100_01001100_11110000_0;
      patterns[42063] = 25'b10100100_01001101_11110001_0;
      patterns[42064] = 25'b10100100_01001110_11110010_0;
      patterns[42065] = 25'b10100100_01001111_11110011_0;
      patterns[42066] = 25'b10100100_01010000_11110100_0;
      patterns[42067] = 25'b10100100_01010001_11110101_0;
      patterns[42068] = 25'b10100100_01010010_11110110_0;
      patterns[42069] = 25'b10100100_01010011_11110111_0;
      patterns[42070] = 25'b10100100_01010100_11111000_0;
      patterns[42071] = 25'b10100100_01010101_11111001_0;
      patterns[42072] = 25'b10100100_01010110_11111010_0;
      patterns[42073] = 25'b10100100_01010111_11111011_0;
      patterns[42074] = 25'b10100100_01011000_11111100_0;
      patterns[42075] = 25'b10100100_01011001_11111101_0;
      patterns[42076] = 25'b10100100_01011010_11111110_0;
      patterns[42077] = 25'b10100100_01011011_11111111_0;
      patterns[42078] = 25'b10100100_01011100_00000000_1;
      patterns[42079] = 25'b10100100_01011101_00000001_1;
      patterns[42080] = 25'b10100100_01011110_00000010_1;
      patterns[42081] = 25'b10100100_01011111_00000011_1;
      patterns[42082] = 25'b10100100_01100000_00000100_1;
      patterns[42083] = 25'b10100100_01100001_00000101_1;
      patterns[42084] = 25'b10100100_01100010_00000110_1;
      patterns[42085] = 25'b10100100_01100011_00000111_1;
      patterns[42086] = 25'b10100100_01100100_00001000_1;
      patterns[42087] = 25'b10100100_01100101_00001001_1;
      patterns[42088] = 25'b10100100_01100110_00001010_1;
      patterns[42089] = 25'b10100100_01100111_00001011_1;
      patterns[42090] = 25'b10100100_01101000_00001100_1;
      patterns[42091] = 25'b10100100_01101001_00001101_1;
      patterns[42092] = 25'b10100100_01101010_00001110_1;
      patterns[42093] = 25'b10100100_01101011_00001111_1;
      patterns[42094] = 25'b10100100_01101100_00010000_1;
      patterns[42095] = 25'b10100100_01101101_00010001_1;
      patterns[42096] = 25'b10100100_01101110_00010010_1;
      patterns[42097] = 25'b10100100_01101111_00010011_1;
      patterns[42098] = 25'b10100100_01110000_00010100_1;
      patterns[42099] = 25'b10100100_01110001_00010101_1;
      patterns[42100] = 25'b10100100_01110010_00010110_1;
      patterns[42101] = 25'b10100100_01110011_00010111_1;
      patterns[42102] = 25'b10100100_01110100_00011000_1;
      patterns[42103] = 25'b10100100_01110101_00011001_1;
      patterns[42104] = 25'b10100100_01110110_00011010_1;
      patterns[42105] = 25'b10100100_01110111_00011011_1;
      patterns[42106] = 25'b10100100_01111000_00011100_1;
      patterns[42107] = 25'b10100100_01111001_00011101_1;
      patterns[42108] = 25'b10100100_01111010_00011110_1;
      patterns[42109] = 25'b10100100_01111011_00011111_1;
      patterns[42110] = 25'b10100100_01111100_00100000_1;
      patterns[42111] = 25'b10100100_01111101_00100001_1;
      patterns[42112] = 25'b10100100_01111110_00100010_1;
      patterns[42113] = 25'b10100100_01111111_00100011_1;
      patterns[42114] = 25'b10100100_10000000_00100100_1;
      patterns[42115] = 25'b10100100_10000001_00100101_1;
      patterns[42116] = 25'b10100100_10000010_00100110_1;
      patterns[42117] = 25'b10100100_10000011_00100111_1;
      patterns[42118] = 25'b10100100_10000100_00101000_1;
      patterns[42119] = 25'b10100100_10000101_00101001_1;
      patterns[42120] = 25'b10100100_10000110_00101010_1;
      patterns[42121] = 25'b10100100_10000111_00101011_1;
      patterns[42122] = 25'b10100100_10001000_00101100_1;
      patterns[42123] = 25'b10100100_10001001_00101101_1;
      patterns[42124] = 25'b10100100_10001010_00101110_1;
      patterns[42125] = 25'b10100100_10001011_00101111_1;
      patterns[42126] = 25'b10100100_10001100_00110000_1;
      patterns[42127] = 25'b10100100_10001101_00110001_1;
      patterns[42128] = 25'b10100100_10001110_00110010_1;
      patterns[42129] = 25'b10100100_10001111_00110011_1;
      patterns[42130] = 25'b10100100_10010000_00110100_1;
      patterns[42131] = 25'b10100100_10010001_00110101_1;
      patterns[42132] = 25'b10100100_10010010_00110110_1;
      patterns[42133] = 25'b10100100_10010011_00110111_1;
      patterns[42134] = 25'b10100100_10010100_00111000_1;
      patterns[42135] = 25'b10100100_10010101_00111001_1;
      patterns[42136] = 25'b10100100_10010110_00111010_1;
      patterns[42137] = 25'b10100100_10010111_00111011_1;
      patterns[42138] = 25'b10100100_10011000_00111100_1;
      patterns[42139] = 25'b10100100_10011001_00111101_1;
      patterns[42140] = 25'b10100100_10011010_00111110_1;
      patterns[42141] = 25'b10100100_10011011_00111111_1;
      patterns[42142] = 25'b10100100_10011100_01000000_1;
      patterns[42143] = 25'b10100100_10011101_01000001_1;
      patterns[42144] = 25'b10100100_10011110_01000010_1;
      patterns[42145] = 25'b10100100_10011111_01000011_1;
      patterns[42146] = 25'b10100100_10100000_01000100_1;
      patterns[42147] = 25'b10100100_10100001_01000101_1;
      patterns[42148] = 25'b10100100_10100010_01000110_1;
      patterns[42149] = 25'b10100100_10100011_01000111_1;
      patterns[42150] = 25'b10100100_10100100_01001000_1;
      patterns[42151] = 25'b10100100_10100101_01001001_1;
      patterns[42152] = 25'b10100100_10100110_01001010_1;
      patterns[42153] = 25'b10100100_10100111_01001011_1;
      patterns[42154] = 25'b10100100_10101000_01001100_1;
      patterns[42155] = 25'b10100100_10101001_01001101_1;
      patterns[42156] = 25'b10100100_10101010_01001110_1;
      patterns[42157] = 25'b10100100_10101011_01001111_1;
      patterns[42158] = 25'b10100100_10101100_01010000_1;
      patterns[42159] = 25'b10100100_10101101_01010001_1;
      patterns[42160] = 25'b10100100_10101110_01010010_1;
      patterns[42161] = 25'b10100100_10101111_01010011_1;
      patterns[42162] = 25'b10100100_10110000_01010100_1;
      patterns[42163] = 25'b10100100_10110001_01010101_1;
      patterns[42164] = 25'b10100100_10110010_01010110_1;
      patterns[42165] = 25'b10100100_10110011_01010111_1;
      patterns[42166] = 25'b10100100_10110100_01011000_1;
      patterns[42167] = 25'b10100100_10110101_01011001_1;
      patterns[42168] = 25'b10100100_10110110_01011010_1;
      patterns[42169] = 25'b10100100_10110111_01011011_1;
      patterns[42170] = 25'b10100100_10111000_01011100_1;
      patterns[42171] = 25'b10100100_10111001_01011101_1;
      patterns[42172] = 25'b10100100_10111010_01011110_1;
      patterns[42173] = 25'b10100100_10111011_01011111_1;
      patterns[42174] = 25'b10100100_10111100_01100000_1;
      patterns[42175] = 25'b10100100_10111101_01100001_1;
      patterns[42176] = 25'b10100100_10111110_01100010_1;
      patterns[42177] = 25'b10100100_10111111_01100011_1;
      patterns[42178] = 25'b10100100_11000000_01100100_1;
      patterns[42179] = 25'b10100100_11000001_01100101_1;
      patterns[42180] = 25'b10100100_11000010_01100110_1;
      patterns[42181] = 25'b10100100_11000011_01100111_1;
      patterns[42182] = 25'b10100100_11000100_01101000_1;
      patterns[42183] = 25'b10100100_11000101_01101001_1;
      patterns[42184] = 25'b10100100_11000110_01101010_1;
      patterns[42185] = 25'b10100100_11000111_01101011_1;
      patterns[42186] = 25'b10100100_11001000_01101100_1;
      patterns[42187] = 25'b10100100_11001001_01101101_1;
      patterns[42188] = 25'b10100100_11001010_01101110_1;
      patterns[42189] = 25'b10100100_11001011_01101111_1;
      patterns[42190] = 25'b10100100_11001100_01110000_1;
      patterns[42191] = 25'b10100100_11001101_01110001_1;
      patterns[42192] = 25'b10100100_11001110_01110010_1;
      patterns[42193] = 25'b10100100_11001111_01110011_1;
      patterns[42194] = 25'b10100100_11010000_01110100_1;
      patterns[42195] = 25'b10100100_11010001_01110101_1;
      patterns[42196] = 25'b10100100_11010010_01110110_1;
      patterns[42197] = 25'b10100100_11010011_01110111_1;
      patterns[42198] = 25'b10100100_11010100_01111000_1;
      patterns[42199] = 25'b10100100_11010101_01111001_1;
      patterns[42200] = 25'b10100100_11010110_01111010_1;
      patterns[42201] = 25'b10100100_11010111_01111011_1;
      patterns[42202] = 25'b10100100_11011000_01111100_1;
      patterns[42203] = 25'b10100100_11011001_01111101_1;
      patterns[42204] = 25'b10100100_11011010_01111110_1;
      patterns[42205] = 25'b10100100_11011011_01111111_1;
      patterns[42206] = 25'b10100100_11011100_10000000_1;
      patterns[42207] = 25'b10100100_11011101_10000001_1;
      patterns[42208] = 25'b10100100_11011110_10000010_1;
      patterns[42209] = 25'b10100100_11011111_10000011_1;
      patterns[42210] = 25'b10100100_11100000_10000100_1;
      patterns[42211] = 25'b10100100_11100001_10000101_1;
      patterns[42212] = 25'b10100100_11100010_10000110_1;
      patterns[42213] = 25'b10100100_11100011_10000111_1;
      patterns[42214] = 25'b10100100_11100100_10001000_1;
      patterns[42215] = 25'b10100100_11100101_10001001_1;
      patterns[42216] = 25'b10100100_11100110_10001010_1;
      patterns[42217] = 25'b10100100_11100111_10001011_1;
      patterns[42218] = 25'b10100100_11101000_10001100_1;
      patterns[42219] = 25'b10100100_11101001_10001101_1;
      patterns[42220] = 25'b10100100_11101010_10001110_1;
      patterns[42221] = 25'b10100100_11101011_10001111_1;
      patterns[42222] = 25'b10100100_11101100_10010000_1;
      patterns[42223] = 25'b10100100_11101101_10010001_1;
      patterns[42224] = 25'b10100100_11101110_10010010_1;
      patterns[42225] = 25'b10100100_11101111_10010011_1;
      patterns[42226] = 25'b10100100_11110000_10010100_1;
      patterns[42227] = 25'b10100100_11110001_10010101_1;
      patterns[42228] = 25'b10100100_11110010_10010110_1;
      patterns[42229] = 25'b10100100_11110011_10010111_1;
      patterns[42230] = 25'b10100100_11110100_10011000_1;
      patterns[42231] = 25'b10100100_11110101_10011001_1;
      patterns[42232] = 25'b10100100_11110110_10011010_1;
      patterns[42233] = 25'b10100100_11110111_10011011_1;
      patterns[42234] = 25'b10100100_11111000_10011100_1;
      patterns[42235] = 25'b10100100_11111001_10011101_1;
      patterns[42236] = 25'b10100100_11111010_10011110_1;
      patterns[42237] = 25'b10100100_11111011_10011111_1;
      patterns[42238] = 25'b10100100_11111100_10100000_1;
      patterns[42239] = 25'b10100100_11111101_10100001_1;
      patterns[42240] = 25'b10100100_11111110_10100010_1;
      patterns[42241] = 25'b10100100_11111111_10100011_1;
      patterns[42242] = 25'b10100101_00000000_10100101_0;
      patterns[42243] = 25'b10100101_00000001_10100110_0;
      patterns[42244] = 25'b10100101_00000010_10100111_0;
      patterns[42245] = 25'b10100101_00000011_10101000_0;
      patterns[42246] = 25'b10100101_00000100_10101001_0;
      patterns[42247] = 25'b10100101_00000101_10101010_0;
      patterns[42248] = 25'b10100101_00000110_10101011_0;
      patterns[42249] = 25'b10100101_00000111_10101100_0;
      patterns[42250] = 25'b10100101_00001000_10101101_0;
      patterns[42251] = 25'b10100101_00001001_10101110_0;
      patterns[42252] = 25'b10100101_00001010_10101111_0;
      patterns[42253] = 25'b10100101_00001011_10110000_0;
      patterns[42254] = 25'b10100101_00001100_10110001_0;
      patterns[42255] = 25'b10100101_00001101_10110010_0;
      patterns[42256] = 25'b10100101_00001110_10110011_0;
      patterns[42257] = 25'b10100101_00001111_10110100_0;
      patterns[42258] = 25'b10100101_00010000_10110101_0;
      patterns[42259] = 25'b10100101_00010001_10110110_0;
      patterns[42260] = 25'b10100101_00010010_10110111_0;
      patterns[42261] = 25'b10100101_00010011_10111000_0;
      patterns[42262] = 25'b10100101_00010100_10111001_0;
      patterns[42263] = 25'b10100101_00010101_10111010_0;
      patterns[42264] = 25'b10100101_00010110_10111011_0;
      patterns[42265] = 25'b10100101_00010111_10111100_0;
      patterns[42266] = 25'b10100101_00011000_10111101_0;
      patterns[42267] = 25'b10100101_00011001_10111110_0;
      patterns[42268] = 25'b10100101_00011010_10111111_0;
      patterns[42269] = 25'b10100101_00011011_11000000_0;
      patterns[42270] = 25'b10100101_00011100_11000001_0;
      patterns[42271] = 25'b10100101_00011101_11000010_0;
      patterns[42272] = 25'b10100101_00011110_11000011_0;
      patterns[42273] = 25'b10100101_00011111_11000100_0;
      patterns[42274] = 25'b10100101_00100000_11000101_0;
      patterns[42275] = 25'b10100101_00100001_11000110_0;
      patterns[42276] = 25'b10100101_00100010_11000111_0;
      patterns[42277] = 25'b10100101_00100011_11001000_0;
      patterns[42278] = 25'b10100101_00100100_11001001_0;
      patterns[42279] = 25'b10100101_00100101_11001010_0;
      patterns[42280] = 25'b10100101_00100110_11001011_0;
      patterns[42281] = 25'b10100101_00100111_11001100_0;
      patterns[42282] = 25'b10100101_00101000_11001101_0;
      patterns[42283] = 25'b10100101_00101001_11001110_0;
      patterns[42284] = 25'b10100101_00101010_11001111_0;
      patterns[42285] = 25'b10100101_00101011_11010000_0;
      patterns[42286] = 25'b10100101_00101100_11010001_0;
      patterns[42287] = 25'b10100101_00101101_11010010_0;
      patterns[42288] = 25'b10100101_00101110_11010011_0;
      patterns[42289] = 25'b10100101_00101111_11010100_0;
      patterns[42290] = 25'b10100101_00110000_11010101_0;
      patterns[42291] = 25'b10100101_00110001_11010110_0;
      patterns[42292] = 25'b10100101_00110010_11010111_0;
      patterns[42293] = 25'b10100101_00110011_11011000_0;
      patterns[42294] = 25'b10100101_00110100_11011001_0;
      patterns[42295] = 25'b10100101_00110101_11011010_0;
      patterns[42296] = 25'b10100101_00110110_11011011_0;
      patterns[42297] = 25'b10100101_00110111_11011100_0;
      patterns[42298] = 25'b10100101_00111000_11011101_0;
      patterns[42299] = 25'b10100101_00111001_11011110_0;
      patterns[42300] = 25'b10100101_00111010_11011111_0;
      patterns[42301] = 25'b10100101_00111011_11100000_0;
      patterns[42302] = 25'b10100101_00111100_11100001_0;
      patterns[42303] = 25'b10100101_00111101_11100010_0;
      patterns[42304] = 25'b10100101_00111110_11100011_0;
      patterns[42305] = 25'b10100101_00111111_11100100_0;
      patterns[42306] = 25'b10100101_01000000_11100101_0;
      patterns[42307] = 25'b10100101_01000001_11100110_0;
      patterns[42308] = 25'b10100101_01000010_11100111_0;
      patterns[42309] = 25'b10100101_01000011_11101000_0;
      patterns[42310] = 25'b10100101_01000100_11101001_0;
      patterns[42311] = 25'b10100101_01000101_11101010_0;
      patterns[42312] = 25'b10100101_01000110_11101011_0;
      patterns[42313] = 25'b10100101_01000111_11101100_0;
      patterns[42314] = 25'b10100101_01001000_11101101_0;
      patterns[42315] = 25'b10100101_01001001_11101110_0;
      patterns[42316] = 25'b10100101_01001010_11101111_0;
      patterns[42317] = 25'b10100101_01001011_11110000_0;
      patterns[42318] = 25'b10100101_01001100_11110001_0;
      patterns[42319] = 25'b10100101_01001101_11110010_0;
      patterns[42320] = 25'b10100101_01001110_11110011_0;
      patterns[42321] = 25'b10100101_01001111_11110100_0;
      patterns[42322] = 25'b10100101_01010000_11110101_0;
      patterns[42323] = 25'b10100101_01010001_11110110_0;
      patterns[42324] = 25'b10100101_01010010_11110111_0;
      patterns[42325] = 25'b10100101_01010011_11111000_0;
      patterns[42326] = 25'b10100101_01010100_11111001_0;
      patterns[42327] = 25'b10100101_01010101_11111010_0;
      patterns[42328] = 25'b10100101_01010110_11111011_0;
      patterns[42329] = 25'b10100101_01010111_11111100_0;
      patterns[42330] = 25'b10100101_01011000_11111101_0;
      patterns[42331] = 25'b10100101_01011001_11111110_0;
      patterns[42332] = 25'b10100101_01011010_11111111_0;
      patterns[42333] = 25'b10100101_01011011_00000000_1;
      patterns[42334] = 25'b10100101_01011100_00000001_1;
      patterns[42335] = 25'b10100101_01011101_00000010_1;
      patterns[42336] = 25'b10100101_01011110_00000011_1;
      patterns[42337] = 25'b10100101_01011111_00000100_1;
      patterns[42338] = 25'b10100101_01100000_00000101_1;
      patterns[42339] = 25'b10100101_01100001_00000110_1;
      patterns[42340] = 25'b10100101_01100010_00000111_1;
      patterns[42341] = 25'b10100101_01100011_00001000_1;
      patterns[42342] = 25'b10100101_01100100_00001001_1;
      patterns[42343] = 25'b10100101_01100101_00001010_1;
      patterns[42344] = 25'b10100101_01100110_00001011_1;
      patterns[42345] = 25'b10100101_01100111_00001100_1;
      patterns[42346] = 25'b10100101_01101000_00001101_1;
      patterns[42347] = 25'b10100101_01101001_00001110_1;
      patterns[42348] = 25'b10100101_01101010_00001111_1;
      patterns[42349] = 25'b10100101_01101011_00010000_1;
      patterns[42350] = 25'b10100101_01101100_00010001_1;
      patterns[42351] = 25'b10100101_01101101_00010010_1;
      patterns[42352] = 25'b10100101_01101110_00010011_1;
      patterns[42353] = 25'b10100101_01101111_00010100_1;
      patterns[42354] = 25'b10100101_01110000_00010101_1;
      patterns[42355] = 25'b10100101_01110001_00010110_1;
      patterns[42356] = 25'b10100101_01110010_00010111_1;
      patterns[42357] = 25'b10100101_01110011_00011000_1;
      patterns[42358] = 25'b10100101_01110100_00011001_1;
      patterns[42359] = 25'b10100101_01110101_00011010_1;
      patterns[42360] = 25'b10100101_01110110_00011011_1;
      patterns[42361] = 25'b10100101_01110111_00011100_1;
      patterns[42362] = 25'b10100101_01111000_00011101_1;
      patterns[42363] = 25'b10100101_01111001_00011110_1;
      patterns[42364] = 25'b10100101_01111010_00011111_1;
      patterns[42365] = 25'b10100101_01111011_00100000_1;
      patterns[42366] = 25'b10100101_01111100_00100001_1;
      patterns[42367] = 25'b10100101_01111101_00100010_1;
      patterns[42368] = 25'b10100101_01111110_00100011_1;
      patterns[42369] = 25'b10100101_01111111_00100100_1;
      patterns[42370] = 25'b10100101_10000000_00100101_1;
      patterns[42371] = 25'b10100101_10000001_00100110_1;
      patterns[42372] = 25'b10100101_10000010_00100111_1;
      patterns[42373] = 25'b10100101_10000011_00101000_1;
      patterns[42374] = 25'b10100101_10000100_00101001_1;
      patterns[42375] = 25'b10100101_10000101_00101010_1;
      patterns[42376] = 25'b10100101_10000110_00101011_1;
      patterns[42377] = 25'b10100101_10000111_00101100_1;
      patterns[42378] = 25'b10100101_10001000_00101101_1;
      patterns[42379] = 25'b10100101_10001001_00101110_1;
      patterns[42380] = 25'b10100101_10001010_00101111_1;
      patterns[42381] = 25'b10100101_10001011_00110000_1;
      patterns[42382] = 25'b10100101_10001100_00110001_1;
      patterns[42383] = 25'b10100101_10001101_00110010_1;
      patterns[42384] = 25'b10100101_10001110_00110011_1;
      patterns[42385] = 25'b10100101_10001111_00110100_1;
      patterns[42386] = 25'b10100101_10010000_00110101_1;
      patterns[42387] = 25'b10100101_10010001_00110110_1;
      patterns[42388] = 25'b10100101_10010010_00110111_1;
      patterns[42389] = 25'b10100101_10010011_00111000_1;
      patterns[42390] = 25'b10100101_10010100_00111001_1;
      patterns[42391] = 25'b10100101_10010101_00111010_1;
      patterns[42392] = 25'b10100101_10010110_00111011_1;
      patterns[42393] = 25'b10100101_10010111_00111100_1;
      patterns[42394] = 25'b10100101_10011000_00111101_1;
      patterns[42395] = 25'b10100101_10011001_00111110_1;
      patterns[42396] = 25'b10100101_10011010_00111111_1;
      patterns[42397] = 25'b10100101_10011011_01000000_1;
      patterns[42398] = 25'b10100101_10011100_01000001_1;
      patterns[42399] = 25'b10100101_10011101_01000010_1;
      patterns[42400] = 25'b10100101_10011110_01000011_1;
      patterns[42401] = 25'b10100101_10011111_01000100_1;
      patterns[42402] = 25'b10100101_10100000_01000101_1;
      patterns[42403] = 25'b10100101_10100001_01000110_1;
      patterns[42404] = 25'b10100101_10100010_01000111_1;
      patterns[42405] = 25'b10100101_10100011_01001000_1;
      patterns[42406] = 25'b10100101_10100100_01001001_1;
      patterns[42407] = 25'b10100101_10100101_01001010_1;
      patterns[42408] = 25'b10100101_10100110_01001011_1;
      patterns[42409] = 25'b10100101_10100111_01001100_1;
      patterns[42410] = 25'b10100101_10101000_01001101_1;
      patterns[42411] = 25'b10100101_10101001_01001110_1;
      patterns[42412] = 25'b10100101_10101010_01001111_1;
      patterns[42413] = 25'b10100101_10101011_01010000_1;
      patterns[42414] = 25'b10100101_10101100_01010001_1;
      patterns[42415] = 25'b10100101_10101101_01010010_1;
      patterns[42416] = 25'b10100101_10101110_01010011_1;
      patterns[42417] = 25'b10100101_10101111_01010100_1;
      patterns[42418] = 25'b10100101_10110000_01010101_1;
      patterns[42419] = 25'b10100101_10110001_01010110_1;
      patterns[42420] = 25'b10100101_10110010_01010111_1;
      patterns[42421] = 25'b10100101_10110011_01011000_1;
      patterns[42422] = 25'b10100101_10110100_01011001_1;
      patterns[42423] = 25'b10100101_10110101_01011010_1;
      patterns[42424] = 25'b10100101_10110110_01011011_1;
      patterns[42425] = 25'b10100101_10110111_01011100_1;
      patterns[42426] = 25'b10100101_10111000_01011101_1;
      patterns[42427] = 25'b10100101_10111001_01011110_1;
      patterns[42428] = 25'b10100101_10111010_01011111_1;
      patterns[42429] = 25'b10100101_10111011_01100000_1;
      patterns[42430] = 25'b10100101_10111100_01100001_1;
      patterns[42431] = 25'b10100101_10111101_01100010_1;
      patterns[42432] = 25'b10100101_10111110_01100011_1;
      patterns[42433] = 25'b10100101_10111111_01100100_1;
      patterns[42434] = 25'b10100101_11000000_01100101_1;
      patterns[42435] = 25'b10100101_11000001_01100110_1;
      patterns[42436] = 25'b10100101_11000010_01100111_1;
      patterns[42437] = 25'b10100101_11000011_01101000_1;
      patterns[42438] = 25'b10100101_11000100_01101001_1;
      patterns[42439] = 25'b10100101_11000101_01101010_1;
      patterns[42440] = 25'b10100101_11000110_01101011_1;
      patterns[42441] = 25'b10100101_11000111_01101100_1;
      patterns[42442] = 25'b10100101_11001000_01101101_1;
      patterns[42443] = 25'b10100101_11001001_01101110_1;
      patterns[42444] = 25'b10100101_11001010_01101111_1;
      patterns[42445] = 25'b10100101_11001011_01110000_1;
      patterns[42446] = 25'b10100101_11001100_01110001_1;
      patterns[42447] = 25'b10100101_11001101_01110010_1;
      patterns[42448] = 25'b10100101_11001110_01110011_1;
      patterns[42449] = 25'b10100101_11001111_01110100_1;
      patterns[42450] = 25'b10100101_11010000_01110101_1;
      patterns[42451] = 25'b10100101_11010001_01110110_1;
      patterns[42452] = 25'b10100101_11010010_01110111_1;
      patterns[42453] = 25'b10100101_11010011_01111000_1;
      patterns[42454] = 25'b10100101_11010100_01111001_1;
      patterns[42455] = 25'b10100101_11010101_01111010_1;
      patterns[42456] = 25'b10100101_11010110_01111011_1;
      patterns[42457] = 25'b10100101_11010111_01111100_1;
      patterns[42458] = 25'b10100101_11011000_01111101_1;
      patterns[42459] = 25'b10100101_11011001_01111110_1;
      patterns[42460] = 25'b10100101_11011010_01111111_1;
      patterns[42461] = 25'b10100101_11011011_10000000_1;
      patterns[42462] = 25'b10100101_11011100_10000001_1;
      patterns[42463] = 25'b10100101_11011101_10000010_1;
      patterns[42464] = 25'b10100101_11011110_10000011_1;
      patterns[42465] = 25'b10100101_11011111_10000100_1;
      patterns[42466] = 25'b10100101_11100000_10000101_1;
      patterns[42467] = 25'b10100101_11100001_10000110_1;
      patterns[42468] = 25'b10100101_11100010_10000111_1;
      patterns[42469] = 25'b10100101_11100011_10001000_1;
      patterns[42470] = 25'b10100101_11100100_10001001_1;
      patterns[42471] = 25'b10100101_11100101_10001010_1;
      patterns[42472] = 25'b10100101_11100110_10001011_1;
      patterns[42473] = 25'b10100101_11100111_10001100_1;
      patterns[42474] = 25'b10100101_11101000_10001101_1;
      patterns[42475] = 25'b10100101_11101001_10001110_1;
      patterns[42476] = 25'b10100101_11101010_10001111_1;
      patterns[42477] = 25'b10100101_11101011_10010000_1;
      patterns[42478] = 25'b10100101_11101100_10010001_1;
      patterns[42479] = 25'b10100101_11101101_10010010_1;
      patterns[42480] = 25'b10100101_11101110_10010011_1;
      patterns[42481] = 25'b10100101_11101111_10010100_1;
      patterns[42482] = 25'b10100101_11110000_10010101_1;
      patterns[42483] = 25'b10100101_11110001_10010110_1;
      patterns[42484] = 25'b10100101_11110010_10010111_1;
      patterns[42485] = 25'b10100101_11110011_10011000_1;
      patterns[42486] = 25'b10100101_11110100_10011001_1;
      patterns[42487] = 25'b10100101_11110101_10011010_1;
      patterns[42488] = 25'b10100101_11110110_10011011_1;
      patterns[42489] = 25'b10100101_11110111_10011100_1;
      patterns[42490] = 25'b10100101_11111000_10011101_1;
      patterns[42491] = 25'b10100101_11111001_10011110_1;
      patterns[42492] = 25'b10100101_11111010_10011111_1;
      patterns[42493] = 25'b10100101_11111011_10100000_1;
      patterns[42494] = 25'b10100101_11111100_10100001_1;
      patterns[42495] = 25'b10100101_11111101_10100010_1;
      patterns[42496] = 25'b10100101_11111110_10100011_1;
      patterns[42497] = 25'b10100101_11111111_10100100_1;
      patterns[42498] = 25'b10100110_00000000_10100110_0;
      patterns[42499] = 25'b10100110_00000001_10100111_0;
      patterns[42500] = 25'b10100110_00000010_10101000_0;
      patterns[42501] = 25'b10100110_00000011_10101001_0;
      patterns[42502] = 25'b10100110_00000100_10101010_0;
      patterns[42503] = 25'b10100110_00000101_10101011_0;
      patterns[42504] = 25'b10100110_00000110_10101100_0;
      patterns[42505] = 25'b10100110_00000111_10101101_0;
      patterns[42506] = 25'b10100110_00001000_10101110_0;
      patterns[42507] = 25'b10100110_00001001_10101111_0;
      patterns[42508] = 25'b10100110_00001010_10110000_0;
      patterns[42509] = 25'b10100110_00001011_10110001_0;
      patterns[42510] = 25'b10100110_00001100_10110010_0;
      patterns[42511] = 25'b10100110_00001101_10110011_0;
      patterns[42512] = 25'b10100110_00001110_10110100_0;
      patterns[42513] = 25'b10100110_00001111_10110101_0;
      patterns[42514] = 25'b10100110_00010000_10110110_0;
      patterns[42515] = 25'b10100110_00010001_10110111_0;
      patterns[42516] = 25'b10100110_00010010_10111000_0;
      patterns[42517] = 25'b10100110_00010011_10111001_0;
      patterns[42518] = 25'b10100110_00010100_10111010_0;
      patterns[42519] = 25'b10100110_00010101_10111011_0;
      patterns[42520] = 25'b10100110_00010110_10111100_0;
      patterns[42521] = 25'b10100110_00010111_10111101_0;
      patterns[42522] = 25'b10100110_00011000_10111110_0;
      patterns[42523] = 25'b10100110_00011001_10111111_0;
      patterns[42524] = 25'b10100110_00011010_11000000_0;
      patterns[42525] = 25'b10100110_00011011_11000001_0;
      patterns[42526] = 25'b10100110_00011100_11000010_0;
      patterns[42527] = 25'b10100110_00011101_11000011_0;
      patterns[42528] = 25'b10100110_00011110_11000100_0;
      patterns[42529] = 25'b10100110_00011111_11000101_0;
      patterns[42530] = 25'b10100110_00100000_11000110_0;
      patterns[42531] = 25'b10100110_00100001_11000111_0;
      patterns[42532] = 25'b10100110_00100010_11001000_0;
      patterns[42533] = 25'b10100110_00100011_11001001_0;
      patterns[42534] = 25'b10100110_00100100_11001010_0;
      patterns[42535] = 25'b10100110_00100101_11001011_0;
      patterns[42536] = 25'b10100110_00100110_11001100_0;
      patterns[42537] = 25'b10100110_00100111_11001101_0;
      patterns[42538] = 25'b10100110_00101000_11001110_0;
      patterns[42539] = 25'b10100110_00101001_11001111_0;
      patterns[42540] = 25'b10100110_00101010_11010000_0;
      patterns[42541] = 25'b10100110_00101011_11010001_0;
      patterns[42542] = 25'b10100110_00101100_11010010_0;
      patterns[42543] = 25'b10100110_00101101_11010011_0;
      patterns[42544] = 25'b10100110_00101110_11010100_0;
      patterns[42545] = 25'b10100110_00101111_11010101_0;
      patterns[42546] = 25'b10100110_00110000_11010110_0;
      patterns[42547] = 25'b10100110_00110001_11010111_0;
      patterns[42548] = 25'b10100110_00110010_11011000_0;
      patterns[42549] = 25'b10100110_00110011_11011001_0;
      patterns[42550] = 25'b10100110_00110100_11011010_0;
      patterns[42551] = 25'b10100110_00110101_11011011_0;
      patterns[42552] = 25'b10100110_00110110_11011100_0;
      patterns[42553] = 25'b10100110_00110111_11011101_0;
      patterns[42554] = 25'b10100110_00111000_11011110_0;
      patterns[42555] = 25'b10100110_00111001_11011111_0;
      patterns[42556] = 25'b10100110_00111010_11100000_0;
      patterns[42557] = 25'b10100110_00111011_11100001_0;
      patterns[42558] = 25'b10100110_00111100_11100010_0;
      patterns[42559] = 25'b10100110_00111101_11100011_0;
      patterns[42560] = 25'b10100110_00111110_11100100_0;
      patterns[42561] = 25'b10100110_00111111_11100101_0;
      patterns[42562] = 25'b10100110_01000000_11100110_0;
      patterns[42563] = 25'b10100110_01000001_11100111_0;
      patterns[42564] = 25'b10100110_01000010_11101000_0;
      patterns[42565] = 25'b10100110_01000011_11101001_0;
      patterns[42566] = 25'b10100110_01000100_11101010_0;
      patterns[42567] = 25'b10100110_01000101_11101011_0;
      patterns[42568] = 25'b10100110_01000110_11101100_0;
      patterns[42569] = 25'b10100110_01000111_11101101_0;
      patterns[42570] = 25'b10100110_01001000_11101110_0;
      patterns[42571] = 25'b10100110_01001001_11101111_0;
      patterns[42572] = 25'b10100110_01001010_11110000_0;
      patterns[42573] = 25'b10100110_01001011_11110001_0;
      patterns[42574] = 25'b10100110_01001100_11110010_0;
      patterns[42575] = 25'b10100110_01001101_11110011_0;
      patterns[42576] = 25'b10100110_01001110_11110100_0;
      patterns[42577] = 25'b10100110_01001111_11110101_0;
      patterns[42578] = 25'b10100110_01010000_11110110_0;
      patterns[42579] = 25'b10100110_01010001_11110111_0;
      patterns[42580] = 25'b10100110_01010010_11111000_0;
      patterns[42581] = 25'b10100110_01010011_11111001_0;
      patterns[42582] = 25'b10100110_01010100_11111010_0;
      patterns[42583] = 25'b10100110_01010101_11111011_0;
      patterns[42584] = 25'b10100110_01010110_11111100_0;
      patterns[42585] = 25'b10100110_01010111_11111101_0;
      patterns[42586] = 25'b10100110_01011000_11111110_0;
      patterns[42587] = 25'b10100110_01011001_11111111_0;
      patterns[42588] = 25'b10100110_01011010_00000000_1;
      patterns[42589] = 25'b10100110_01011011_00000001_1;
      patterns[42590] = 25'b10100110_01011100_00000010_1;
      patterns[42591] = 25'b10100110_01011101_00000011_1;
      patterns[42592] = 25'b10100110_01011110_00000100_1;
      patterns[42593] = 25'b10100110_01011111_00000101_1;
      patterns[42594] = 25'b10100110_01100000_00000110_1;
      patterns[42595] = 25'b10100110_01100001_00000111_1;
      patterns[42596] = 25'b10100110_01100010_00001000_1;
      patterns[42597] = 25'b10100110_01100011_00001001_1;
      patterns[42598] = 25'b10100110_01100100_00001010_1;
      patterns[42599] = 25'b10100110_01100101_00001011_1;
      patterns[42600] = 25'b10100110_01100110_00001100_1;
      patterns[42601] = 25'b10100110_01100111_00001101_1;
      patterns[42602] = 25'b10100110_01101000_00001110_1;
      patterns[42603] = 25'b10100110_01101001_00001111_1;
      patterns[42604] = 25'b10100110_01101010_00010000_1;
      patterns[42605] = 25'b10100110_01101011_00010001_1;
      patterns[42606] = 25'b10100110_01101100_00010010_1;
      patterns[42607] = 25'b10100110_01101101_00010011_1;
      patterns[42608] = 25'b10100110_01101110_00010100_1;
      patterns[42609] = 25'b10100110_01101111_00010101_1;
      patterns[42610] = 25'b10100110_01110000_00010110_1;
      patterns[42611] = 25'b10100110_01110001_00010111_1;
      patterns[42612] = 25'b10100110_01110010_00011000_1;
      patterns[42613] = 25'b10100110_01110011_00011001_1;
      patterns[42614] = 25'b10100110_01110100_00011010_1;
      patterns[42615] = 25'b10100110_01110101_00011011_1;
      patterns[42616] = 25'b10100110_01110110_00011100_1;
      patterns[42617] = 25'b10100110_01110111_00011101_1;
      patterns[42618] = 25'b10100110_01111000_00011110_1;
      patterns[42619] = 25'b10100110_01111001_00011111_1;
      patterns[42620] = 25'b10100110_01111010_00100000_1;
      patterns[42621] = 25'b10100110_01111011_00100001_1;
      patterns[42622] = 25'b10100110_01111100_00100010_1;
      patterns[42623] = 25'b10100110_01111101_00100011_1;
      patterns[42624] = 25'b10100110_01111110_00100100_1;
      patterns[42625] = 25'b10100110_01111111_00100101_1;
      patterns[42626] = 25'b10100110_10000000_00100110_1;
      patterns[42627] = 25'b10100110_10000001_00100111_1;
      patterns[42628] = 25'b10100110_10000010_00101000_1;
      patterns[42629] = 25'b10100110_10000011_00101001_1;
      patterns[42630] = 25'b10100110_10000100_00101010_1;
      patterns[42631] = 25'b10100110_10000101_00101011_1;
      patterns[42632] = 25'b10100110_10000110_00101100_1;
      patterns[42633] = 25'b10100110_10000111_00101101_1;
      patterns[42634] = 25'b10100110_10001000_00101110_1;
      patterns[42635] = 25'b10100110_10001001_00101111_1;
      patterns[42636] = 25'b10100110_10001010_00110000_1;
      patterns[42637] = 25'b10100110_10001011_00110001_1;
      patterns[42638] = 25'b10100110_10001100_00110010_1;
      patterns[42639] = 25'b10100110_10001101_00110011_1;
      patterns[42640] = 25'b10100110_10001110_00110100_1;
      patterns[42641] = 25'b10100110_10001111_00110101_1;
      patterns[42642] = 25'b10100110_10010000_00110110_1;
      patterns[42643] = 25'b10100110_10010001_00110111_1;
      patterns[42644] = 25'b10100110_10010010_00111000_1;
      patterns[42645] = 25'b10100110_10010011_00111001_1;
      patterns[42646] = 25'b10100110_10010100_00111010_1;
      patterns[42647] = 25'b10100110_10010101_00111011_1;
      patterns[42648] = 25'b10100110_10010110_00111100_1;
      patterns[42649] = 25'b10100110_10010111_00111101_1;
      patterns[42650] = 25'b10100110_10011000_00111110_1;
      patterns[42651] = 25'b10100110_10011001_00111111_1;
      patterns[42652] = 25'b10100110_10011010_01000000_1;
      patterns[42653] = 25'b10100110_10011011_01000001_1;
      patterns[42654] = 25'b10100110_10011100_01000010_1;
      patterns[42655] = 25'b10100110_10011101_01000011_1;
      patterns[42656] = 25'b10100110_10011110_01000100_1;
      patterns[42657] = 25'b10100110_10011111_01000101_1;
      patterns[42658] = 25'b10100110_10100000_01000110_1;
      patterns[42659] = 25'b10100110_10100001_01000111_1;
      patterns[42660] = 25'b10100110_10100010_01001000_1;
      patterns[42661] = 25'b10100110_10100011_01001001_1;
      patterns[42662] = 25'b10100110_10100100_01001010_1;
      patterns[42663] = 25'b10100110_10100101_01001011_1;
      patterns[42664] = 25'b10100110_10100110_01001100_1;
      patterns[42665] = 25'b10100110_10100111_01001101_1;
      patterns[42666] = 25'b10100110_10101000_01001110_1;
      patterns[42667] = 25'b10100110_10101001_01001111_1;
      patterns[42668] = 25'b10100110_10101010_01010000_1;
      patterns[42669] = 25'b10100110_10101011_01010001_1;
      patterns[42670] = 25'b10100110_10101100_01010010_1;
      patterns[42671] = 25'b10100110_10101101_01010011_1;
      patterns[42672] = 25'b10100110_10101110_01010100_1;
      patterns[42673] = 25'b10100110_10101111_01010101_1;
      patterns[42674] = 25'b10100110_10110000_01010110_1;
      patterns[42675] = 25'b10100110_10110001_01010111_1;
      patterns[42676] = 25'b10100110_10110010_01011000_1;
      patterns[42677] = 25'b10100110_10110011_01011001_1;
      patterns[42678] = 25'b10100110_10110100_01011010_1;
      patterns[42679] = 25'b10100110_10110101_01011011_1;
      patterns[42680] = 25'b10100110_10110110_01011100_1;
      patterns[42681] = 25'b10100110_10110111_01011101_1;
      patterns[42682] = 25'b10100110_10111000_01011110_1;
      patterns[42683] = 25'b10100110_10111001_01011111_1;
      patterns[42684] = 25'b10100110_10111010_01100000_1;
      patterns[42685] = 25'b10100110_10111011_01100001_1;
      patterns[42686] = 25'b10100110_10111100_01100010_1;
      patterns[42687] = 25'b10100110_10111101_01100011_1;
      patterns[42688] = 25'b10100110_10111110_01100100_1;
      patterns[42689] = 25'b10100110_10111111_01100101_1;
      patterns[42690] = 25'b10100110_11000000_01100110_1;
      patterns[42691] = 25'b10100110_11000001_01100111_1;
      patterns[42692] = 25'b10100110_11000010_01101000_1;
      patterns[42693] = 25'b10100110_11000011_01101001_1;
      patterns[42694] = 25'b10100110_11000100_01101010_1;
      patterns[42695] = 25'b10100110_11000101_01101011_1;
      patterns[42696] = 25'b10100110_11000110_01101100_1;
      patterns[42697] = 25'b10100110_11000111_01101101_1;
      patterns[42698] = 25'b10100110_11001000_01101110_1;
      patterns[42699] = 25'b10100110_11001001_01101111_1;
      patterns[42700] = 25'b10100110_11001010_01110000_1;
      patterns[42701] = 25'b10100110_11001011_01110001_1;
      patterns[42702] = 25'b10100110_11001100_01110010_1;
      patterns[42703] = 25'b10100110_11001101_01110011_1;
      patterns[42704] = 25'b10100110_11001110_01110100_1;
      patterns[42705] = 25'b10100110_11001111_01110101_1;
      patterns[42706] = 25'b10100110_11010000_01110110_1;
      patterns[42707] = 25'b10100110_11010001_01110111_1;
      patterns[42708] = 25'b10100110_11010010_01111000_1;
      patterns[42709] = 25'b10100110_11010011_01111001_1;
      patterns[42710] = 25'b10100110_11010100_01111010_1;
      patterns[42711] = 25'b10100110_11010101_01111011_1;
      patterns[42712] = 25'b10100110_11010110_01111100_1;
      patterns[42713] = 25'b10100110_11010111_01111101_1;
      patterns[42714] = 25'b10100110_11011000_01111110_1;
      patterns[42715] = 25'b10100110_11011001_01111111_1;
      patterns[42716] = 25'b10100110_11011010_10000000_1;
      patterns[42717] = 25'b10100110_11011011_10000001_1;
      patterns[42718] = 25'b10100110_11011100_10000010_1;
      patterns[42719] = 25'b10100110_11011101_10000011_1;
      patterns[42720] = 25'b10100110_11011110_10000100_1;
      patterns[42721] = 25'b10100110_11011111_10000101_1;
      patterns[42722] = 25'b10100110_11100000_10000110_1;
      patterns[42723] = 25'b10100110_11100001_10000111_1;
      patterns[42724] = 25'b10100110_11100010_10001000_1;
      patterns[42725] = 25'b10100110_11100011_10001001_1;
      patterns[42726] = 25'b10100110_11100100_10001010_1;
      patterns[42727] = 25'b10100110_11100101_10001011_1;
      patterns[42728] = 25'b10100110_11100110_10001100_1;
      patterns[42729] = 25'b10100110_11100111_10001101_1;
      patterns[42730] = 25'b10100110_11101000_10001110_1;
      patterns[42731] = 25'b10100110_11101001_10001111_1;
      patterns[42732] = 25'b10100110_11101010_10010000_1;
      patterns[42733] = 25'b10100110_11101011_10010001_1;
      patterns[42734] = 25'b10100110_11101100_10010010_1;
      patterns[42735] = 25'b10100110_11101101_10010011_1;
      patterns[42736] = 25'b10100110_11101110_10010100_1;
      patterns[42737] = 25'b10100110_11101111_10010101_1;
      patterns[42738] = 25'b10100110_11110000_10010110_1;
      patterns[42739] = 25'b10100110_11110001_10010111_1;
      patterns[42740] = 25'b10100110_11110010_10011000_1;
      patterns[42741] = 25'b10100110_11110011_10011001_1;
      patterns[42742] = 25'b10100110_11110100_10011010_1;
      patterns[42743] = 25'b10100110_11110101_10011011_1;
      patterns[42744] = 25'b10100110_11110110_10011100_1;
      patterns[42745] = 25'b10100110_11110111_10011101_1;
      patterns[42746] = 25'b10100110_11111000_10011110_1;
      patterns[42747] = 25'b10100110_11111001_10011111_1;
      patterns[42748] = 25'b10100110_11111010_10100000_1;
      patterns[42749] = 25'b10100110_11111011_10100001_1;
      patterns[42750] = 25'b10100110_11111100_10100010_1;
      patterns[42751] = 25'b10100110_11111101_10100011_1;
      patterns[42752] = 25'b10100110_11111110_10100100_1;
      patterns[42753] = 25'b10100110_11111111_10100101_1;
      patterns[42754] = 25'b10100111_00000000_10100111_0;
      patterns[42755] = 25'b10100111_00000001_10101000_0;
      patterns[42756] = 25'b10100111_00000010_10101001_0;
      patterns[42757] = 25'b10100111_00000011_10101010_0;
      patterns[42758] = 25'b10100111_00000100_10101011_0;
      patterns[42759] = 25'b10100111_00000101_10101100_0;
      patterns[42760] = 25'b10100111_00000110_10101101_0;
      patterns[42761] = 25'b10100111_00000111_10101110_0;
      patterns[42762] = 25'b10100111_00001000_10101111_0;
      patterns[42763] = 25'b10100111_00001001_10110000_0;
      patterns[42764] = 25'b10100111_00001010_10110001_0;
      patterns[42765] = 25'b10100111_00001011_10110010_0;
      patterns[42766] = 25'b10100111_00001100_10110011_0;
      patterns[42767] = 25'b10100111_00001101_10110100_0;
      patterns[42768] = 25'b10100111_00001110_10110101_0;
      patterns[42769] = 25'b10100111_00001111_10110110_0;
      patterns[42770] = 25'b10100111_00010000_10110111_0;
      patterns[42771] = 25'b10100111_00010001_10111000_0;
      patterns[42772] = 25'b10100111_00010010_10111001_0;
      patterns[42773] = 25'b10100111_00010011_10111010_0;
      patterns[42774] = 25'b10100111_00010100_10111011_0;
      patterns[42775] = 25'b10100111_00010101_10111100_0;
      patterns[42776] = 25'b10100111_00010110_10111101_0;
      patterns[42777] = 25'b10100111_00010111_10111110_0;
      patterns[42778] = 25'b10100111_00011000_10111111_0;
      patterns[42779] = 25'b10100111_00011001_11000000_0;
      patterns[42780] = 25'b10100111_00011010_11000001_0;
      patterns[42781] = 25'b10100111_00011011_11000010_0;
      patterns[42782] = 25'b10100111_00011100_11000011_0;
      patterns[42783] = 25'b10100111_00011101_11000100_0;
      patterns[42784] = 25'b10100111_00011110_11000101_0;
      patterns[42785] = 25'b10100111_00011111_11000110_0;
      patterns[42786] = 25'b10100111_00100000_11000111_0;
      patterns[42787] = 25'b10100111_00100001_11001000_0;
      patterns[42788] = 25'b10100111_00100010_11001001_0;
      patterns[42789] = 25'b10100111_00100011_11001010_0;
      patterns[42790] = 25'b10100111_00100100_11001011_0;
      patterns[42791] = 25'b10100111_00100101_11001100_0;
      patterns[42792] = 25'b10100111_00100110_11001101_0;
      patterns[42793] = 25'b10100111_00100111_11001110_0;
      patterns[42794] = 25'b10100111_00101000_11001111_0;
      patterns[42795] = 25'b10100111_00101001_11010000_0;
      patterns[42796] = 25'b10100111_00101010_11010001_0;
      patterns[42797] = 25'b10100111_00101011_11010010_0;
      patterns[42798] = 25'b10100111_00101100_11010011_0;
      patterns[42799] = 25'b10100111_00101101_11010100_0;
      patterns[42800] = 25'b10100111_00101110_11010101_0;
      patterns[42801] = 25'b10100111_00101111_11010110_0;
      patterns[42802] = 25'b10100111_00110000_11010111_0;
      patterns[42803] = 25'b10100111_00110001_11011000_0;
      patterns[42804] = 25'b10100111_00110010_11011001_0;
      patterns[42805] = 25'b10100111_00110011_11011010_0;
      patterns[42806] = 25'b10100111_00110100_11011011_0;
      patterns[42807] = 25'b10100111_00110101_11011100_0;
      patterns[42808] = 25'b10100111_00110110_11011101_0;
      patterns[42809] = 25'b10100111_00110111_11011110_0;
      patterns[42810] = 25'b10100111_00111000_11011111_0;
      patterns[42811] = 25'b10100111_00111001_11100000_0;
      patterns[42812] = 25'b10100111_00111010_11100001_0;
      patterns[42813] = 25'b10100111_00111011_11100010_0;
      patterns[42814] = 25'b10100111_00111100_11100011_0;
      patterns[42815] = 25'b10100111_00111101_11100100_0;
      patterns[42816] = 25'b10100111_00111110_11100101_0;
      patterns[42817] = 25'b10100111_00111111_11100110_0;
      patterns[42818] = 25'b10100111_01000000_11100111_0;
      patterns[42819] = 25'b10100111_01000001_11101000_0;
      patterns[42820] = 25'b10100111_01000010_11101001_0;
      patterns[42821] = 25'b10100111_01000011_11101010_0;
      patterns[42822] = 25'b10100111_01000100_11101011_0;
      patterns[42823] = 25'b10100111_01000101_11101100_0;
      patterns[42824] = 25'b10100111_01000110_11101101_0;
      patterns[42825] = 25'b10100111_01000111_11101110_0;
      patterns[42826] = 25'b10100111_01001000_11101111_0;
      patterns[42827] = 25'b10100111_01001001_11110000_0;
      patterns[42828] = 25'b10100111_01001010_11110001_0;
      patterns[42829] = 25'b10100111_01001011_11110010_0;
      patterns[42830] = 25'b10100111_01001100_11110011_0;
      patterns[42831] = 25'b10100111_01001101_11110100_0;
      patterns[42832] = 25'b10100111_01001110_11110101_0;
      patterns[42833] = 25'b10100111_01001111_11110110_0;
      patterns[42834] = 25'b10100111_01010000_11110111_0;
      patterns[42835] = 25'b10100111_01010001_11111000_0;
      patterns[42836] = 25'b10100111_01010010_11111001_0;
      patterns[42837] = 25'b10100111_01010011_11111010_0;
      patterns[42838] = 25'b10100111_01010100_11111011_0;
      patterns[42839] = 25'b10100111_01010101_11111100_0;
      patterns[42840] = 25'b10100111_01010110_11111101_0;
      patterns[42841] = 25'b10100111_01010111_11111110_0;
      patterns[42842] = 25'b10100111_01011000_11111111_0;
      patterns[42843] = 25'b10100111_01011001_00000000_1;
      patterns[42844] = 25'b10100111_01011010_00000001_1;
      patterns[42845] = 25'b10100111_01011011_00000010_1;
      patterns[42846] = 25'b10100111_01011100_00000011_1;
      patterns[42847] = 25'b10100111_01011101_00000100_1;
      patterns[42848] = 25'b10100111_01011110_00000101_1;
      patterns[42849] = 25'b10100111_01011111_00000110_1;
      patterns[42850] = 25'b10100111_01100000_00000111_1;
      patterns[42851] = 25'b10100111_01100001_00001000_1;
      patterns[42852] = 25'b10100111_01100010_00001001_1;
      patterns[42853] = 25'b10100111_01100011_00001010_1;
      patterns[42854] = 25'b10100111_01100100_00001011_1;
      patterns[42855] = 25'b10100111_01100101_00001100_1;
      patterns[42856] = 25'b10100111_01100110_00001101_1;
      patterns[42857] = 25'b10100111_01100111_00001110_1;
      patterns[42858] = 25'b10100111_01101000_00001111_1;
      patterns[42859] = 25'b10100111_01101001_00010000_1;
      patterns[42860] = 25'b10100111_01101010_00010001_1;
      patterns[42861] = 25'b10100111_01101011_00010010_1;
      patterns[42862] = 25'b10100111_01101100_00010011_1;
      patterns[42863] = 25'b10100111_01101101_00010100_1;
      patterns[42864] = 25'b10100111_01101110_00010101_1;
      patterns[42865] = 25'b10100111_01101111_00010110_1;
      patterns[42866] = 25'b10100111_01110000_00010111_1;
      patterns[42867] = 25'b10100111_01110001_00011000_1;
      patterns[42868] = 25'b10100111_01110010_00011001_1;
      patterns[42869] = 25'b10100111_01110011_00011010_1;
      patterns[42870] = 25'b10100111_01110100_00011011_1;
      patterns[42871] = 25'b10100111_01110101_00011100_1;
      patterns[42872] = 25'b10100111_01110110_00011101_1;
      patterns[42873] = 25'b10100111_01110111_00011110_1;
      patterns[42874] = 25'b10100111_01111000_00011111_1;
      patterns[42875] = 25'b10100111_01111001_00100000_1;
      patterns[42876] = 25'b10100111_01111010_00100001_1;
      patterns[42877] = 25'b10100111_01111011_00100010_1;
      patterns[42878] = 25'b10100111_01111100_00100011_1;
      patterns[42879] = 25'b10100111_01111101_00100100_1;
      patterns[42880] = 25'b10100111_01111110_00100101_1;
      patterns[42881] = 25'b10100111_01111111_00100110_1;
      patterns[42882] = 25'b10100111_10000000_00100111_1;
      patterns[42883] = 25'b10100111_10000001_00101000_1;
      patterns[42884] = 25'b10100111_10000010_00101001_1;
      patterns[42885] = 25'b10100111_10000011_00101010_1;
      patterns[42886] = 25'b10100111_10000100_00101011_1;
      patterns[42887] = 25'b10100111_10000101_00101100_1;
      patterns[42888] = 25'b10100111_10000110_00101101_1;
      patterns[42889] = 25'b10100111_10000111_00101110_1;
      patterns[42890] = 25'b10100111_10001000_00101111_1;
      patterns[42891] = 25'b10100111_10001001_00110000_1;
      patterns[42892] = 25'b10100111_10001010_00110001_1;
      patterns[42893] = 25'b10100111_10001011_00110010_1;
      patterns[42894] = 25'b10100111_10001100_00110011_1;
      patterns[42895] = 25'b10100111_10001101_00110100_1;
      patterns[42896] = 25'b10100111_10001110_00110101_1;
      patterns[42897] = 25'b10100111_10001111_00110110_1;
      patterns[42898] = 25'b10100111_10010000_00110111_1;
      patterns[42899] = 25'b10100111_10010001_00111000_1;
      patterns[42900] = 25'b10100111_10010010_00111001_1;
      patterns[42901] = 25'b10100111_10010011_00111010_1;
      patterns[42902] = 25'b10100111_10010100_00111011_1;
      patterns[42903] = 25'b10100111_10010101_00111100_1;
      patterns[42904] = 25'b10100111_10010110_00111101_1;
      patterns[42905] = 25'b10100111_10010111_00111110_1;
      patterns[42906] = 25'b10100111_10011000_00111111_1;
      patterns[42907] = 25'b10100111_10011001_01000000_1;
      patterns[42908] = 25'b10100111_10011010_01000001_1;
      patterns[42909] = 25'b10100111_10011011_01000010_1;
      patterns[42910] = 25'b10100111_10011100_01000011_1;
      patterns[42911] = 25'b10100111_10011101_01000100_1;
      patterns[42912] = 25'b10100111_10011110_01000101_1;
      patterns[42913] = 25'b10100111_10011111_01000110_1;
      patterns[42914] = 25'b10100111_10100000_01000111_1;
      patterns[42915] = 25'b10100111_10100001_01001000_1;
      patterns[42916] = 25'b10100111_10100010_01001001_1;
      patterns[42917] = 25'b10100111_10100011_01001010_1;
      patterns[42918] = 25'b10100111_10100100_01001011_1;
      patterns[42919] = 25'b10100111_10100101_01001100_1;
      patterns[42920] = 25'b10100111_10100110_01001101_1;
      patterns[42921] = 25'b10100111_10100111_01001110_1;
      patterns[42922] = 25'b10100111_10101000_01001111_1;
      patterns[42923] = 25'b10100111_10101001_01010000_1;
      patterns[42924] = 25'b10100111_10101010_01010001_1;
      patterns[42925] = 25'b10100111_10101011_01010010_1;
      patterns[42926] = 25'b10100111_10101100_01010011_1;
      patterns[42927] = 25'b10100111_10101101_01010100_1;
      patterns[42928] = 25'b10100111_10101110_01010101_1;
      patterns[42929] = 25'b10100111_10101111_01010110_1;
      patterns[42930] = 25'b10100111_10110000_01010111_1;
      patterns[42931] = 25'b10100111_10110001_01011000_1;
      patterns[42932] = 25'b10100111_10110010_01011001_1;
      patterns[42933] = 25'b10100111_10110011_01011010_1;
      patterns[42934] = 25'b10100111_10110100_01011011_1;
      patterns[42935] = 25'b10100111_10110101_01011100_1;
      patterns[42936] = 25'b10100111_10110110_01011101_1;
      patterns[42937] = 25'b10100111_10110111_01011110_1;
      patterns[42938] = 25'b10100111_10111000_01011111_1;
      patterns[42939] = 25'b10100111_10111001_01100000_1;
      patterns[42940] = 25'b10100111_10111010_01100001_1;
      patterns[42941] = 25'b10100111_10111011_01100010_1;
      patterns[42942] = 25'b10100111_10111100_01100011_1;
      patterns[42943] = 25'b10100111_10111101_01100100_1;
      patterns[42944] = 25'b10100111_10111110_01100101_1;
      patterns[42945] = 25'b10100111_10111111_01100110_1;
      patterns[42946] = 25'b10100111_11000000_01100111_1;
      patterns[42947] = 25'b10100111_11000001_01101000_1;
      patterns[42948] = 25'b10100111_11000010_01101001_1;
      patterns[42949] = 25'b10100111_11000011_01101010_1;
      patterns[42950] = 25'b10100111_11000100_01101011_1;
      patterns[42951] = 25'b10100111_11000101_01101100_1;
      patterns[42952] = 25'b10100111_11000110_01101101_1;
      patterns[42953] = 25'b10100111_11000111_01101110_1;
      patterns[42954] = 25'b10100111_11001000_01101111_1;
      patterns[42955] = 25'b10100111_11001001_01110000_1;
      patterns[42956] = 25'b10100111_11001010_01110001_1;
      patterns[42957] = 25'b10100111_11001011_01110010_1;
      patterns[42958] = 25'b10100111_11001100_01110011_1;
      patterns[42959] = 25'b10100111_11001101_01110100_1;
      patterns[42960] = 25'b10100111_11001110_01110101_1;
      patterns[42961] = 25'b10100111_11001111_01110110_1;
      patterns[42962] = 25'b10100111_11010000_01110111_1;
      patterns[42963] = 25'b10100111_11010001_01111000_1;
      patterns[42964] = 25'b10100111_11010010_01111001_1;
      patterns[42965] = 25'b10100111_11010011_01111010_1;
      patterns[42966] = 25'b10100111_11010100_01111011_1;
      patterns[42967] = 25'b10100111_11010101_01111100_1;
      patterns[42968] = 25'b10100111_11010110_01111101_1;
      patterns[42969] = 25'b10100111_11010111_01111110_1;
      patterns[42970] = 25'b10100111_11011000_01111111_1;
      patterns[42971] = 25'b10100111_11011001_10000000_1;
      patterns[42972] = 25'b10100111_11011010_10000001_1;
      patterns[42973] = 25'b10100111_11011011_10000010_1;
      patterns[42974] = 25'b10100111_11011100_10000011_1;
      patterns[42975] = 25'b10100111_11011101_10000100_1;
      patterns[42976] = 25'b10100111_11011110_10000101_1;
      patterns[42977] = 25'b10100111_11011111_10000110_1;
      patterns[42978] = 25'b10100111_11100000_10000111_1;
      patterns[42979] = 25'b10100111_11100001_10001000_1;
      patterns[42980] = 25'b10100111_11100010_10001001_1;
      patterns[42981] = 25'b10100111_11100011_10001010_1;
      patterns[42982] = 25'b10100111_11100100_10001011_1;
      patterns[42983] = 25'b10100111_11100101_10001100_1;
      patterns[42984] = 25'b10100111_11100110_10001101_1;
      patterns[42985] = 25'b10100111_11100111_10001110_1;
      patterns[42986] = 25'b10100111_11101000_10001111_1;
      patterns[42987] = 25'b10100111_11101001_10010000_1;
      patterns[42988] = 25'b10100111_11101010_10010001_1;
      patterns[42989] = 25'b10100111_11101011_10010010_1;
      patterns[42990] = 25'b10100111_11101100_10010011_1;
      patterns[42991] = 25'b10100111_11101101_10010100_1;
      patterns[42992] = 25'b10100111_11101110_10010101_1;
      patterns[42993] = 25'b10100111_11101111_10010110_1;
      patterns[42994] = 25'b10100111_11110000_10010111_1;
      patterns[42995] = 25'b10100111_11110001_10011000_1;
      patterns[42996] = 25'b10100111_11110010_10011001_1;
      patterns[42997] = 25'b10100111_11110011_10011010_1;
      patterns[42998] = 25'b10100111_11110100_10011011_1;
      patterns[42999] = 25'b10100111_11110101_10011100_1;
      patterns[43000] = 25'b10100111_11110110_10011101_1;
      patterns[43001] = 25'b10100111_11110111_10011110_1;
      patterns[43002] = 25'b10100111_11111000_10011111_1;
      patterns[43003] = 25'b10100111_11111001_10100000_1;
      patterns[43004] = 25'b10100111_11111010_10100001_1;
      patterns[43005] = 25'b10100111_11111011_10100010_1;
      patterns[43006] = 25'b10100111_11111100_10100011_1;
      patterns[43007] = 25'b10100111_11111101_10100100_1;
      patterns[43008] = 25'b10100111_11111110_10100101_1;
      patterns[43009] = 25'b10100111_11111111_10100110_1;
      patterns[43010] = 25'b10101000_00000000_10101000_0;
      patterns[43011] = 25'b10101000_00000001_10101001_0;
      patterns[43012] = 25'b10101000_00000010_10101010_0;
      patterns[43013] = 25'b10101000_00000011_10101011_0;
      patterns[43014] = 25'b10101000_00000100_10101100_0;
      patterns[43015] = 25'b10101000_00000101_10101101_0;
      patterns[43016] = 25'b10101000_00000110_10101110_0;
      patterns[43017] = 25'b10101000_00000111_10101111_0;
      patterns[43018] = 25'b10101000_00001000_10110000_0;
      patterns[43019] = 25'b10101000_00001001_10110001_0;
      patterns[43020] = 25'b10101000_00001010_10110010_0;
      patterns[43021] = 25'b10101000_00001011_10110011_0;
      patterns[43022] = 25'b10101000_00001100_10110100_0;
      patterns[43023] = 25'b10101000_00001101_10110101_0;
      patterns[43024] = 25'b10101000_00001110_10110110_0;
      patterns[43025] = 25'b10101000_00001111_10110111_0;
      patterns[43026] = 25'b10101000_00010000_10111000_0;
      patterns[43027] = 25'b10101000_00010001_10111001_0;
      patterns[43028] = 25'b10101000_00010010_10111010_0;
      patterns[43029] = 25'b10101000_00010011_10111011_0;
      patterns[43030] = 25'b10101000_00010100_10111100_0;
      patterns[43031] = 25'b10101000_00010101_10111101_0;
      patterns[43032] = 25'b10101000_00010110_10111110_0;
      patterns[43033] = 25'b10101000_00010111_10111111_0;
      patterns[43034] = 25'b10101000_00011000_11000000_0;
      patterns[43035] = 25'b10101000_00011001_11000001_0;
      patterns[43036] = 25'b10101000_00011010_11000010_0;
      patterns[43037] = 25'b10101000_00011011_11000011_0;
      patterns[43038] = 25'b10101000_00011100_11000100_0;
      patterns[43039] = 25'b10101000_00011101_11000101_0;
      patterns[43040] = 25'b10101000_00011110_11000110_0;
      patterns[43041] = 25'b10101000_00011111_11000111_0;
      patterns[43042] = 25'b10101000_00100000_11001000_0;
      patterns[43043] = 25'b10101000_00100001_11001001_0;
      patterns[43044] = 25'b10101000_00100010_11001010_0;
      patterns[43045] = 25'b10101000_00100011_11001011_0;
      patterns[43046] = 25'b10101000_00100100_11001100_0;
      patterns[43047] = 25'b10101000_00100101_11001101_0;
      patterns[43048] = 25'b10101000_00100110_11001110_0;
      patterns[43049] = 25'b10101000_00100111_11001111_0;
      patterns[43050] = 25'b10101000_00101000_11010000_0;
      patterns[43051] = 25'b10101000_00101001_11010001_0;
      patterns[43052] = 25'b10101000_00101010_11010010_0;
      patterns[43053] = 25'b10101000_00101011_11010011_0;
      patterns[43054] = 25'b10101000_00101100_11010100_0;
      patterns[43055] = 25'b10101000_00101101_11010101_0;
      patterns[43056] = 25'b10101000_00101110_11010110_0;
      patterns[43057] = 25'b10101000_00101111_11010111_0;
      patterns[43058] = 25'b10101000_00110000_11011000_0;
      patterns[43059] = 25'b10101000_00110001_11011001_0;
      patterns[43060] = 25'b10101000_00110010_11011010_0;
      patterns[43061] = 25'b10101000_00110011_11011011_0;
      patterns[43062] = 25'b10101000_00110100_11011100_0;
      patterns[43063] = 25'b10101000_00110101_11011101_0;
      patterns[43064] = 25'b10101000_00110110_11011110_0;
      patterns[43065] = 25'b10101000_00110111_11011111_0;
      patterns[43066] = 25'b10101000_00111000_11100000_0;
      patterns[43067] = 25'b10101000_00111001_11100001_0;
      patterns[43068] = 25'b10101000_00111010_11100010_0;
      patterns[43069] = 25'b10101000_00111011_11100011_0;
      patterns[43070] = 25'b10101000_00111100_11100100_0;
      patterns[43071] = 25'b10101000_00111101_11100101_0;
      patterns[43072] = 25'b10101000_00111110_11100110_0;
      patterns[43073] = 25'b10101000_00111111_11100111_0;
      patterns[43074] = 25'b10101000_01000000_11101000_0;
      patterns[43075] = 25'b10101000_01000001_11101001_0;
      patterns[43076] = 25'b10101000_01000010_11101010_0;
      patterns[43077] = 25'b10101000_01000011_11101011_0;
      patterns[43078] = 25'b10101000_01000100_11101100_0;
      patterns[43079] = 25'b10101000_01000101_11101101_0;
      patterns[43080] = 25'b10101000_01000110_11101110_0;
      patterns[43081] = 25'b10101000_01000111_11101111_0;
      patterns[43082] = 25'b10101000_01001000_11110000_0;
      patterns[43083] = 25'b10101000_01001001_11110001_0;
      patterns[43084] = 25'b10101000_01001010_11110010_0;
      patterns[43085] = 25'b10101000_01001011_11110011_0;
      patterns[43086] = 25'b10101000_01001100_11110100_0;
      patterns[43087] = 25'b10101000_01001101_11110101_0;
      patterns[43088] = 25'b10101000_01001110_11110110_0;
      patterns[43089] = 25'b10101000_01001111_11110111_0;
      patterns[43090] = 25'b10101000_01010000_11111000_0;
      patterns[43091] = 25'b10101000_01010001_11111001_0;
      patterns[43092] = 25'b10101000_01010010_11111010_0;
      patterns[43093] = 25'b10101000_01010011_11111011_0;
      patterns[43094] = 25'b10101000_01010100_11111100_0;
      patterns[43095] = 25'b10101000_01010101_11111101_0;
      patterns[43096] = 25'b10101000_01010110_11111110_0;
      patterns[43097] = 25'b10101000_01010111_11111111_0;
      patterns[43098] = 25'b10101000_01011000_00000000_1;
      patterns[43099] = 25'b10101000_01011001_00000001_1;
      patterns[43100] = 25'b10101000_01011010_00000010_1;
      patterns[43101] = 25'b10101000_01011011_00000011_1;
      patterns[43102] = 25'b10101000_01011100_00000100_1;
      patterns[43103] = 25'b10101000_01011101_00000101_1;
      patterns[43104] = 25'b10101000_01011110_00000110_1;
      patterns[43105] = 25'b10101000_01011111_00000111_1;
      patterns[43106] = 25'b10101000_01100000_00001000_1;
      patterns[43107] = 25'b10101000_01100001_00001001_1;
      patterns[43108] = 25'b10101000_01100010_00001010_1;
      patterns[43109] = 25'b10101000_01100011_00001011_1;
      patterns[43110] = 25'b10101000_01100100_00001100_1;
      patterns[43111] = 25'b10101000_01100101_00001101_1;
      patterns[43112] = 25'b10101000_01100110_00001110_1;
      patterns[43113] = 25'b10101000_01100111_00001111_1;
      patterns[43114] = 25'b10101000_01101000_00010000_1;
      patterns[43115] = 25'b10101000_01101001_00010001_1;
      patterns[43116] = 25'b10101000_01101010_00010010_1;
      patterns[43117] = 25'b10101000_01101011_00010011_1;
      patterns[43118] = 25'b10101000_01101100_00010100_1;
      patterns[43119] = 25'b10101000_01101101_00010101_1;
      patterns[43120] = 25'b10101000_01101110_00010110_1;
      patterns[43121] = 25'b10101000_01101111_00010111_1;
      patterns[43122] = 25'b10101000_01110000_00011000_1;
      patterns[43123] = 25'b10101000_01110001_00011001_1;
      patterns[43124] = 25'b10101000_01110010_00011010_1;
      patterns[43125] = 25'b10101000_01110011_00011011_1;
      patterns[43126] = 25'b10101000_01110100_00011100_1;
      patterns[43127] = 25'b10101000_01110101_00011101_1;
      patterns[43128] = 25'b10101000_01110110_00011110_1;
      patterns[43129] = 25'b10101000_01110111_00011111_1;
      patterns[43130] = 25'b10101000_01111000_00100000_1;
      patterns[43131] = 25'b10101000_01111001_00100001_1;
      patterns[43132] = 25'b10101000_01111010_00100010_1;
      patterns[43133] = 25'b10101000_01111011_00100011_1;
      patterns[43134] = 25'b10101000_01111100_00100100_1;
      patterns[43135] = 25'b10101000_01111101_00100101_1;
      patterns[43136] = 25'b10101000_01111110_00100110_1;
      patterns[43137] = 25'b10101000_01111111_00100111_1;
      patterns[43138] = 25'b10101000_10000000_00101000_1;
      patterns[43139] = 25'b10101000_10000001_00101001_1;
      patterns[43140] = 25'b10101000_10000010_00101010_1;
      patterns[43141] = 25'b10101000_10000011_00101011_1;
      patterns[43142] = 25'b10101000_10000100_00101100_1;
      patterns[43143] = 25'b10101000_10000101_00101101_1;
      patterns[43144] = 25'b10101000_10000110_00101110_1;
      patterns[43145] = 25'b10101000_10000111_00101111_1;
      patterns[43146] = 25'b10101000_10001000_00110000_1;
      patterns[43147] = 25'b10101000_10001001_00110001_1;
      patterns[43148] = 25'b10101000_10001010_00110010_1;
      patterns[43149] = 25'b10101000_10001011_00110011_1;
      patterns[43150] = 25'b10101000_10001100_00110100_1;
      patterns[43151] = 25'b10101000_10001101_00110101_1;
      patterns[43152] = 25'b10101000_10001110_00110110_1;
      patterns[43153] = 25'b10101000_10001111_00110111_1;
      patterns[43154] = 25'b10101000_10010000_00111000_1;
      patterns[43155] = 25'b10101000_10010001_00111001_1;
      patterns[43156] = 25'b10101000_10010010_00111010_1;
      patterns[43157] = 25'b10101000_10010011_00111011_1;
      patterns[43158] = 25'b10101000_10010100_00111100_1;
      patterns[43159] = 25'b10101000_10010101_00111101_1;
      patterns[43160] = 25'b10101000_10010110_00111110_1;
      patterns[43161] = 25'b10101000_10010111_00111111_1;
      patterns[43162] = 25'b10101000_10011000_01000000_1;
      patterns[43163] = 25'b10101000_10011001_01000001_1;
      patterns[43164] = 25'b10101000_10011010_01000010_1;
      patterns[43165] = 25'b10101000_10011011_01000011_1;
      patterns[43166] = 25'b10101000_10011100_01000100_1;
      patterns[43167] = 25'b10101000_10011101_01000101_1;
      patterns[43168] = 25'b10101000_10011110_01000110_1;
      patterns[43169] = 25'b10101000_10011111_01000111_1;
      patterns[43170] = 25'b10101000_10100000_01001000_1;
      patterns[43171] = 25'b10101000_10100001_01001001_1;
      patterns[43172] = 25'b10101000_10100010_01001010_1;
      patterns[43173] = 25'b10101000_10100011_01001011_1;
      patterns[43174] = 25'b10101000_10100100_01001100_1;
      patterns[43175] = 25'b10101000_10100101_01001101_1;
      patterns[43176] = 25'b10101000_10100110_01001110_1;
      patterns[43177] = 25'b10101000_10100111_01001111_1;
      patterns[43178] = 25'b10101000_10101000_01010000_1;
      patterns[43179] = 25'b10101000_10101001_01010001_1;
      patterns[43180] = 25'b10101000_10101010_01010010_1;
      patterns[43181] = 25'b10101000_10101011_01010011_1;
      patterns[43182] = 25'b10101000_10101100_01010100_1;
      patterns[43183] = 25'b10101000_10101101_01010101_1;
      patterns[43184] = 25'b10101000_10101110_01010110_1;
      patterns[43185] = 25'b10101000_10101111_01010111_1;
      patterns[43186] = 25'b10101000_10110000_01011000_1;
      patterns[43187] = 25'b10101000_10110001_01011001_1;
      patterns[43188] = 25'b10101000_10110010_01011010_1;
      patterns[43189] = 25'b10101000_10110011_01011011_1;
      patterns[43190] = 25'b10101000_10110100_01011100_1;
      patterns[43191] = 25'b10101000_10110101_01011101_1;
      patterns[43192] = 25'b10101000_10110110_01011110_1;
      patterns[43193] = 25'b10101000_10110111_01011111_1;
      patterns[43194] = 25'b10101000_10111000_01100000_1;
      patterns[43195] = 25'b10101000_10111001_01100001_1;
      patterns[43196] = 25'b10101000_10111010_01100010_1;
      patterns[43197] = 25'b10101000_10111011_01100011_1;
      patterns[43198] = 25'b10101000_10111100_01100100_1;
      patterns[43199] = 25'b10101000_10111101_01100101_1;
      patterns[43200] = 25'b10101000_10111110_01100110_1;
      patterns[43201] = 25'b10101000_10111111_01100111_1;
      patterns[43202] = 25'b10101000_11000000_01101000_1;
      patterns[43203] = 25'b10101000_11000001_01101001_1;
      patterns[43204] = 25'b10101000_11000010_01101010_1;
      patterns[43205] = 25'b10101000_11000011_01101011_1;
      patterns[43206] = 25'b10101000_11000100_01101100_1;
      patterns[43207] = 25'b10101000_11000101_01101101_1;
      patterns[43208] = 25'b10101000_11000110_01101110_1;
      patterns[43209] = 25'b10101000_11000111_01101111_1;
      patterns[43210] = 25'b10101000_11001000_01110000_1;
      patterns[43211] = 25'b10101000_11001001_01110001_1;
      patterns[43212] = 25'b10101000_11001010_01110010_1;
      patterns[43213] = 25'b10101000_11001011_01110011_1;
      patterns[43214] = 25'b10101000_11001100_01110100_1;
      patterns[43215] = 25'b10101000_11001101_01110101_1;
      patterns[43216] = 25'b10101000_11001110_01110110_1;
      patterns[43217] = 25'b10101000_11001111_01110111_1;
      patterns[43218] = 25'b10101000_11010000_01111000_1;
      patterns[43219] = 25'b10101000_11010001_01111001_1;
      patterns[43220] = 25'b10101000_11010010_01111010_1;
      patterns[43221] = 25'b10101000_11010011_01111011_1;
      patterns[43222] = 25'b10101000_11010100_01111100_1;
      patterns[43223] = 25'b10101000_11010101_01111101_1;
      patterns[43224] = 25'b10101000_11010110_01111110_1;
      patterns[43225] = 25'b10101000_11010111_01111111_1;
      patterns[43226] = 25'b10101000_11011000_10000000_1;
      patterns[43227] = 25'b10101000_11011001_10000001_1;
      patterns[43228] = 25'b10101000_11011010_10000010_1;
      patterns[43229] = 25'b10101000_11011011_10000011_1;
      patterns[43230] = 25'b10101000_11011100_10000100_1;
      patterns[43231] = 25'b10101000_11011101_10000101_1;
      patterns[43232] = 25'b10101000_11011110_10000110_1;
      patterns[43233] = 25'b10101000_11011111_10000111_1;
      patterns[43234] = 25'b10101000_11100000_10001000_1;
      patterns[43235] = 25'b10101000_11100001_10001001_1;
      patterns[43236] = 25'b10101000_11100010_10001010_1;
      patterns[43237] = 25'b10101000_11100011_10001011_1;
      patterns[43238] = 25'b10101000_11100100_10001100_1;
      patterns[43239] = 25'b10101000_11100101_10001101_1;
      patterns[43240] = 25'b10101000_11100110_10001110_1;
      patterns[43241] = 25'b10101000_11100111_10001111_1;
      patterns[43242] = 25'b10101000_11101000_10010000_1;
      patterns[43243] = 25'b10101000_11101001_10010001_1;
      patterns[43244] = 25'b10101000_11101010_10010010_1;
      patterns[43245] = 25'b10101000_11101011_10010011_1;
      patterns[43246] = 25'b10101000_11101100_10010100_1;
      patterns[43247] = 25'b10101000_11101101_10010101_1;
      patterns[43248] = 25'b10101000_11101110_10010110_1;
      patterns[43249] = 25'b10101000_11101111_10010111_1;
      patterns[43250] = 25'b10101000_11110000_10011000_1;
      patterns[43251] = 25'b10101000_11110001_10011001_1;
      patterns[43252] = 25'b10101000_11110010_10011010_1;
      patterns[43253] = 25'b10101000_11110011_10011011_1;
      patterns[43254] = 25'b10101000_11110100_10011100_1;
      patterns[43255] = 25'b10101000_11110101_10011101_1;
      patterns[43256] = 25'b10101000_11110110_10011110_1;
      patterns[43257] = 25'b10101000_11110111_10011111_1;
      patterns[43258] = 25'b10101000_11111000_10100000_1;
      patterns[43259] = 25'b10101000_11111001_10100001_1;
      patterns[43260] = 25'b10101000_11111010_10100010_1;
      patterns[43261] = 25'b10101000_11111011_10100011_1;
      patterns[43262] = 25'b10101000_11111100_10100100_1;
      patterns[43263] = 25'b10101000_11111101_10100101_1;
      patterns[43264] = 25'b10101000_11111110_10100110_1;
      patterns[43265] = 25'b10101000_11111111_10100111_1;
      patterns[43266] = 25'b10101001_00000000_10101001_0;
      patterns[43267] = 25'b10101001_00000001_10101010_0;
      patterns[43268] = 25'b10101001_00000010_10101011_0;
      patterns[43269] = 25'b10101001_00000011_10101100_0;
      patterns[43270] = 25'b10101001_00000100_10101101_0;
      patterns[43271] = 25'b10101001_00000101_10101110_0;
      patterns[43272] = 25'b10101001_00000110_10101111_0;
      patterns[43273] = 25'b10101001_00000111_10110000_0;
      patterns[43274] = 25'b10101001_00001000_10110001_0;
      patterns[43275] = 25'b10101001_00001001_10110010_0;
      patterns[43276] = 25'b10101001_00001010_10110011_0;
      patterns[43277] = 25'b10101001_00001011_10110100_0;
      patterns[43278] = 25'b10101001_00001100_10110101_0;
      patterns[43279] = 25'b10101001_00001101_10110110_0;
      patterns[43280] = 25'b10101001_00001110_10110111_0;
      patterns[43281] = 25'b10101001_00001111_10111000_0;
      patterns[43282] = 25'b10101001_00010000_10111001_0;
      patterns[43283] = 25'b10101001_00010001_10111010_0;
      patterns[43284] = 25'b10101001_00010010_10111011_0;
      patterns[43285] = 25'b10101001_00010011_10111100_0;
      patterns[43286] = 25'b10101001_00010100_10111101_0;
      patterns[43287] = 25'b10101001_00010101_10111110_0;
      patterns[43288] = 25'b10101001_00010110_10111111_0;
      patterns[43289] = 25'b10101001_00010111_11000000_0;
      patterns[43290] = 25'b10101001_00011000_11000001_0;
      patterns[43291] = 25'b10101001_00011001_11000010_0;
      patterns[43292] = 25'b10101001_00011010_11000011_0;
      patterns[43293] = 25'b10101001_00011011_11000100_0;
      patterns[43294] = 25'b10101001_00011100_11000101_0;
      patterns[43295] = 25'b10101001_00011101_11000110_0;
      patterns[43296] = 25'b10101001_00011110_11000111_0;
      patterns[43297] = 25'b10101001_00011111_11001000_0;
      patterns[43298] = 25'b10101001_00100000_11001001_0;
      patterns[43299] = 25'b10101001_00100001_11001010_0;
      patterns[43300] = 25'b10101001_00100010_11001011_0;
      patterns[43301] = 25'b10101001_00100011_11001100_0;
      patterns[43302] = 25'b10101001_00100100_11001101_0;
      patterns[43303] = 25'b10101001_00100101_11001110_0;
      patterns[43304] = 25'b10101001_00100110_11001111_0;
      patterns[43305] = 25'b10101001_00100111_11010000_0;
      patterns[43306] = 25'b10101001_00101000_11010001_0;
      patterns[43307] = 25'b10101001_00101001_11010010_0;
      patterns[43308] = 25'b10101001_00101010_11010011_0;
      patterns[43309] = 25'b10101001_00101011_11010100_0;
      patterns[43310] = 25'b10101001_00101100_11010101_0;
      patterns[43311] = 25'b10101001_00101101_11010110_0;
      patterns[43312] = 25'b10101001_00101110_11010111_0;
      patterns[43313] = 25'b10101001_00101111_11011000_0;
      patterns[43314] = 25'b10101001_00110000_11011001_0;
      patterns[43315] = 25'b10101001_00110001_11011010_0;
      patterns[43316] = 25'b10101001_00110010_11011011_0;
      patterns[43317] = 25'b10101001_00110011_11011100_0;
      patterns[43318] = 25'b10101001_00110100_11011101_0;
      patterns[43319] = 25'b10101001_00110101_11011110_0;
      patterns[43320] = 25'b10101001_00110110_11011111_0;
      patterns[43321] = 25'b10101001_00110111_11100000_0;
      patterns[43322] = 25'b10101001_00111000_11100001_0;
      patterns[43323] = 25'b10101001_00111001_11100010_0;
      patterns[43324] = 25'b10101001_00111010_11100011_0;
      patterns[43325] = 25'b10101001_00111011_11100100_0;
      patterns[43326] = 25'b10101001_00111100_11100101_0;
      patterns[43327] = 25'b10101001_00111101_11100110_0;
      patterns[43328] = 25'b10101001_00111110_11100111_0;
      patterns[43329] = 25'b10101001_00111111_11101000_0;
      patterns[43330] = 25'b10101001_01000000_11101001_0;
      patterns[43331] = 25'b10101001_01000001_11101010_0;
      patterns[43332] = 25'b10101001_01000010_11101011_0;
      patterns[43333] = 25'b10101001_01000011_11101100_0;
      patterns[43334] = 25'b10101001_01000100_11101101_0;
      patterns[43335] = 25'b10101001_01000101_11101110_0;
      patterns[43336] = 25'b10101001_01000110_11101111_0;
      patterns[43337] = 25'b10101001_01000111_11110000_0;
      patterns[43338] = 25'b10101001_01001000_11110001_0;
      patterns[43339] = 25'b10101001_01001001_11110010_0;
      patterns[43340] = 25'b10101001_01001010_11110011_0;
      patterns[43341] = 25'b10101001_01001011_11110100_0;
      patterns[43342] = 25'b10101001_01001100_11110101_0;
      patterns[43343] = 25'b10101001_01001101_11110110_0;
      patterns[43344] = 25'b10101001_01001110_11110111_0;
      patterns[43345] = 25'b10101001_01001111_11111000_0;
      patterns[43346] = 25'b10101001_01010000_11111001_0;
      patterns[43347] = 25'b10101001_01010001_11111010_0;
      patterns[43348] = 25'b10101001_01010010_11111011_0;
      patterns[43349] = 25'b10101001_01010011_11111100_0;
      patterns[43350] = 25'b10101001_01010100_11111101_0;
      patterns[43351] = 25'b10101001_01010101_11111110_0;
      patterns[43352] = 25'b10101001_01010110_11111111_0;
      patterns[43353] = 25'b10101001_01010111_00000000_1;
      patterns[43354] = 25'b10101001_01011000_00000001_1;
      patterns[43355] = 25'b10101001_01011001_00000010_1;
      patterns[43356] = 25'b10101001_01011010_00000011_1;
      patterns[43357] = 25'b10101001_01011011_00000100_1;
      patterns[43358] = 25'b10101001_01011100_00000101_1;
      patterns[43359] = 25'b10101001_01011101_00000110_1;
      patterns[43360] = 25'b10101001_01011110_00000111_1;
      patterns[43361] = 25'b10101001_01011111_00001000_1;
      patterns[43362] = 25'b10101001_01100000_00001001_1;
      patterns[43363] = 25'b10101001_01100001_00001010_1;
      patterns[43364] = 25'b10101001_01100010_00001011_1;
      patterns[43365] = 25'b10101001_01100011_00001100_1;
      patterns[43366] = 25'b10101001_01100100_00001101_1;
      patterns[43367] = 25'b10101001_01100101_00001110_1;
      patterns[43368] = 25'b10101001_01100110_00001111_1;
      patterns[43369] = 25'b10101001_01100111_00010000_1;
      patterns[43370] = 25'b10101001_01101000_00010001_1;
      patterns[43371] = 25'b10101001_01101001_00010010_1;
      patterns[43372] = 25'b10101001_01101010_00010011_1;
      patterns[43373] = 25'b10101001_01101011_00010100_1;
      patterns[43374] = 25'b10101001_01101100_00010101_1;
      patterns[43375] = 25'b10101001_01101101_00010110_1;
      patterns[43376] = 25'b10101001_01101110_00010111_1;
      patterns[43377] = 25'b10101001_01101111_00011000_1;
      patterns[43378] = 25'b10101001_01110000_00011001_1;
      patterns[43379] = 25'b10101001_01110001_00011010_1;
      patterns[43380] = 25'b10101001_01110010_00011011_1;
      patterns[43381] = 25'b10101001_01110011_00011100_1;
      patterns[43382] = 25'b10101001_01110100_00011101_1;
      patterns[43383] = 25'b10101001_01110101_00011110_1;
      patterns[43384] = 25'b10101001_01110110_00011111_1;
      patterns[43385] = 25'b10101001_01110111_00100000_1;
      patterns[43386] = 25'b10101001_01111000_00100001_1;
      patterns[43387] = 25'b10101001_01111001_00100010_1;
      patterns[43388] = 25'b10101001_01111010_00100011_1;
      patterns[43389] = 25'b10101001_01111011_00100100_1;
      patterns[43390] = 25'b10101001_01111100_00100101_1;
      patterns[43391] = 25'b10101001_01111101_00100110_1;
      patterns[43392] = 25'b10101001_01111110_00100111_1;
      patterns[43393] = 25'b10101001_01111111_00101000_1;
      patterns[43394] = 25'b10101001_10000000_00101001_1;
      patterns[43395] = 25'b10101001_10000001_00101010_1;
      patterns[43396] = 25'b10101001_10000010_00101011_1;
      patterns[43397] = 25'b10101001_10000011_00101100_1;
      patterns[43398] = 25'b10101001_10000100_00101101_1;
      patterns[43399] = 25'b10101001_10000101_00101110_1;
      patterns[43400] = 25'b10101001_10000110_00101111_1;
      patterns[43401] = 25'b10101001_10000111_00110000_1;
      patterns[43402] = 25'b10101001_10001000_00110001_1;
      patterns[43403] = 25'b10101001_10001001_00110010_1;
      patterns[43404] = 25'b10101001_10001010_00110011_1;
      patterns[43405] = 25'b10101001_10001011_00110100_1;
      patterns[43406] = 25'b10101001_10001100_00110101_1;
      patterns[43407] = 25'b10101001_10001101_00110110_1;
      patterns[43408] = 25'b10101001_10001110_00110111_1;
      patterns[43409] = 25'b10101001_10001111_00111000_1;
      patterns[43410] = 25'b10101001_10010000_00111001_1;
      patterns[43411] = 25'b10101001_10010001_00111010_1;
      patterns[43412] = 25'b10101001_10010010_00111011_1;
      patterns[43413] = 25'b10101001_10010011_00111100_1;
      patterns[43414] = 25'b10101001_10010100_00111101_1;
      patterns[43415] = 25'b10101001_10010101_00111110_1;
      patterns[43416] = 25'b10101001_10010110_00111111_1;
      patterns[43417] = 25'b10101001_10010111_01000000_1;
      patterns[43418] = 25'b10101001_10011000_01000001_1;
      patterns[43419] = 25'b10101001_10011001_01000010_1;
      patterns[43420] = 25'b10101001_10011010_01000011_1;
      patterns[43421] = 25'b10101001_10011011_01000100_1;
      patterns[43422] = 25'b10101001_10011100_01000101_1;
      patterns[43423] = 25'b10101001_10011101_01000110_1;
      patterns[43424] = 25'b10101001_10011110_01000111_1;
      patterns[43425] = 25'b10101001_10011111_01001000_1;
      patterns[43426] = 25'b10101001_10100000_01001001_1;
      patterns[43427] = 25'b10101001_10100001_01001010_1;
      patterns[43428] = 25'b10101001_10100010_01001011_1;
      patterns[43429] = 25'b10101001_10100011_01001100_1;
      patterns[43430] = 25'b10101001_10100100_01001101_1;
      patterns[43431] = 25'b10101001_10100101_01001110_1;
      patterns[43432] = 25'b10101001_10100110_01001111_1;
      patterns[43433] = 25'b10101001_10100111_01010000_1;
      patterns[43434] = 25'b10101001_10101000_01010001_1;
      patterns[43435] = 25'b10101001_10101001_01010010_1;
      patterns[43436] = 25'b10101001_10101010_01010011_1;
      patterns[43437] = 25'b10101001_10101011_01010100_1;
      patterns[43438] = 25'b10101001_10101100_01010101_1;
      patterns[43439] = 25'b10101001_10101101_01010110_1;
      patterns[43440] = 25'b10101001_10101110_01010111_1;
      patterns[43441] = 25'b10101001_10101111_01011000_1;
      patterns[43442] = 25'b10101001_10110000_01011001_1;
      patterns[43443] = 25'b10101001_10110001_01011010_1;
      patterns[43444] = 25'b10101001_10110010_01011011_1;
      patterns[43445] = 25'b10101001_10110011_01011100_1;
      patterns[43446] = 25'b10101001_10110100_01011101_1;
      patterns[43447] = 25'b10101001_10110101_01011110_1;
      patterns[43448] = 25'b10101001_10110110_01011111_1;
      patterns[43449] = 25'b10101001_10110111_01100000_1;
      patterns[43450] = 25'b10101001_10111000_01100001_1;
      patterns[43451] = 25'b10101001_10111001_01100010_1;
      patterns[43452] = 25'b10101001_10111010_01100011_1;
      patterns[43453] = 25'b10101001_10111011_01100100_1;
      patterns[43454] = 25'b10101001_10111100_01100101_1;
      patterns[43455] = 25'b10101001_10111101_01100110_1;
      patterns[43456] = 25'b10101001_10111110_01100111_1;
      patterns[43457] = 25'b10101001_10111111_01101000_1;
      patterns[43458] = 25'b10101001_11000000_01101001_1;
      patterns[43459] = 25'b10101001_11000001_01101010_1;
      patterns[43460] = 25'b10101001_11000010_01101011_1;
      patterns[43461] = 25'b10101001_11000011_01101100_1;
      patterns[43462] = 25'b10101001_11000100_01101101_1;
      patterns[43463] = 25'b10101001_11000101_01101110_1;
      patterns[43464] = 25'b10101001_11000110_01101111_1;
      patterns[43465] = 25'b10101001_11000111_01110000_1;
      patterns[43466] = 25'b10101001_11001000_01110001_1;
      patterns[43467] = 25'b10101001_11001001_01110010_1;
      patterns[43468] = 25'b10101001_11001010_01110011_1;
      patterns[43469] = 25'b10101001_11001011_01110100_1;
      patterns[43470] = 25'b10101001_11001100_01110101_1;
      patterns[43471] = 25'b10101001_11001101_01110110_1;
      patterns[43472] = 25'b10101001_11001110_01110111_1;
      patterns[43473] = 25'b10101001_11001111_01111000_1;
      patterns[43474] = 25'b10101001_11010000_01111001_1;
      patterns[43475] = 25'b10101001_11010001_01111010_1;
      patterns[43476] = 25'b10101001_11010010_01111011_1;
      patterns[43477] = 25'b10101001_11010011_01111100_1;
      patterns[43478] = 25'b10101001_11010100_01111101_1;
      patterns[43479] = 25'b10101001_11010101_01111110_1;
      patterns[43480] = 25'b10101001_11010110_01111111_1;
      patterns[43481] = 25'b10101001_11010111_10000000_1;
      patterns[43482] = 25'b10101001_11011000_10000001_1;
      patterns[43483] = 25'b10101001_11011001_10000010_1;
      patterns[43484] = 25'b10101001_11011010_10000011_1;
      patterns[43485] = 25'b10101001_11011011_10000100_1;
      patterns[43486] = 25'b10101001_11011100_10000101_1;
      patterns[43487] = 25'b10101001_11011101_10000110_1;
      patterns[43488] = 25'b10101001_11011110_10000111_1;
      patterns[43489] = 25'b10101001_11011111_10001000_1;
      patterns[43490] = 25'b10101001_11100000_10001001_1;
      patterns[43491] = 25'b10101001_11100001_10001010_1;
      patterns[43492] = 25'b10101001_11100010_10001011_1;
      patterns[43493] = 25'b10101001_11100011_10001100_1;
      patterns[43494] = 25'b10101001_11100100_10001101_1;
      patterns[43495] = 25'b10101001_11100101_10001110_1;
      patterns[43496] = 25'b10101001_11100110_10001111_1;
      patterns[43497] = 25'b10101001_11100111_10010000_1;
      patterns[43498] = 25'b10101001_11101000_10010001_1;
      patterns[43499] = 25'b10101001_11101001_10010010_1;
      patterns[43500] = 25'b10101001_11101010_10010011_1;
      patterns[43501] = 25'b10101001_11101011_10010100_1;
      patterns[43502] = 25'b10101001_11101100_10010101_1;
      patterns[43503] = 25'b10101001_11101101_10010110_1;
      patterns[43504] = 25'b10101001_11101110_10010111_1;
      patterns[43505] = 25'b10101001_11101111_10011000_1;
      patterns[43506] = 25'b10101001_11110000_10011001_1;
      patterns[43507] = 25'b10101001_11110001_10011010_1;
      patterns[43508] = 25'b10101001_11110010_10011011_1;
      patterns[43509] = 25'b10101001_11110011_10011100_1;
      patterns[43510] = 25'b10101001_11110100_10011101_1;
      patterns[43511] = 25'b10101001_11110101_10011110_1;
      patterns[43512] = 25'b10101001_11110110_10011111_1;
      patterns[43513] = 25'b10101001_11110111_10100000_1;
      patterns[43514] = 25'b10101001_11111000_10100001_1;
      patterns[43515] = 25'b10101001_11111001_10100010_1;
      patterns[43516] = 25'b10101001_11111010_10100011_1;
      patterns[43517] = 25'b10101001_11111011_10100100_1;
      patterns[43518] = 25'b10101001_11111100_10100101_1;
      patterns[43519] = 25'b10101001_11111101_10100110_1;
      patterns[43520] = 25'b10101001_11111110_10100111_1;
      patterns[43521] = 25'b10101001_11111111_10101000_1;
      patterns[43522] = 25'b10101010_00000000_10101010_0;
      patterns[43523] = 25'b10101010_00000001_10101011_0;
      patterns[43524] = 25'b10101010_00000010_10101100_0;
      patterns[43525] = 25'b10101010_00000011_10101101_0;
      patterns[43526] = 25'b10101010_00000100_10101110_0;
      patterns[43527] = 25'b10101010_00000101_10101111_0;
      patterns[43528] = 25'b10101010_00000110_10110000_0;
      patterns[43529] = 25'b10101010_00000111_10110001_0;
      patterns[43530] = 25'b10101010_00001000_10110010_0;
      patterns[43531] = 25'b10101010_00001001_10110011_0;
      patterns[43532] = 25'b10101010_00001010_10110100_0;
      patterns[43533] = 25'b10101010_00001011_10110101_0;
      patterns[43534] = 25'b10101010_00001100_10110110_0;
      patterns[43535] = 25'b10101010_00001101_10110111_0;
      patterns[43536] = 25'b10101010_00001110_10111000_0;
      patterns[43537] = 25'b10101010_00001111_10111001_0;
      patterns[43538] = 25'b10101010_00010000_10111010_0;
      patterns[43539] = 25'b10101010_00010001_10111011_0;
      patterns[43540] = 25'b10101010_00010010_10111100_0;
      patterns[43541] = 25'b10101010_00010011_10111101_0;
      patterns[43542] = 25'b10101010_00010100_10111110_0;
      patterns[43543] = 25'b10101010_00010101_10111111_0;
      patterns[43544] = 25'b10101010_00010110_11000000_0;
      patterns[43545] = 25'b10101010_00010111_11000001_0;
      patterns[43546] = 25'b10101010_00011000_11000010_0;
      patterns[43547] = 25'b10101010_00011001_11000011_0;
      patterns[43548] = 25'b10101010_00011010_11000100_0;
      patterns[43549] = 25'b10101010_00011011_11000101_0;
      patterns[43550] = 25'b10101010_00011100_11000110_0;
      patterns[43551] = 25'b10101010_00011101_11000111_0;
      patterns[43552] = 25'b10101010_00011110_11001000_0;
      patterns[43553] = 25'b10101010_00011111_11001001_0;
      patterns[43554] = 25'b10101010_00100000_11001010_0;
      patterns[43555] = 25'b10101010_00100001_11001011_0;
      patterns[43556] = 25'b10101010_00100010_11001100_0;
      patterns[43557] = 25'b10101010_00100011_11001101_0;
      patterns[43558] = 25'b10101010_00100100_11001110_0;
      patterns[43559] = 25'b10101010_00100101_11001111_0;
      patterns[43560] = 25'b10101010_00100110_11010000_0;
      patterns[43561] = 25'b10101010_00100111_11010001_0;
      patterns[43562] = 25'b10101010_00101000_11010010_0;
      patterns[43563] = 25'b10101010_00101001_11010011_0;
      patterns[43564] = 25'b10101010_00101010_11010100_0;
      patterns[43565] = 25'b10101010_00101011_11010101_0;
      patterns[43566] = 25'b10101010_00101100_11010110_0;
      patterns[43567] = 25'b10101010_00101101_11010111_0;
      patterns[43568] = 25'b10101010_00101110_11011000_0;
      patterns[43569] = 25'b10101010_00101111_11011001_0;
      patterns[43570] = 25'b10101010_00110000_11011010_0;
      patterns[43571] = 25'b10101010_00110001_11011011_0;
      patterns[43572] = 25'b10101010_00110010_11011100_0;
      patterns[43573] = 25'b10101010_00110011_11011101_0;
      patterns[43574] = 25'b10101010_00110100_11011110_0;
      patterns[43575] = 25'b10101010_00110101_11011111_0;
      patterns[43576] = 25'b10101010_00110110_11100000_0;
      patterns[43577] = 25'b10101010_00110111_11100001_0;
      patterns[43578] = 25'b10101010_00111000_11100010_0;
      patterns[43579] = 25'b10101010_00111001_11100011_0;
      patterns[43580] = 25'b10101010_00111010_11100100_0;
      patterns[43581] = 25'b10101010_00111011_11100101_0;
      patterns[43582] = 25'b10101010_00111100_11100110_0;
      patterns[43583] = 25'b10101010_00111101_11100111_0;
      patterns[43584] = 25'b10101010_00111110_11101000_0;
      patterns[43585] = 25'b10101010_00111111_11101001_0;
      patterns[43586] = 25'b10101010_01000000_11101010_0;
      patterns[43587] = 25'b10101010_01000001_11101011_0;
      patterns[43588] = 25'b10101010_01000010_11101100_0;
      patterns[43589] = 25'b10101010_01000011_11101101_0;
      patterns[43590] = 25'b10101010_01000100_11101110_0;
      patterns[43591] = 25'b10101010_01000101_11101111_0;
      patterns[43592] = 25'b10101010_01000110_11110000_0;
      patterns[43593] = 25'b10101010_01000111_11110001_0;
      patterns[43594] = 25'b10101010_01001000_11110010_0;
      patterns[43595] = 25'b10101010_01001001_11110011_0;
      patterns[43596] = 25'b10101010_01001010_11110100_0;
      patterns[43597] = 25'b10101010_01001011_11110101_0;
      patterns[43598] = 25'b10101010_01001100_11110110_0;
      patterns[43599] = 25'b10101010_01001101_11110111_0;
      patterns[43600] = 25'b10101010_01001110_11111000_0;
      patterns[43601] = 25'b10101010_01001111_11111001_0;
      patterns[43602] = 25'b10101010_01010000_11111010_0;
      patterns[43603] = 25'b10101010_01010001_11111011_0;
      patterns[43604] = 25'b10101010_01010010_11111100_0;
      patterns[43605] = 25'b10101010_01010011_11111101_0;
      patterns[43606] = 25'b10101010_01010100_11111110_0;
      patterns[43607] = 25'b10101010_01010101_11111111_0;
      patterns[43608] = 25'b10101010_01010110_00000000_1;
      patterns[43609] = 25'b10101010_01010111_00000001_1;
      patterns[43610] = 25'b10101010_01011000_00000010_1;
      patterns[43611] = 25'b10101010_01011001_00000011_1;
      patterns[43612] = 25'b10101010_01011010_00000100_1;
      patterns[43613] = 25'b10101010_01011011_00000101_1;
      patterns[43614] = 25'b10101010_01011100_00000110_1;
      patterns[43615] = 25'b10101010_01011101_00000111_1;
      patterns[43616] = 25'b10101010_01011110_00001000_1;
      patterns[43617] = 25'b10101010_01011111_00001001_1;
      patterns[43618] = 25'b10101010_01100000_00001010_1;
      patterns[43619] = 25'b10101010_01100001_00001011_1;
      patterns[43620] = 25'b10101010_01100010_00001100_1;
      patterns[43621] = 25'b10101010_01100011_00001101_1;
      patterns[43622] = 25'b10101010_01100100_00001110_1;
      patterns[43623] = 25'b10101010_01100101_00001111_1;
      patterns[43624] = 25'b10101010_01100110_00010000_1;
      patterns[43625] = 25'b10101010_01100111_00010001_1;
      patterns[43626] = 25'b10101010_01101000_00010010_1;
      patterns[43627] = 25'b10101010_01101001_00010011_1;
      patterns[43628] = 25'b10101010_01101010_00010100_1;
      patterns[43629] = 25'b10101010_01101011_00010101_1;
      patterns[43630] = 25'b10101010_01101100_00010110_1;
      patterns[43631] = 25'b10101010_01101101_00010111_1;
      patterns[43632] = 25'b10101010_01101110_00011000_1;
      patterns[43633] = 25'b10101010_01101111_00011001_1;
      patterns[43634] = 25'b10101010_01110000_00011010_1;
      patterns[43635] = 25'b10101010_01110001_00011011_1;
      patterns[43636] = 25'b10101010_01110010_00011100_1;
      patterns[43637] = 25'b10101010_01110011_00011101_1;
      patterns[43638] = 25'b10101010_01110100_00011110_1;
      patterns[43639] = 25'b10101010_01110101_00011111_1;
      patterns[43640] = 25'b10101010_01110110_00100000_1;
      patterns[43641] = 25'b10101010_01110111_00100001_1;
      patterns[43642] = 25'b10101010_01111000_00100010_1;
      patterns[43643] = 25'b10101010_01111001_00100011_1;
      patterns[43644] = 25'b10101010_01111010_00100100_1;
      patterns[43645] = 25'b10101010_01111011_00100101_1;
      patterns[43646] = 25'b10101010_01111100_00100110_1;
      patterns[43647] = 25'b10101010_01111101_00100111_1;
      patterns[43648] = 25'b10101010_01111110_00101000_1;
      patterns[43649] = 25'b10101010_01111111_00101001_1;
      patterns[43650] = 25'b10101010_10000000_00101010_1;
      patterns[43651] = 25'b10101010_10000001_00101011_1;
      patterns[43652] = 25'b10101010_10000010_00101100_1;
      patterns[43653] = 25'b10101010_10000011_00101101_1;
      patterns[43654] = 25'b10101010_10000100_00101110_1;
      patterns[43655] = 25'b10101010_10000101_00101111_1;
      patterns[43656] = 25'b10101010_10000110_00110000_1;
      patterns[43657] = 25'b10101010_10000111_00110001_1;
      patterns[43658] = 25'b10101010_10001000_00110010_1;
      patterns[43659] = 25'b10101010_10001001_00110011_1;
      patterns[43660] = 25'b10101010_10001010_00110100_1;
      patterns[43661] = 25'b10101010_10001011_00110101_1;
      patterns[43662] = 25'b10101010_10001100_00110110_1;
      patterns[43663] = 25'b10101010_10001101_00110111_1;
      patterns[43664] = 25'b10101010_10001110_00111000_1;
      patterns[43665] = 25'b10101010_10001111_00111001_1;
      patterns[43666] = 25'b10101010_10010000_00111010_1;
      patterns[43667] = 25'b10101010_10010001_00111011_1;
      patterns[43668] = 25'b10101010_10010010_00111100_1;
      patterns[43669] = 25'b10101010_10010011_00111101_1;
      patterns[43670] = 25'b10101010_10010100_00111110_1;
      patterns[43671] = 25'b10101010_10010101_00111111_1;
      patterns[43672] = 25'b10101010_10010110_01000000_1;
      patterns[43673] = 25'b10101010_10010111_01000001_1;
      patterns[43674] = 25'b10101010_10011000_01000010_1;
      patterns[43675] = 25'b10101010_10011001_01000011_1;
      patterns[43676] = 25'b10101010_10011010_01000100_1;
      patterns[43677] = 25'b10101010_10011011_01000101_1;
      patterns[43678] = 25'b10101010_10011100_01000110_1;
      patterns[43679] = 25'b10101010_10011101_01000111_1;
      patterns[43680] = 25'b10101010_10011110_01001000_1;
      patterns[43681] = 25'b10101010_10011111_01001001_1;
      patterns[43682] = 25'b10101010_10100000_01001010_1;
      patterns[43683] = 25'b10101010_10100001_01001011_1;
      patterns[43684] = 25'b10101010_10100010_01001100_1;
      patterns[43685] = 25'b10101010_10100011_01001101_1;
      patterns[43686] = 25'b10101010_10100100_01001110_1;
      patterns[43687] = 25'b10101010_10100101_01001111_1;
      patterns[43688] = 25'b10101010_10100110_01010000_1;
      patterns[43689] = 25'b10101010_10100111_01010001_1;
      patterns[43690] = 25'b10101010_10101000_01010010_1;
      patterns[43691] = 25'b10101010_10101001_01010011_1;
      patterns[43692] = 25'b10101010_10101010_01010100_1;
      patterns[43693] = 25'b10101010_10101011_01010101_1;
      patterns[43694] = 25'b10101010_10101100_01010110_1;
      patterns[43695] = 25'b10101010_10101101_01010111_1;
      patterns[43696] = 25'b10101010_10101110_01011000_1;
      patterns[43697] = 25'b10101010_10101111_01011001_1;
      patterns[43698] = 25'b10101010_10110000_01011010_1;
      patterns[43699] = 25'b10101010_10110001_01011011_1;
      patterns[43700] = 25'b10101010_10110010_01011100_1;
      patterns[43701] = 25'b10101010_10110011_01011101_1;
      patterns[43702] = 25'b10101010_10110100_01011110_1;
      patterns[43703] = 25'b10101010_10110101_01011111_1;
      patterns[43704] = 25'b10101010_10110110_01100000_1;
      patterns[43705] = 25'b10101010_10110111_01100001_1;
      patterns[43706] = 25'b10101010_10111000_01100010_1;
      patterns[43707] = 25'b10101010_10111001_01100011_1;
      patterns[43708] = 25'b10101010_10111010_01100100_1;
      patterns[43709] = 25'b10101010_10111011_01100101_1;
      patterns[43710] = 25'b10101010_10111100_01100110_1;
      patterns[43711] = 25'b10101010_10111101_01100111_1;
      patterns[43712] = 25'b10101010_10111110_01101000_1;
      patterns[43713] = 25'b10101010_10111111_01101001_1;
      patterns[43714] = 25'b10101010_11000000_01101010_1;
      patterns[43715] = 25'b10101010_11000001_01101011_1;
      patterns[43716] = 25'b10101010_11000010_01101100_1;
      patterns[43717] = 25'b10101010_11000011_01101101_1;
      patterns[43718] = 25'b10101010_11000100_01101110_1;
      patterns[43719] = 25'b10101010_11000101_01101111_1;
      patterns[43720] = 25'b10101010_11000110_01110000_1;
      patterns[43721] = 25'b10101010_11000111_01110001_1;
      patterns[43722] = 25'b10101010_11001000_01110010_1;
      patterns[43723] = 25'b10101010_11001001_01110011_1;
      patterns[43724] = 25'b10101010_11001010_01110100_1;
      patterns[43725] = 25'b10101010_11001011_01110101_1;
      patterns[43726] = 25'b10101010_11001100_01110110_1;
      patterns[43727] = 25'b10101010_11001101_01110111_1;
      patterns[43728] = 25'b10101010_11001110_01111000_1;
      patterns[43729] = 25'b10101010_11001111_01111001_1;
      patterns[43730] = 25'b10101010_11010000_01111010_1;
      patterns[43731] = 25'b10101010_11010001_01111011_1;
      patterns[43732] = 25'b10101010_11010010_01111100_1;
      patterns[43733] = 25'b10101010_11010011_01111101_1;
      patterns[43734] = 25'b10101010_11010100_01111110_1;
      patterns[43735] = 25'b10101010_11010101_01111111_1;
      patterns[43736] = 25'b10101010_11010110_10000000_1;
      patterns[43737] = 25'b10101010_11010111_10000001_1;
      patterns[43738] = 25'b10101010_11011000_10000010_1;
      patterns[43739] = 25'b10101010_11011001_10000011_1;
      patterns[43740] = 25'b10101010_11011010_10000100_1;
      patterns[43741] = 25'b10101010_11011011_10000101_1;
      patterns[43742] = 25'b10101010_11011100_10000110_1;
      patterns[43743] = 25'b10101010_11011101_10000111_1;
      patterns[43744] = 25'b10101010_11011110_10001000_1;
      patterns[43745] = 25'b10101010_11011111_10001001_1;
      patterns[43746] = 25'b10101010_11100000_10001010_1;
      patterns[43747] = 25'b10101010_11100001_10001011_1;
      patterns[43748] = 25'b10101010_11100010_10001100_1;
      patterns[43749] = 25'b10101010_11100011_10001101_1;
      patterns[43750] = 25'b10101010_11100100_10001110_1;
      patterns[43751] = 25'b10101010_11100101_10001111_1;
      patterns[43752] = 25'b10101010_11100110_10010000_1;
      patterns[43753] = 25'b10101010_11100111_10010001_1;
      patterns[43754] = 25'b10101010_11101000_10010010_1;
      patterns[43755] = 25'b10101010_11101001_10010011_1;
      patterns[43756] = 25'b10101010_11101010_10010100_1;
      patterns[43757] = 25'b10101010_11101011_10010101_1;
      patterns[43758] = 25'b10101010_11101100_10010110_1;
      patterns[43759] = 25'b10101010_11101101_10010111_1;
      patterns[43760] = 25'b10101010_11101110_10011000_1;
      patterns[43761] = 25'b10101010_11101111_10011001_1;
      patterns[43762] = 25'b10101010_11110000_10011010_1;
      patterns[43763] = 25'b10101010_11110001_10011011_1;
      patterns[43764] = 25'b10101010_11110010_10011100_1;
      patterns[43765] = 25'b10101010_11110011_10011101_1;
      patterns[43766] = 25'b10101010_11110100_10011110_1;
      patterns[43767] = 25'b10101010_11110101_10011111_1;
      patterns[43768] = 25'b10101010_11110110_10100000_1;
      patterns[43769] = 25'b10101010_11110111_10100001_1;
      patterns[43770] = 25'b10101010_11111000_10100010_1;
      patterns[43771] = 25'b10101010_11111001_10100011_1;
      patterns[43772] = 25'b10101010_11111010_10100100_1;
      patterns[43773] = 25'b10101010_11111011_10100101_1;
      patterns[43774] = 25'b10101010_11111100_10100110_1;
      patterns[43775] = 25'b10101010_11111101_10100111_1;
      patterns[43776] = 25'b10101010_11111110_10101000_1;
      patterns[43777] = 25'b10101010_11111111_10101001_1;
      patterns[43778] = 25'b10101011_00000000_10101011_0;
      patterns[43779] = 25'b10101011_00000001_10101100_0;
      patterns[43780] = 25'b10101011_00000010_10101101_0;
      patterns[43781] = 25'b10101011_00000011_10101110_0;
      patterns[43782] = 25'b10101011_00000100_10101111_0;
      patterns[43783] = 25'b10101011_00000101_10110000_0;
      patterns[43784] = 25'b10101011_00000110_10110001_0;
      patterns[43785] = 25'b10101011_00000111_10110010_0;
      patterns[43786] = 25'b10101011_00001000_10110011_0;
      patterns[43787] = 25'b10101011_00001001_10110100_0;
      patterns[43788] = 25'b10101011_00001010_10110101_0;
      patterns[43789] = 25'b10101011_00001011_10110110_0;
      patterns[43790] = 25'b10101011_00001100_10110111_0;
      patterns[43791] = 25'b10101011_00001101_10111000_0;
      patterns[43792] = 25'b10101011_00001110_10111001_0;
      patterns[43793] = 25'b10101011_00001111_10111010_0;
      patterns[43794] = 25'b10101011_00010000_10111011_0;
      patterns[43795] = 25'b10101011_00010001_10111100_0;
      patterns[43796] = 25'b10101011_00010010_10111101_0;
      patterns[43797] = 25'b10101011_00010011_10111110_0;
      patterns[43798] = 25'b10101011_00010100_10111111_0;
      patterns[43799] = 25'b10101011_00010101_11000000_0;
      patterns[43800] = 25'b10101011_00010110_11000001_0;
      patterns[43801] = 25'b10101011_00010111_11000010_0;
      patterns[43802] = 25'b10101011_00011000_11000011_0;
      patterns[43803] = 25'b10101011_00011001_11000100_0;
      patterns[43804] = 25'b10101011_00011010_11000101_0;
      patterns[43805] = 25'b10101011_00011011_11000110_0;
      patterns[43806] = 25'b10101011_00011100_11000111_0;
      patterns[43807] = 25'b10101011_00011101_11001000_0;
      patterns[43808] = 25'b10101011_00011110_11001001_0;
      patterns[43809] = 25'b10101011_00011111_11001010_0;
      patterns[43810] = 25'b10101011_00100000_11001011_0;
      patterns[43811] = 25'b10101011_00100001_11001100_0;
      patterns[43812] = 25'b10101011_00100010_11001101_0;
      patterns[43813] = 25'b10101011_00100011_11001110_0;
      patterns[43814] = 25'b10101011_00100100_11001111_0;
      patterns[43815] = 25'b10101011_00100101_11010000_0;
      patterns[43816] = 25'b10101011_00100110_11010001_0;
      patterns[43817] = 25'b10101011_00100111_11010010_0;
      patterns[43818] = 25'b10101011_00101000_11010011_0;
      patterns[43819] = 25'b10101011_00101001_11010100_0;
      patterns[43820] = 25'b10101011_00101010_11010101_0;
      patterns[43821] = 25'b10101011_00101011_11010110_0;
      patterns[43822] = 25'b10101011_00101100_11010111_0;
      patterns[43823] = 25'b10101011_00101101_11011000_0;
      patterns[43824] = 25'b10101011_00101110_11011001_0;
      patterns[43825] = 25'b10101011_00101111_11011010_0;
      patterns[43826] = 25'b10101011_00110000_11011011_0;
      patterns[43827] = 25'b10101011_00110001_11011100_0;
      patterns[43828] = 25'b10101011_00110010_11011101_0;
      patterns[43829] = 25'b10101011_00110011_11011110_0;
      patterns[43830] = 25'b10101011_00110100_11011111_0;
      patterns[43831] = 25'b10101011_00110101_11100000_0;
      patterns[43832] = 25'b10101011_00110110_11100001_0;
      patterns[43833] = 25'b10101011_00110111_11100010_0;
      patterns[43834] = 25'b10101011_00111000_11100011_0;
      patterns[43835] = 25'b10101011_00111001_11100100_0;
      patterns[43836] = 25'b10101011_00111010_11100101_0;
      patterns[43837] = 25'b10101011_00111011_11100110_0;
      patterns[43838] = 25'b10101011_00111100_11100111_0;
      patterns[43839] = 25'b10101011_00111101_11101000_0;
      patterns[43840] = 25'b10101011_00111110_11101001_0;
      patterns[43841] = 25'b10101011_00111111_11101010_0;
      patterns[43842] = 25'b10101011_01000000_11101011_0;
      patterns[43843] = 25'b10101011_01000001_11101100_0;
      patterns[43844] = 25'b10101011_01000010_11101101_0;
      patterns[43845] = 25'b10101011_01000011_11101110_0;
      patterns[43846] = 25'b10101011_01000100_11101111_0;
      patterns[43847] = 25'b10101011_01000101_11110000_0;
      patterns[43848] = 25'b10101011_01000110_11110001_0;
      patterns[43849] = 25'b10101011_01000111_11110010_0;
      patterns[43850] = 25'b10101011_01001000_11110011_0;
      patterns[43851] = 25'b10101011_01001001_11110100_0;
      patterns[43852] = 25'b10101011_01001010_11110101_0;
      patterns[43853] = 25'b10101011_01001011_11110110_0;
      patterns[43854] = 25'b10101011_01001100_11110111_0;
      patterns[43855] = 25'b10101011_01001101_11111000_0;
      patterns[43856] = 25'b10101011_01001110_11111001_0;
      patterns[43857] = 25'b10101011_01001111_11111010_0;
      patterns[43858] = 25'b10101011_01010000_11111011_0;
      patterns[43859] = 25'b10101011_01010001_11111100_0;
      patterns[43860] = 25'b10101011_01010010_11111101_0;
      patterns[43861] = 25'b10101011_01010011_11111110_0;
      patterns[43862] = 25'b10101011_01010100_11111111_0;
      patterns[43863] = 25'b10101011_01010101_00000000_1;
      patterns[43864] = 25'b10101011_01010110_00000001_1;
      patterns[43865] = 25'b10101011_01010111_00000010_1;
      patterns[43866] = 25'b10101011_01011000_00000011_1;
      patterns[43867] = 25'b10101011_01011001_00000100_1;
      patterns[43868] = 25'b10101011_01011010_00000101_1;
      patterns[43869] = 25'b10101011_01011011_00000110_1;
      patterns[43870] = 25'b10101011_01011100_00000111_1;
      patterns[43871] = 25'b10101011_01011101_00001000_1;
      patterns[43872] = 25'b10101011_01011110_00001001_1;
      patterns[43873] = 25'b10101011_01011111_00001010_1;
      patterns[43874] = 25'b10101011_01100000_00001011_1;
      patterns[43875] = 25'b10101011_01100001_00001100_1;
      patterns[43876] = 25'b10101011_01100010_00001101_1;
      patterns[43877] = 25'b10101011_01100011_00001110_1;
      patterns[43878] = 25'b10101011_01100100_00001111_1;
      patterns[43879] = 25'b10101011_01100101_00010000_1;
      patterns[43880] = 25'b10101011_01100110_00010001_1;
      patterns[43881] = 25'b10101011_01100111_00010010_1;
      patterns[43882] = 25'b10101011_01101000_00010011_1;
      patterns[43883] = 25'b10101011_01101001_00010100_1;
      patterns[43884] = 25'b10101011_01101010_00010101_1;
      patterns[43885] = 25'b10101011_01101011_00010110_1;
      patterns[43886] = 25'b10101011_01101100_00010111_1;
      patterns[43887] = 25'b10101011_01101101_00011000_1;
      patterns[43888] = 25'b10101011_01101110_00011001_1;
      patterns[43889] = 25'b10101011_01101111_00011010_1;
      patterns[43890] = 25'b10101011_01110000_00011011_1;
      patterns[43891] = 25'b10101011_01110001_00011100_1;
      patterns[43892] = 25'b10101011_01110010_00011101_1;
      patterns[43893] = 25'b10101011_01110011_00011110_1;
      patterns[43894] = 25'b10101011_01110100_00011111_1;
      patterns[43895] = 25'b10101011_01110101_00100000_1;
      patterns[43896] = 25'b10101011_01110110_00100001_1;
      patterns[43897] = 25'b10101011_01110111_00100010_1;
      patterns[43898] = 25'b10101011_01111000_00100011_1;
      patterns[43899] = 25'b10101011_01111001_00100100_1;
      patterns[43900] = 25'b10101011_01111010_00100101_1;
      patterns[43901] = 25'b10101011_01111011_00100110_1;
      patterns[43902] = 25'b10101011_01111100_00100111_1;
      patterns[43903] = 25'b10101011_01111101_00101000_1;
      patterns[43904] = 25'b10101011_01111110_00101001_1;
      patterns[43905] = 25'b10101011_01111111_00101010_1;
      patterns[43906] = 25'b10101011_10000000_00101011_1;
      patterns[43907] = 25'b10101011_10000001_00101100_1;
      patterns[43908] = 25'b10101011_10000010_00101101_1;
      patterns[43909] = 25'b10101011_10000011_00101110_1;
      patterns[43910] = 25'b10101011_10000100_00101111_1;
      patterns[43911] = 25'b10101011_10000101_00110000_1;
      patterns[43912] = 25'b10101011_10000110_00110001_1;
      patterns[43913] = 25'b10101011_10000111_00110010_1;
      patterns[43914] = 25'b10101011_10001000_00110011_1;
      patterns[43915] = 25'b10101011_10001001_00110100_1;
      patterns[43916] = 25'b10101011_10001010_00110101_1;
      patterns[43917] = 25'b10101011_10001011_00110110_1;
      patterns[43918] = 25'b10101011_10001100_00110111_1;
      patterns[43919] = 25'b10101011_10001101_00111000_1;
      patterns[43920] = 25'b10101011_10001110_00111001_1;
      patterns[43921] = 25'b10101011_10001111_00111010_1;
      patterns[43922] = 25'b10101011_10010000_00111011_1;
      patterns[43923] = 25'b10101011_10010001_00111100_1;
      patterns[43924] = 25'b10101011_10010010_00111101_1;
      patterns[43925] = 25'b10101011_10010011_00111110_1;
      patterns[43926] = 25'b10101011_10010100_00111111_1;
      patterns[43927] = 25'b10101011_10010101_01000000_1;
      patterns[43928] = 25'b10101011_10010110_01000001_1;
      patterns[43929] = 25'b10101011_10010111_01000010_1;
      patterns[43930] = 25'b10101011_10011000_01000011_1;
      patterns[43931] = 25'b10101011_10011001_01000100_1;
      patterns[43932] = 25'b10101011_10011010_01000101_1;
      patterns[43933] = 25'b10101011_10011011_01000110_1;
      patterns[43934] = 25'b10101011_10011100_01000111_1;
      patterns[43935] = 25'b10101011_10011101_01001000_1;
      patterns[43936] = 25'b10101011_10011110_01001001_1;
      patterns[43937] = 25'b10101011_10011111_01001010_1;
      patterns[43938] = 25'b10101011_10100000_01001011_1;
      patterns[43939] = 25'b10101011_10100001_01001100_1;
      patterns[43940] = 25'b10101011_10100010_01001101_1;
      patterns[43941] = 25'b10101011_10100011_01001110_1;
      patterns[43942] = 25'b10101011_10100100_01001111_1;
      patterns[43943] = 25'b10101011_10100101_01010000_1;
      patterns[43944] = 25'b10101011_10100110_01010001_1;
      patterns[43945] = 25'b10101011_10100111_01010010_1;
      patterns[43946] = 25'b10101011_10101000_01010011_1;
      patterns[43947] = 25'b10101011_10101001_01010100_1;
      patterns[43948] = 25'b10101011_10101010_01010101_1;
      patterns[43949] = 25'b10101011_10101011_01010110_1;
      patterns[43950] = 25'b10101011_10101100_01010111_1;
      patterns[43951] = 25'b10101011_10101101_01011000_1;
      patterns[43952] = 25'b10101011_10101110_01011001_1;
      patterns[43953] = 25'b10101011_10101111_01011010_1;
      patterns[43954] = 25'b10101011_10110000_01011011_1;
      patterns[43955] = 25'b10101011_10110001_01011100_1;
      patterns[43956] = 25'b10101011_10110010_01011101_1;
      patterns[43957] = 25'b10101011_10110011_01011110_1;
      patterns[43958] = 25'b10101011_10110100_01011111_1;
      patterns[43959] = 25'b10101011_10110101_01100000_1;
      patterns[43960] = 25'b10101011_10110110_01100001_1;
      patterns[43961] = 25'b10101011_10110111_01100010_1;
      patterns[43962] = 25'b10101011_10111000_01100011_1;
      patterns[43963] = 25'b10101011_10111001_01100100_1;
      patterns[43964] = 25'b10101011_10111010_01100101_1;
      patterns[43965] = 25'b10101011_10111011_01100110_1;
      patterns[43966] = 25'b10101011_10111100_01100111_1;
      patterns[43967] = 25'b10101011_10111101_01101000_1;
      patterns[43968] = 25'b10101011_10111110_01101001_1;
      patterns[43969] = 25'b10101011_10111111_01101010_1;
      patterns[43970] = 25'b10101011_11000000_01101011_1;
      patterns[43971] = 25'b10101011_11000001_01101100_1;
      patterns[43972] = 25'b10101011_11000010_01101101_1;
      patterns[43973] = 25'b10101011_11000011_01101110_1;
      patterns[43974] = 25'b10101011_11000100_01101111_1;
      patterns[43975] = 25'b10101011_11000101_01110000_1;
      patterns[43976] = 25'b10101011_11000110_01110001_1;
      patterns[43977] = 25'b10101011_11000111_01110010_1;
      patterns[43978] = 25'b10101011_11001000_01110011_1;
      patterns[43979] = 25'b10101011_11001001_01110100_1;
      patterns[43980] = 25'b10101011_11001010_01110101_1;
      patterns[43981] = 25'b10101011_11001011_01110110_1;
      patterns[43982] = 25'b10101011_11001100_01110111_1;
      patterns[43983] = 25'b10101011_11001101_01111000_1;
      patterns[43984] = 25'b10101011_11001110_01111001_1;
      patterns[43985] = 25'b10101011_11001111_01111010_1;
      patterns[43986] = 25'b10101011_11010000_01111011_1;
      patterns[43987] = 25'b10101011_11010001_01111100_1;
      patterns[43988] = 25'b10101011_11010010_01111101_1;
      patterns[43989] = 25'b10101011_11010011_01111110_1;
      patterns[43990] = 25'b10101011_11010100_01111111_1;
      patterns[43991] = 25'b10101011_11010101_10000000_1;
      patterns[43992] = 25'b10101011_11010110_10000001_1;
      patterns[43993] = 25'b10101011_11010111_10000010_1;
      patterns[43994] = 25'b10101011_11011000_10000011_1;
      patterns[43995] = 25'b10101011_11011001_10000100_1;
      patterns[43996] = 25'b10101011_11011010_10000101_1;
      patterns[43997] = 25'b10101011_11011011_10000110_1;
      patterns[43998] = 25'b10101011_11011100_10000111_1;
      patterns[43999] = 25'b10101011_11011101_10001000_1;
      patterns[44000] = 25'b10101011_11011110_10001001_1;
      patterns[44001] = 25'b10101011_11011111_10001010_1;
      patterns[44002] = 25'b10101011_11100000_10001011_1;
      patterns[44003] = 25'b10101011_11100001_10001100_1;
      patterns[44004] = 25'b10101011_11100010_10001101_1;
      patterns[44005] = 25'b10101011_11100011_10001110_1;
      patterns[44006] = 25'b10101011_11100100_10001111_1;
      patterns[44007] = 25'b10101011_11100101_10010000_1;
      patterns[44008] = 25'b10101011_11100110_10010001_1;
      patterns[44009] = 25'b10101011_11100111_10010010_1;
      patterns[44010] = 25'b10101011_11101000_10010011_1;
      patterns[44011] = 25'b10101011_11101001_10010100_1;
      patterns[44012] = 25'b10101011_11101010_10010101_1;
      patterns[44013] = 25'b10101011_11101011_10010110_1;
      patterns[44014] = 25'b10101011_11101100_10010111_1;
      patterns[44015] = 25'b10101011_11101101_10011000_1;
      patterns[44016] = 25'b10101011_11101110_10011001_1;
      patterns[44017] = 25'b10101011_11101111_10011010_1;
      patterns[44018] = 25'b10101011_11110000_10011011_1;
      patterns[44019] = 25'b10101011_11110001_10011100_1;
      patterns[44020] = 25'b10101011_11110010_10011101_1;
      patterns[44021] = 25'b10101011_11110011_10011110_1;
      patterns[44022] = 25'b10101011_11110100_10011111_1;
      patterns[44023] = 25'b10101011_11110101_10100000_1;
      patterns[44024] = 25'b10101011_11110110_10100001_1;
      patterns[44025] = 25'b10101011_11110111_10100010_1;
      patterns[44026] = 25'b10101011_11111000_10100011_1;
      patterns[44027] = 25'b10101011_11111001_10100100_1;
      patterns[44028] = 25'b10101011_11111010_10100101_1;
      patterns[44029] = 25'b10101011_11111011_10100110_1;
      patterns[44030] = 25'b10101011_11111100_10100111_1;
      patterns[44031] = 25'b10101011_11111101_10101000_1;
      patterns[44032] = 25'b10101011_11111110_10101001_1;
      patterns[44033] = 25'b10101011_11111111_10101010_1;
      patterns[44034] = 25'b10101100_00000000_10101100_0;
      patterns[44035] = 25'b10101100_00000001_10101101_0;
      patterns[44036] = 25'b10101100_00000010_10101110_0;
      patterns[44037] = 25'b10101100_00000011_10101111_0;
      patterns[44038] = 25'b10101100_00000100_10110000_0;
      patterns[44039] = 25'b10101100_00000101_10110001_0;
      patterns[44040] = 25'b10101100_00000110_10110010_0;
      patterns[44041] = 25'b10101100_00000111_10110011_0;
      patterns[44042] = 25'b10101100_00001000_10110100_0;
      patterns[44043] = 25'b10101100_00001001_10110101_0;
      patterns[44044] = 25'b10101100_00001010_10110110_0;
      patterns[44045] = 25'b10101100_00001011_10110111_0;
      patterns[44046] = 25'b10101100_00001100_10111000_0;
      patterns[44047] = 25'b10101100_00001101_10111001_0;
      patterns[44048] = 25'b10101100_00001110_10111010_0;
      patterns[44049] = 25'b10101100_00001111_10111011_0;
      patterns[44050] = 25'b10101100_00010000_10111100_0;
      patterns[44051] = 25'b10101100_00010001_10111101_0;
      patterns[44052] = 25'b10101100_00010010_10111110_0;
      patterns[44053] = 25'b10101100_00010011_10111111_0;
      patterns[44054] = 25'b10101100_00010100_11000000_0;
      patterns[44055] = 25'b10101100_00010101_11000001_0;
      patterns[44056] = 25'b10101100_00010110_11000010_0;
      patterns[44057] = 25'b10101100_00010111_11000011_0;
      patterns[44058] = 25'b10101100_00011000_11000100_0;
      patterns[44059] = 25'b10101100_00011001_11000101_0;
      patterns[44060] = 25'b10101100_00011010_11000110_0;
      patterns[44061] = 25'b10101100_00011011_11000111_0;
      patterns[44062] = 25'b10101100_00011100_11001000_0;
      patterns[44063] = 25'b10101100_00011101_11001001_0;
      patterns[44064] = 25'b10101100_00011110_11001010_0;
      patterns[44065] = 25'b10101100_00011111_11001011_0;
      patterns[44066] = 25'b10101100_00100000_11001100_0;
      patterns[44067] = 25'b10101100_00100001_11001101_0;
      patterns[44068] = 25'b10101100_00100010_11001110_0;
      patterns[44069] = 25'b10101100_00100011_11001111_0;
      patterns[44070] = 25'b10101100_00100100_11010000_0;
      patterns[44071] = 25'b10101100_00100101_11010001_0;
      patterns[44072] = 25'b10101100_00100110_11010010_0;
      patterns[44073] = 25'b10101100_00100111_11010011_0;
      patterns[44074] = 25'b10101100_00101000_11010100_0;
      patterns[44075] = 25'b10101100_00101001_11010101_0;
      patterns[44076] = 25'b10101100_00101010_11010110_0;
      patterns[44077] = 25'b10101100_00101011_11010111_0;
      patterns[44078] = 25'b10101100_00101100_11011000_0;
      patterns[44079] = 25'b10101100_00101101_11011001_0;
      patterns[44080] = 25'b10101100_00101110_11011010_0;
      patterns[44081] = 25'b10101100_00101111_11011011_0;
      patterns[44082] = 25'b10101100_00110000_11011100_0;
      patterns[44083] = 25'b10101100_00110001_11011101_0;
      patterns[44084] = 25'b10101100_00110010_11011110_0;
      patterns[44085] = 25'b10101100_00110011_11011111_0;
      patterns[44086] = 25'b10101100_00110100_11100000_0;
      patterns[44087] = 25'b10101100_00110101_11100001_0;
      patterns[44088] = 25'b10101100_00110110_11100010_0;
      patterns[44089] = 25'b10101100_00110111_11100011_0;
      patterns[44090] = 25'b10101100_00111000_11100100_0;
      patterns[44091] = 25'b10101100_00111001_11100101_0;
      patterns[44092] = 25'b10101100_00111010_11100110_0;
      patterns[44093] = 25'b10101100_00111011_11100111_0;
      patterns[44094] = 25'b10101100_00111100_11101000_0;
      patterns[44095] = 25'b10101100_00111101_11101001_0;
      patterns[44096] = 25'b10101100_00111110_11101010_0;
      patterns[44097] = 25'b10101100_00111111_11101011_0;
      patterns[44098] = 25'b10101100_01000000_11101100_0;
      patterns[44099] = 25'b10101100_01000001_11101101_0;
      patterns[44100] = 25'b10101100_01000010_11101110_0;
      patterns[44101] = 25'b10101100_01000011_11101111_0;
      patterns[44102] = 25'b10101100_01000100_11110000_0;
      patterns[44103] = 25'b10101100_01000101_11110001_0;
      patterns[44104] = 25'b10101100_01000110_11110010_0;
      patterns[44105] = 25'b10101100_01000111_11110011_0;
      patterns[44106] = 25'b10101100_01001000_11110100_0;
      patterns[44107] = 25'b10101100_01001001_11110101_0;
      patterns[44108] = 25'b10101100_01001010_11110110_0;
      patterns[44109] = 25'b10101100_01001011_11110111_0;
      patterns[44110] = 25'b10101100_01001100_11111000_0;
      patterns[44111] = 25'b10101100_01001101_11111001_0;
      patterns[44112] = 25'b10101100_01001110_11111010_0;
      patterns[44113] = 25'b10101100_01001111_11111011_0;
      patterns[44114] = 25'b10101100_01010000_11111100_0;
      patterns[44115] = 25'b10101100_01010001_11111101_0;
      patterns[44116] = 25'b10101100_01010010_11111110_0;
      patterns[44117] = 25'b10101100_01010011_11111111_0;
      patterns[44118] = 25'b10101100_01010100_00000000_1;
      patterns[44119] = 25'b10101100_01010101_00000001_1;
      patterns[44120] = 25'b10101100_01010110_00000010_1;
      patterns[44121] = 25'b10101100_01010111_00000011_1;
      patterns[44122] = 25'b10101100_01011000_00000100_1;
      patterns[44123] = 25'b10101100_01011001_00000101_1;
      patterns[44124] = 25'b10101100_01011010_00000110_1;
      patterns[44125] = 25'b10101100_01011011_00000111_1;
      patterns[44126] = 25'b10101100_01011100_00001000_1;
      patterns[44127] = 25'b10101100_01011101_00001001_1;
      patterns[44128] = 25'b10101100_01011110_00001010_1;
      patterns[44129] = 25'b10101100_01011111_00001011_1;
      patterns[44130] = 25'b10101100_01100000_00001100_1;
      patterns[44131] = 25'b10101100_01100001_00001101_1;
      patterns[44132] = 25'b10101100_01100010_00001110_1;
      patterns[44133] = 25'b10101100_01100011_00001111_1;
      patterns[44134] = 25'b10101100_01100100_00010000_1;
      patterns[44135] = 25'b10101100_01100101_00010001_1;
      patterns[44136] = 25'b10101100_01100110_00010010_1;
      patterns[44137] = 25'b10101100_01100111_00010011_1;
      patterns[44138] = 25'b10101100_01101000_00010100_1;
      patterns[44139] = 25'b10101100_01101001_00010101_1;
      patterns[44140] = 25'b10101100_01101010_00010110_1;
      patterns[44141] = 25'b10101100_01101011_00010111_1;
      patterns[44142] = 25'b10101100_01101100_00011000_1;
      patterns[44143] = 25'b10101100_01101101_00011001_1;
      patterns[44144] = 25'b10101100_01101110_00011010_1;
      patterns[44145] = 25'b10101100_01101111_00011011_1;
      patterns[44146] = 25'b10101100_01110000_00011100_1;
      patterns[44147] = 25'b10101100_01110001_00011101_1;
      patterns[44148] = 25'b10101100_01110010_00011110_1;
      patterns[44149] = 25'b10101100_01110011_00011111_1;
      patterns[44150] = 25'b10101100_01110100_00100000_1;
      patterns[44151] = 25'b10101100_01110101_00100001_1;
      patterns[44152] = 25'b10101100_01110110_00100010_1;
      patterns[44153] = 25'b10101100_01110111_00100011_1;
      patterns[44154] = 25'b10101100_01111000_00100100_1;
      patterns[44155] = 25'b10101100_01111001_00100101_1;
      patterns[44156] = 25'b10101100_01111010_00100110_1;
      patterns[44157] = 25'b10101100_01111011_00100111_1;
      patterns[44158] = 25'b10101100_01111100_00101000_1;
      patterns[44159] = 25'b10101100_01111101_00101001_1;
      patterns[44160] = 25'b10101100_01111110_00101010_1;
      patterns[44161] = 25'b10101100_01111111_00101011_1;
      patterns[44162] = 25'b10101100_10000000_00101100_1;
      patterns[44163] = 25'b10101100_10000001_00101101_1;
      patterns[44164] = 25'b10101100_10000010_00101110_1;
      patterns[44165] = 25'b10101100_10000011_00101111_1;
      patterns[44166] = 25'b10101100_10000100_00110000_1;
      patterns[44167] = 25'b10101100_10000101_00110001_1;
      patterns[44168] = 25'b10101100_10000110_00110010_1;
      patterns[44169] = 25'b10101100_10000111_00110011_1;
      patterns[44170] = 25'b10101100_10001000_00110100_1;
      patterns[44171] = 25'b10101100_10001001_00110101_1;
      patterns[44172] = 25'b10101100_10001010_00110110_1;
      patterns[44173] = 25'b10101100_10001011_00110111_1;
      patterns[44174] = 25'b10101100_10001100_00111000_1;
      patterns[44175] = 25'b10101100_10001101_00111001_1;
      patterns[44176] = 25'b10101100_10001110_00111010_1;
      patterns[44177] = 25'b10101100_10001111_00111011_1;
      patterns[44178] = 25'b10101100_10010000_00111100_1;
      patterns[44179] = 25'b10101100_10010001_00111101_1;
      patterns[44180] = 25'b10101100_10010010_00111110_1;
      patterns[44181] = 25'b10101100_10010011_00111111_1;
      patterns[44182] = 25'b10101100_10010100_01000000_1;
      patterns[44183] = 25'b10101100_10010101_01000001_1;
      patterns[44184] = 25'b10101100_10010110_01000010_1;
      patterns[44185] = 25'b10101100_10010111_01000011_1;
      patterns[44186] = 25'b10101100_10011000_01000100_1;
      patterns[44187] = 25'b10101100_10011001_01000101_1;
      patterns[44188] = 25'b10101100_10011010_01000110_1;
      patterns[44189] = 25'b10101100_10011011_01000111_1;
      patterns[44190] = 25'b10101100_10011100_01001000_1;
      patterns[44191] = 25'b10101100_10011101_01001001_1;
      patterns[44192] = 25'b10101100_10011110_01001010_1;
      patterns[44193] = 25'b10101100_10011111_01001011_1;
      patterns[44194] = 25'b10101100_10100000_01001100_1;
      patterns[44195] = 25'b10101100_10100001_01001101_1;
      patterns[44196] = 25'b10101100_10100010_01001110_1;
      patterns[44197] = 25'b10101100_10100011_01001111_1;
      patterns[44198] = 25'b10101100_10100100_01010000_1;
      patterns[44199] = 25'b10101100_10100101_01010001_1;
      patterns[44200] = 25'b10101100_10100110_01010010_1;
      patterns[44201] = 25'b10101100_10100111_01010011_1;
      patterns[44202] = 25'b10101100_10101000_01010100_1;
      patterns[44203] = 25'b10101100_10101001_01010101_1;
      patterns[44204] = 25'b10101100_10101010_01010110_1;
      patterns[44205] = 25'b10101100_10101011_01010111_1;
      patterns[44206] = 25'b10101100_10101100_01011000_1;
      patterns[44207] = 25'b10101100_10101101_01011001_1;
      patterns[44208] = 25'b10101100_10101110_01011010_1;
      patterns[44209] = 25'b10101100_10101111_01011011_1;
      patterns[44210] = 25'b10101100_10110000_01011100_1;
      patterns[44211] = 25'b10101100_10110001_01011101_1;
      patterns[44212] = 25'b10101100_10110010_01011110_1;
      patterns[44213] = 25'b10101100_10110011_01011111_1;
      patterns[44214] = 25'b10101100_10110100_01100000_1;
      patterns[44215] = 25'b10101100_10110101_01100001_1;
      patterns[44216] = 25'b10101100_10110110_01100010_1;
      patterns[44217] = 25'b10101100_10110111_01100011_1;
      patterns[44218] = 25'b10101100_10111000_01100100_1;
      patterns[44219] = 25'b10101100_10111001_01100101_1;
      patterns[44220] = 25'b10101100_10111010_01100110_1;
      patterns[44221] = 25'b10101100_10111011_01100111_1;
      patterns[44222] = 25'b10101100_10111100_01101000_1;
      patterns[44223] = 25'b10101100_10111101_01101001_1;
      patterns[44224] = 25'b10101100_10111110_01101010_1;
      patterns[44225] = 25'b10101100_10111111_01101011_1;
      patterns[44226] = 25'b10101100_11000000_01101100_1;
      patterns[44227] = 25'b10101100_11000001_01101101_1;
      patterns[44228] = 25'b10101100_11000010_01101110_1;
      patterns[44229] = 25'b10101100_11000011_01101111_1;
      patterns[44230] = 25'b10101100_11000100_01110000_1;
      patterns[44231] = 25'b10101100_11000101_01110001_1;
      patterns[44232] = 25'b10101100_11000110_01110010_1;
      patterns[44233] = 25'b10101100_11000111_01110011_1;
      patterns[44234] = 25'b10101100_11001000_01110100_1;
      patterns[44235] = 25'b10101100_11001001_01110101_1;
      patterns[44236] = 25'b10101100_11001010_01110110_1;
      patterns[44237] = 25'b10101100_11001011_01110111_1;
      patterns[44238] = 25'b10101100_11001100_01111000_1;
      patterns[44239] = 25'b10101100_11001101_01111001_1;
      patterns[44240] = 25'b10101100_11001110_01111010_1;
      patterns[44241] = 25'b10101100_11001111_01111011_1;
      patterns[44242] = 25'b10101100_11010000_01111100_1;
      patterns[44243] = 25'b10101100_11010001_01111101_1;
      patterns[44244] = 25'b10101100_11010010_01111110_1;
      patterns[44245] = 25'b10101100_11010011_01111111_1;
      patterns[44246] = 25'b10101100_11010100_10000000_1;
      patterns[44247] = 25'b10101100_11010101_10000001_1;
      patterns[44248] = 25'b10101100_11010110_10000010_1;
      patterns[44249] = 25'b10101100_11010111_10000011_1;
      patterns[44250] = 25'b10101100_11011000_10000100_1;
      patterns[44251] = 25'b10101100_11011001_10000101_1;
      patterns[44252] = 25'b10101100_11011010_10000110_1;
      patterns[44253] = 25'b10101100_11011011_10000111_1;
      patterns[44254] = 25'b10101100_11011100_10001000_1;
      patterns[44255] = 25'b10101100_11011101_10001001_1;
      patterns[44256] = 25'b10101100_11011110_10001010_1;
      patterns[44257] = 25'b10101100_11011111_10001011_1;
      patterns[44258] = 25'b10101100_11100000_10001100_1;
      patterns[44259] = 25'b10101100_11100001_10001101_1;
      patterns[44260] = 25'b10101100_11100010_10001110_1;
      patterns[44261] = 25'b10101100_11100011_10001111_1;
      patterns[44262] = 25'b10101100_11100100_10010000_1;
      patterns[44263] = 25'b10101100_11100101_10010001_1;
      patterns[44264] = 25'b10101100_11100110_10010010_1;
      patterns[44265] = 25'b10101100_11100111_10010011_1;
      patterns[44266] = 25'b10101100_11101000_10010100_1;
      patterns[44267] = 25'b10101100_11101001_10010101_1;
      patterns[44268] = 25'b10101100_11101010_10010110_1;
      patterns[44269] = 25'b10101100_11101011_10010111_1;
      patterns[44270] = 25'b10101100_11101100_10011000_1;
      patterns[44271] = 25'b10101100_11101101_10011001_1;
      patterns[44272] = 25'b10101100_11101110_10011010_1;
      patterns[44273] = 25'b10101100_11101111_10011011_1;
      patterns[44274] = 25'b10101100_11110000_10011100_1;
      patterns[44275] = 25'b10101100_11110001_10011101_1;
      patterns[44276] = 25'b10101100_11110010_10011110_1;
      patterns[44277] = 25'b10101100_11110011_10011111_1;
      patterns[44278] = 25'b10101100_11110100_10100000_1;
      patterns[44279] = 25'b10101100_11110101_10100001_1;
      patterns[44280] = 25'b10101100_11110110_10100010_1;
      patterns[44281] = 25'b10101100_11110111_10100011_1;
      patterns[44282] = 25'b10101100_11111000_10100100_1;
      patterns[44283] = 25'b10101100_11111001_10100101_1;
      patterns[44284] = 25'b10101100_11111010_10100110_1;
      patterns[44285] = 25'b10101100_11111011_10100111_1;
      patterns[44286] = 25'b10101100_11111100_10101000_1;
      patterns[44287] = 25'b10101100_11111101_10101001_1;
      patterns[44288] = 25'b10101100_11111110_10101010_1;
      patterns[44289] = 25'b10101100_11111111_10101011_1;
      patterns[44290] = 25'b10101101_00000000_10101101_0;
      patterns[44291] = 25'b10101101_00000001_10101110_0;
      patterns[44292] = 25'b10101101_00000010_10101111_0;
      patterns[44293] = 25'b10101101_00000011_10110000_0;
      patterns[44294] = 25'b10101101_00000100_10110001_0;
      patterns[44295] = 25'b10101101_00000101_10110010_0;
      patterns[44296] = 25'b10101101_00000110_10110011_0;
      patterns[44297] = 25'b10101101_00000111_10110100_0;
      patterns[44298] = 25'b10101101_00001000_10110101_0;
      patterns[44299] = 25'b10101101_00001001_10110110_0;
      patterns[44300] = 25'b10101101_00001010_10110111_0;
      patterns[44301] = 25'b10101101_00001011_10111000_0;
      patterns[44302] = 25'b10101101_00001100_10111001_0;
      patterns[44303] = 25'b10101101_00001101_10111010_0;
      patterns[44304] = 25'b10101101_00001110_10111011_0;
      patterns[44305] = 25'b10101101_00001111_10111100_0;
      patterns[44306] = 25'b10101101_00010000_10111101_0;
      patterns[44307] = 25'b10101101_00010001_10111110_0;
      patterns[44308] = 25'b10101101_00010010_10111111_0;
      patterns[44309] = 25'b10101101_00010011_11000000_0;
      patterns[44310] = 25'b10101101_00010100_11000001_0;
      patterns[44311] = 25'b10101101_00010101_11000010_0;
      patterns[44312] = 25'b10101101_00010110_11000011_0;
      patterns[44313] = 25'b10101101_00010111_11000100_0;
      patterns[44314] = 25'b10101101_00011000_11000101_0;
      patterns[44315] = 25'b10101101_00011001_11000110_0;
      patterns[44316] = 25'b10101101_00011010_11000111_0;
      patterns[44317] = 25'b10101101_00011011_11001000_0;
      patterns[44318] = 25'b10101101_00011100_11001001_0;
      patterns[44319] = 25'b10101101_00011101_11001010_0;
      patterns[44320] = 25'b10101101_00011110_11001011_0;
      patterns[44321] = 25'b10101101_00011111_11001100_0;
      patterns[44322] = 25'b10101101_00100000_11001101_0;
      patterns[44323] = 25'b10101101_00100001_11001110_0;
      patterns[44324] = 25'b10101101_00100010_11001111_0;
      patterns[44325] = 25'b10101101_00100011_11010000_0;
      patterns[44326] = 25'b10101101_00100100_11010001_0;
      patterns[44327] = 25'b10101101_00100101_11010010_0;
      patterns[44328] = 25'b10101101_00100110_11010011_0;
      patterns[44329] = 25'b10101101_00100111_11010100_0;
      patterns[44330] = 25'b10101101_00101000_11010101_0;
      patterns[44331] = 25'b10101101_00101001_11010110_0;
      patterns[44332] = 25'b10101101_00101010_11010111_0;
      patterns[44333] = 25'b10101101_00101011_11011000_0;
      patterns[44334] = 25'b10101101_00101100_11011001_0;
      patterns[44335] = 25'b10101101_00101101_11011010_0;
      patterns[44336] = 25'b10101101_00101110_11011011_0;
      patterns[44337] = 25'b10101101_00101111_11011100_0;
      patterns[44338] = 25'b10101101_00110000_11011101_0;
      patterns[44339] = 25'b10101101_00110001_11011110_0;
      patterns[44340] = 25'b10101101_00110010_11011111_0;
      patterns[44341] = 25'b10101101_00110011_11100000_0;
      patterns[44342] = 25'b10101101_00110100_11100001_0;
      patterns[44343] = 25'b10101101_00110101_11100010_0;
      patterns[44344] = 25'b10101101_00110110_11100011_0;
      patterns[44345] = 25'b10101101_00110111_11100100_0;
      patterns[44346] = 25'b10101101_00111000_11100101_0;
      patterns[44347] = 25'b10101101_00111001_11100110_0;
      patterns[44348] = 25'b10101101_00111010_11100111_0;
      patterns[44349] = 25'b10101101_00111011_11101000_0;
      patterns[44350] = 25'b10101101_00111100_11101001_0;
      patterns[44351] = 25'b10101101_00111101_11101010_0;
      patterns[44352] = 25'b10101101_00111110_11101011_0;
      patterns[44353] = 25'b10101101_00111111_11101100_0;
      patterns[44354] = 25'b10101101_01000000_11101101_0;
      patterns[44355] = 25'b10101101_01000001_11101110_0;
      patterns[44356] = 25'b10101101_01000010_11101111_0;
      patterns[44357] = 25'b10101101_01000011_11110000_0;
      patterns[44358] = 25'b10101101_01000100_11110001_0;
      patterns[44359] = 25'b10101101_01000101_11110010_0;
      patterns[44360] = 25'b10101101_01000110_11110011_0;
      patterns[44361] = 25'b10101101_01000111_11110100_0;
      patterns[44362] = 25'b10101101_01001000_11110101_0;
      patterns[44363] = 25'b10101101_01001001_11110110_0;
      patterns[44364] = 25'b10101101_01001010_11110111_0;
      patterns[44365] = 25'b10101101_01001011_11111000_0;
      patterns[44366] = 25'b10101101_01001100_11111001_0;
      patterns[44367] = 25'b10101101_01001101_11111010_0;
      patterns[44368] = 25'b10101101_01001110_11111011_0;
      patterns[44369] = 25'b10101101_01001111_11111100_0;
      patterns[44370] = 25'b10101101_01010000_11111101_0;
      patterns[44371] = 25'b10101101_01010001_11111110_0;
      patterns[44372] = 25'b10101101_01010010_11111111_0;
      patterns[44373] = 25'b10101101_01010011_00000000_1;
      patterns[44374] = 25'b10101101_01010100_00000001_1;
      patterns[44375] = 25'b10101101_01010101_00000010_1;
      patterns[44376] = 25'b10101101_01010110_00000011_1;
      patterns[44377] = 25'b10101101_01010111_00000100_1;
      patterns[44378] = 25'b10101101_01011000_00000101_1;
      patterns[44379] = 25'b10101101_01011001_00000110_1;
      patterns[44380] = 25'b10101101_01011010_00000111_1;
      patterns[44381] = 25'b10101101_01011011_00001000_1;
      patterns[44382] = 25'b10101101_01011100_00001001_1;
      patterns[44383] = 25'b10101101_01011101_00001010_1;
      patterns[44384] = 25'b10101101_01011110_00001011_1;
      patterns[44385] = 25'b10101101_01011111_00001100_1;
      patterns[44386] = 25'b10101101_01100000_00001101_1;
      patterns[44387] = 25'b10101101_01100001_00001110_1;
      patterns[44388] = 25'b10101101_01100010_00001111_1;
      patterns[44389] = 25'b10101101_01100011_00010000_1;
      patterns[44390] = 25'b10101101_01100100_00010001_1;
      patterns[44391] = 25'b10101101_01100101_00010010_1;
      patterns[44392] = 25'b10101101_01100110_00010011_1;
      patterns[44393] = 25'b10101101_01100111_00010100_1;
      patterns[44394] = 25'b10101101_01101000_00010101_1;
      patterns[44395] = 25'b10101101_01101001_00010110_1;
      patterns[44396] = 25'b10101101_01101010_00010111_1;
      patterns[44397] = 25'b10101101_01101011_00011000_1;
      patterns[44398] = 25'b10101101_01101100_00011001_1;
      patterns[44399] = 25'b10101101_01101101_00011010_1;
      patterns[44400] = 25'b10101101_01101110_00011011_1;
      patterns[44401] = 25'b10101101_01101111_00011100_1;
      patterns[44402] = 25'b10101101_01110000_00011101_1;
      patterns[44403] = 25'b10101101_01110001_00011110_1;
      patterns[44404] = 25'b10101101_01110010_00011111_1;
      patterns[44405] = 25'b10101101_01110011_00100000_1;
      patterns[44406] = 25'b10101101_01110100_00100001_1;
      patterns[44407] = 25'b10101101_01110101_00100010_1;
      patterns[44408] = 25'b10101101_01110110_00100011_1;
      patterns[44409] = 25'b10101101_01110111_00100100_1;
      patterns[44410] = 25'b10101101_01111000_00100101_1;
      patterns[44411] = 25'b10101101_01111001_00100110_1;
      patterns[44412] = 25'b10101101_01111010_00100111_1;
      patterns[44413] = 25'b10101101_01111011_00101000_1;
      patterns[44414] = 25'b10101101_01111100_00101001_1;
      patterns[44415] = 25'b10101101_01111101_00101010_1;
      patterns[44416] = 25'b10101101_01111110_00101011_1;
      patterns[44417] = 25'b10101101_01111111_00101100_1;
      patterns[44418] = 25'b10101101_10000000_00101101_1;
      patterns[44419] = 25'b10101101_10000001_00101110_1;
      patterns[44420] = 25'b10101101_10000010_00101111_1;
      patterns[44421] = 25'b10101101_10000011_00110000_1;
      patterns[44422] = 25'b10101101_10000100_00110001_1;
      patterns[44423] = 25'b10101101_10000101_00110010_1;
      patterns[44424] = 25'b10101101_10000110_00110011_1;
      patterns[44425] = 25'b10101101_10000111_00110100_1;
      patterns[44426] = 25'b10101101_10001000_00110101_1;
      patterns[44427] = 25'b10101101_10001001_00110110_1;
      patterns[44428] = 25'b10101101_10001010_00110111_1;
      patterns[44429] = 25'b10101101_10001011_00111000_1;
      patterns[44430] = 25'b10101101_10001100_00111001_1;
      patterns[44431] = 25'b10101101_10001101_00111010_1;
      patterns[44432] = 25'b10101101_10001110_00111011_1;
      patterns[44433] = 25'b10101101_10001111_00111100_1;
      patterns[44434] = 25'b10101101_10010000_00111101_1;
      patterns[44435] = 25'b10101101_10010001_00111110_1;
      patterns[44436] = 25'b10101101_10010010_00111111_1;
      patterns[44437] = 25'b10101101_10010011_01000000_1;
      patterns[44438] = 25'b10101101_10010100_01000001_1;
      patterns[44439] = 25'b10101101_10010101_01000010_1;
      patterns[44440] = 25'b10101101_10010110_01000011_1;
      patterns[44441] = 25'b10101101_10010111_01000100_1;
      patterns[44442] = 25'b10101101_10011000_01000101_1;
      patterns[44443] = 25'b10101101_10011001_01000110_1;
      patterns[44444] = 25'b10101101_10011010_01000111_1;
      patterns[44445] = 25'b10101101_10011011_01001000_1;
      patterns[44446] = 25'b10101101_10011100_01001001_1;
      patterns[44447] = 25'b10101101_10011101_01001010_1;
      patterns[44448] = 25'b10101101_10011110_01001011_1;
      patterns[44449] = 25'b10101101_10011111_01001100_1;
      patterns[44450] = 25'b10101101_10100000_01001101_1;
      patterns[44451] = 25'b10101101_10100001_01001110_1;
      patterns[44452] = 25'b10101101_10100010_01001111_1;
      patterns[44453] = 25'b10101101_10100011_01010000_1;
      patterns[44454] = 25'b10101101_10100100_01010001_1;
      patterns[44455] = 25'b10101101_10100101_01010010_1;
      patterns[44456] = 25'b10101101_10100110_01010011_1;
      patterns[44457] = 25'b10101101_10100111_01010100_1;
      patterns[44458] = 25'b10101101_10101000_01010101_1;
      patterns[44459] = 25'b10101101_10101001_01010110_1;
      patterns[44460] = 25'b10101101_10101010_01010111_1;
      patterns[44461] = 25'b10101101_10101011_01011000_1;
      patterns[44462] = 25'b10101101_10101100_01011001_1;
      patterns[44463] = 25'b10101101_10101101_01011010_1;
      patterns[44464] = 25'b10101101_10101110_01011011_1;
      patterns[44465] = 25'b10101101_10101111_01011100_1;
      patterns[44466] = 25'b10101101_10110000_01011101_1;
      patterns[44467] = 25'b10101101_10110001_01011110_1;
      patterns[44468] = 25'b10101101_10110010_01011111_1;
      patterns[44469] = 25'b10101101_10110011_01100000_1;
      patterns[44470] = 25'b10101101_10110100_01100001_1;
      patterns[44471] = 25'b10101101_10110101_01100010_1;
      patterns[44472] = 25'b10101101_10110110_01100011_1;
      patterns[44473] = 25'b10101101_10110111_01100100_1;
      patterns[44474] = 25'b10101101_10111000_01100101_1;
      patterns[44475] = 25'b10101101_10111001_01100110_1;
      patterns[44476] = 25'b10101101_10111010_01100111_1;
      patterns[44477] = 25'b10101101_10111011_01101000_1;
      patterns[44478] = 25'b10101101_10111100_01101001_1;
      patterns[44479] = 25'b10101101_10111101_01101010_1;
      patterns[44480] = 25'b10101101_10111110_01101011_1;
      patterns[44481] = 25'b10101101_10111111_01101100_1;
      patterns[44482] = 25'b10101101_11000000_01101101_1;
      patterns[44483] = 25'b10101101_11000001_01101110_1;
      patterns[44484] = 25'b10101101_11000010_01101111_1;
      patterns[44485] = 25'b10101101_11000011_01110000_1;
      patterns[44486] = 25'b10101101_11000100_01110001_1;
      patterns[44487] = 25'b10101101_11000101_01110010_1;
      patterns[44488] = 25'b10101101_11000110_01110011_1;
      patterns[44489] = 25'b10101101_11000111_01110100_1;
      patterns[44490] = 25'b10101101_11001000_01110101_1;
      patterns[44491] = 25'b10101101_11001001_01110110_1;
      patterns[44492] = 25'b10101101_11001010_01110111_1;
      patterns[44493] = 25'b10101101_11001011_01111000_1;
      patterns[44494] = 25'b10101101_11001100_01111001_1;
      patterns[44495] = 25'b10101101_11001101_01111010_1;
      patterns[44496] = 25'b10101101_11001110_01111011_1;
      patterns[44497] = 25'b10101101_11001111_01111100_1;
      patterns[44498] = 25'b10101101_11010000_01111101_1;
      patterns[44499] = 25'b10101101_11010001_01111110_1;
      patterns[44500] = 25'b10101101_11010010_01111111_1;
      patterns[44501] = 25'b10101101_11010011_10000000_1;
      patterns[44502] = 25'b10101101_11010100_10000001_1;
      patterns[44503] = 25'b10101101_11010101_10000010_1;
      patterns[44504] = 25'b10101101_11010110_10000011_1;
      patterns[44505] = 25'b10101101_11010111_10000100_1;
      patterns[44506] = 25'b10101101_11011000_10000101_1;
      patterns[44507] = 25'b10101101_11011001_10000110_1;
      patterns[44508] = 25'b10101101_11011010_10000111_1;
      patterns[44509] = 25'b10101101_11011011_10001000_1;
      patterns[44510] = 25'b10101101_11011100_10001001_1;
      patterns[44511] = 25'b10101101_11011101_10001010_1;
      patterns[44512] = 25'b10101101_11011110_10001011_1;
      patterns[44513] = 25'b10101101_11011111_10001100_1;
      patterns[44514] = 25'b10101101_11100000_10001101_1;
      patterns[44515] = 25'b10101101_11100001_10001110_1;
      patterns[44516] = 25'b10101101_11100010_10001111_1;
      patterns[44517] = 25'b10101101_11100011_10010000_1;
      patterns[44518] = 25'b10101101_11100100_10010001_1;
      patterns[44519] = 25'b10101101_11100101_10010010_1;
      patterns[44520] = 25'b10101101_11100110_10010011_1;
      patterns[44521] = 25'b10101101_11100111_10010100_1;
      patterns[44522] = 25'b10101101_11101000_10010101_1;
      patterns[44523] = 25'b10101101_11101001_10010110_1;
      patterns[44524] = 25'b10101101_11101010_10010111_1;
      patterns[44525] = 25'b10101101_11101011_10011000_1;
      patterns[44526] = 25'b10101101_11101100_10011001_1;
      patterns[44527] = 25'b10101101_11101101_10011010_1;
      patterns[44528] = 25'b10101101_11101110_10011011_1;
      patterns[44529] = 25'b10101101_11101111_10011100_1;
      patterns[44530] = 25'b10101101_11110000_10011101_1;
      patterns[44531] = 25'b10101101_11110001_10011110_1;
      patterns[44532] = 25'b10101101_11110010_10011111_1;
      patterns[44533] = 25'b10101101_11110011_10100000_1;
      patterns[44534] = 25'b10101101_11110100_10100001_1;
      patterns[44535] = 25'b10101101_11110101_10100010_1;
      patterns[44536] = 25'b10101101_11110110_10100011_1;
      patterns[44537] = 25'b10101101_11110111_10100100_1;
      patterns[44538] = 25'b10101101_11111000_10100101_1;
      patterns[44539] = 25'b10101101_11111001_10100110_1;
      patterns[44540] = 25'b10101101_11111010_10100111_1;
      patterns[44541] = 25'b10101101_11111011_10101000_1;
      patterns[44542] = 25'b10101101_11111100_10101001_1;
      patterns[44543] = 25'b10101101_11111101_10101010_1;
      patterns[44544] = 25'b10101101_11111110_10101011_1;
      patterns[44545] = 25'b10101101_11111111_10101100_1;
      patterns[44546] = 25'b10101110_00000000_10101110_0;
      patterns[44547] = 25'b10101110_00000001_10101111_0;
      patterns[44548] = 25'b10101110_00000010_10110000_0;
      patterns[44549] = 25'b10101110_00000011_10110001_0;
      patterns[44550] = 25'b10101110_00000100_10110010_0;
      patterns[44551] = 25'b10101110_00000101_10110011_0;
      patterns[44552] = 25'b10101110_00000110_10110100_0;
      patterns[44553] = 25'b10101110_00000111_10110101_0;
      patterns[44554] = 25'b10101110_00001000_10110110_0;
      patterns[44555] = 25'b10101110_00001001_10110111_0;
      patterns[44556] = 25'b10101110_00001010_10111000_0;
      patterns[44557] = 25'b10101110_00001011_10111001_0;
      patterns[44558] = 25'b10101110_00001100_10111010_0;
      patterns[44559] = 25'b10101110_00001101_10111011_0;
      patterns[44560] = 25'b10101110_00001110_10111100_0;
      patterns[44561] = 25'b10101110_00001111_10111101_0;
      patterns[44562] = 25'b10101110_00010000_10111110_0;
      patterns[44563] = 25'b10101110_00010001_10111111_0;
      patterns[44564] = 25'b10101110_00010010_11000000_0;
      patterns[44565] = 25'b10101110_00010011_11000001_0;
      patterns[44566] = 25'b10101110_00010100_11000010_0;
      patterns[44567] = 25'b10101110_00010101_11000011_0;
      patterns[44568] = 25'b10101110_00010110_11000100_0;
      patterns[44569] = 25'b10101110_00010111_11000101_0;
      patterns[44570] = 25'b10101110_00011000_11000110_0;
      patterns[44571] = 25'b10101110_00011001_11000111_0;
      patterns[44572] = 25'b10101110_00011010_11001000_0;
      patterns[44573] = 25'b10101110_00011011_11001001_0;
      patterns[44574] = 25'b10101110_00011100_11001010_0;
      patterns[44575] = 25'b10101110_00011101_11001011_0;
      patterns[44576] = 25'b10101110_00011110_11001100_0;
      patterns[44577] = 25'b10101110_00011111_11001101_0;
      patterns[44578] = 25'b10101110_00100000_11001110_0;
      patterns[44579] = 25'b10101110_00100001_11001111_0;
      patterns[44580] = 25'b10101110_00100010_11010000_0;
      patterns[44581] = 25'b10101110_00100011_11010001_0;
      patterns[44582] = 25'b10101110_00100100_11010010_0;
      patterns[44583] = 25'b10101110_00100101_11010011_0;
      patterns[44584] = 25'b10101110_00100110_11010100_0;
      patterns[44585] = 25'b10101110_00100111_11010101_0;
      patterns[44586] = 25'b10101110_00101000_11010110_0;
      patterns[44587] = 25'b10101110_00101001_11010111_0;
      patterns[44588] = 25'b10101110_00101010_11011000_0;
      patterns[44589] = 25'b10101110_00101011_11011001_0;
      patterns[44590] = 25'b10101110_00101100_11011010_0;
      patterns[44591] = 25'b10101110_00101101_11011011_0;
      patterns[44592] = 25'b10101110_00101110_11011100_0;
      patterns[44593] = 25'b10101110_00101111_11011101_0;
      patterns[44594] = 25'b10101110_00110000_11011110_0;
      patterns[44595] = 25'b10101110_00110001_11011111_0;
      patterns[44596] = 25'b10101110_00110010_11100000_0;
      patterns[44597] = 25'b10101110_00110011_11100001_0;
      patterns[44598] = 25'b10101110_00110100_11100010_0;
      patterns[44599] = 25'b10101110_00110101_11100011_0;
      patterns[44600] = 25'b10101110_00110110_11100100_0;
      patterns[44601] = 25'b10101110_00110111_11100101_0;
      patterns[44602] = 25'b10101110_00111000_11100110_0;
      patterns[44603] = 25'b10101110_00111001_11100111_0;
      patterns[44604] = 25'b10101110_00111010_11101000_0;
      patterns[44605] = 25'b10101110_00111011_11101001_0;
      patterns[44606] = 25'b10101110_00111100_11101010_0;
      patterns[44607] = 25'b10101110_00111101_11101011_0;
      patterns[44608] = 25'b10101110_00111110_11101100_0;
      patterns[44609] = 25'b10101110_00111111_11101101_0;
      patterns[44610] = 25'b10101110_01000000_11101110_0;
      patterns[44611] = 25'b10101110_01000001_11101111_0;
      patterns[44612] = 25'b10101110_01000010_11110000_0;
      patterns[44613] = 25'b10101110_01000011_11110001_0;
      patterns[44614] = 25'b10101110_01000100_11110010_0;
      patterns[44615] = 25'b10101110_01000101_11110011_0;
      patterns[44616] = 25'b10101110_01000110_11110100_0;
      patterns[44617] = 25'b10101110_01000111_11110101_0;
      patterns[44618] = 25'b10101110_01001000_11110110_0;
      patterns[44619] = 25'b10101110_01001001_11110111_0;
      patterns[44620] = 25'b10101110_01001010_11111000_0;
      patterns[44621] = 25'b10101110_01001011_11111001_0;
      patterns[44622] = 25'b10101110_01001100_11111010_0;
      patterns[44623] = 25'b10101110_01001101_11111011_0;
      patterns[44624] = 25'b10101110_01001110_11111100_0;
      patterns[44625] = 25'b10101110_01001111_11111101_0;
      patterns[44626] = 25'b10101110_01010000_11111110_0;
      patterns[44627] = 25'b10101110_01010001_11111111_0;
      patterns[44628] = 25'b10101110_01010010_00000000_1;
      patterns[44629] = 25'b10101110_01010011_00000001_1;
      patterns[44630] = 25'b10101110_01010100_00000010_1;
      patterns[44631] = 25'b10101110_01010101_00000011_1;
      patterns[44632] = 25'b10101110_01010110_00000100_1;
      patterns[44633] = 25'b10101110_01010111_00000101_1;
      patterns[44634] = 25'b10101110_01011000_00000110_1;
      patterns[44635] = 25'b10101110_01011001_00000111_1;
      patterns[44636] = 25'b10101110_01011010_00001000_1;
      patterns[44637] = 25'b10101110_01011011_00001001_1;
      patterns[44638] = 25'b10101110_01011100_00001010_1;
      patterns[44639] = 25'b10101110_01011101_00001011_1;
      patterns[44640] = 25'b10101110_01011110_00001100_1;
      patterns[44641] = 25'b10101110_01011111_00001101_1;
      patterns[44642] = 25'b10101110_01100000_00001110_1;
      patterns[44643] = 25'b10101110_01100001_00001111_1;
      patterns[44644] = 25'b10101110_01100010_00010000_1;
      patterns[44645] = 25'b10101110_01100011_00010001_1;
      patterns[44646] = 25'b10101110_01100100_00010010_1;
      patterns[44647] = 25'b10101110_01100101_00010011_1;
      patterns[44648] = 25'b10101110_01100110_00010100_1;
      patterns[44649] = 25'b10101110_01100111_00010101_1;
      patterns[44650] = 25'b10101110_01101000_00010110_1;
      patterns[44651] = 25'b10101110_01101001_00010111_1;
      patterns[44652] = 25'b10101110_01101010_00011000_1;
      patterns[44653] = 25'b10101110_01101011_00011001_1;
      patterns[44654] = 25'b10101110_01101100_00011010_1;
      patterns[44655] = 25'b10101110_01101101_00011011_1;
      patterns[44656] = 25'b10101110_01101110_00011100_1;
      patterns[44657] = 25'b10101110_01101111_00011101_1;
      patterns[44658] = 25'b10101110_01110000_00011110_1;
      patterns[44659] = 25'b10101110_01110001_00011111_1;
      patterns[44660] = 25'b10101110_01110010_00100000_1;
      patterns[44661] = 25'b10101110_01110011_00100001_1;
      patterns[44662] = 25'b10101110_01110100_00100010_1;
      patterns[44663] = 25'b10101110_01110101_00100011_1;
      patterns[44664] = 25'b10101110_01110110_00100100_1;
      patterns[44665] = 25'b10101110_01110111_00100101_1;
      patterns[44666] = 25'b10101110_01111000_00100110_1;
      patterns[44667] = 25'b10101110_01111001_00100111_1;
      patterns[44668] = 25'b10101110_01111010_00101000_1;
      patterns[44669] = 25'b10101110_01111011_00101001_1;
      patterns[44670] = 25'b10101110_01111100_00101010_1;
      patterns[44671] = 25'b10101110_01111101_00101011_1;
      patterns[44672] = 25'b10101110_01111110_00101100_1;
      patterns[44673] = 25'b10101110_01111111_00101101_1;
      patterns[44674] = 25'b10101110_10000000_00101110_1;
      patterns[44675] = 25'b10101110_10000001_00101111_1;
      patterns[44676] = 25'b10101110_10000010_00110000_1;
      patterns[44677] = 25'b10101110_10000011_00110001_1;
      patterns[44678] = 25'b10101110_10000100_00110010_1;
      patterns[44679] = 25'b10101110_10000101_00110011_1;
      patterns[44680] = 25'b10101110_10000110_00110100_1;
      patterns[44681] = 25'b10101110_10000111_00110101_1;
      patterns[44682] = 25'b10101110_10001000_00110110_1;
      patterns[44683] = 25'b10101110_10001001_00110111_1;
      patterns[44684] = 25'b10101110_10001010_00111000_1;
      patterns[44685] = 25'b10101110_10001011_00111001_1;
      patterns[44686] = 25'b10101110_10001100_00111010_1;
      patterns[44687] = 25'b10101110_10001101_00111011_1;
      patterns[44688] = 25'b10101110_10001110_00111100_1;
      patterns[44689] = 25'b10101110_10001111_00111101_1;
      patterns[44690] = 25'b10101110_10010000_00111110_1;
      patterns[44691] = 25'b10101110_10010001_00111111_1;
      patterns[44692] = 25'b10101110_10010010_01000000_1;
      patterns[44693] = 25'b10101110_10010011_01000001_1;
      patterns[44694] = 25'b10101110_10010100_01000010_1;
      patterns[44695] = 25'b10101110_10010101_01000011_1;
      patterns[44696] = 25'b10101110_10010110_01000100_1;
      patterns[44697] = 25'b10101110_10010111_01000101_1;
      patterns[44698] = 25'b10101110_10011000_01000110_1;
      patterns[44699] = 25'b10101110_10011001_01000111_1;
      patterns[44700] = 25'b10101110_10011010_01001000_1;
      patterns[44701] = 25'b10101110_10011011_01001001_1;
      patterns[44702] = 25'b10101110_10011100_01001010_1;
      patterns[44703] = 25'b10101110_10011101_01001011_1;
      patterns[44704] = 25'b10101110_10011110_01001100_1;
      patterns[44705] = 25'b10101110_10011111_01001101_1;
      patterns[44706] = 25'b10101110_10100000_01001110_1;
      patterns[44707] = 25'b10101110_10100001_01001111_1;
      patterns[44708] = 25'b10101110_10100010_01010000_1;
      patterns[44709] = 25'b10101110_10100011_01010001_1;
      patterns[44710] = 25'b10101110_10100100_01010010_1;
      patterns[44711] = 25'b10101110_10100101_01010011_1;
      patterns[44712] = 25'b10101110_10100110_01010100_1;
      patterns[44713] = 25'b10101110_10100111_01010101_1;
      patterns[44714] = 25'b10101110_10101000_01010110_1;
      patterns[44715] = 25'b10101110_10101001_01010111_1;
      patterns[44716] = 25'b10101110_10101010_01011000_1;
      patterns[44717] = 25'b10101110_10101011_01011001_1;
      patterns[44718] = 25'b10101110_10101100_01011010_1;
      patterns[44719] = 25'b10101110_10101101_01011011_1;
      patterns[44720] = 25'b10101110_10101110_01011100_1;
      patterns[44721] = 25'b10101110_10101111_01011101_1;
      patterns[44722] = 25'b10101110_10110000_01011110_1;
      patterns[44723] = 25'b10101110_10110001_01011111_1;
      patterns[44724] = 25'b10101110_10110010_01100000_1;
      patterns[44725] = 25'b10101110_10110011_01100001_1;
      patterns[44726] = 25'b10101110_10110100_01100010_1;
      patterns[44727] = 25'b10101110_10110101_01100011_1;
      patterns[44728] = 25'b10101110_10110110_01100100_1;
      patterns[44729] = 25'b10101110_10110111_01100101_1;
      patterns[44730] = 25'b10101110_10111000_01100110_1;
      patterns[44731] = 25'b10101110_10111001_01100111_1;
      patterns[44732] = 25'b10101110_10111010_01101000_1;
      patterns[44733] = 25'b10101110_10111011_01101001_1;
      patterns[44734] = 25'b10101110_10111100_01101010_1;
      patterns[44735] = 25'b10101110_10111101_01101011_1;
      patterns[44736] = 25'b10101110_10111110_01101100_1;
      patterns[44737] = 25'b10101110_10111111_01101101_1;
      patterns[44738] = 25'b10101110_11000000_01101110_1;
      patterns[44739] = 25'b10101110_11000001_01101111_1;
      patterns[44740] = 25'b10101110_11000010_01110000_1;
      patterns[44741] = 25'b10101110_11000011_01110001_1;
      patterns[44742] = 25'b10101110_11000100_01110010_1;
      patterns[44743] = 25'b10101110_11000101_01110011_1;
      patterns[44744] = 25'b10101110_11000110_01110100_1;
      patterns[44745] = 25'b10101110_11000111_01110101_1;
      patterns[44746] = 25'b10101110_11001000_01110110_1;
      patterns[44747] = 25'b10101110_11001001_01110111_1;
      patterns[44748] = 25'b10101110_11001010_01111000_1;
      patterns[44749] = 25'b10101110_11001011_01111001_1;
      patterns[44750] = 25'b10101110_11001100_01111010_1;
      patterns[44751] = 25'b10101110_11001101_01111011_1;
      patterns[44752] = 25'b10101110_11001110_01111100_1;
      patterns[44753] = 25'b10101110_11001111_01111101_1;
      patterns[44754] = 25'b10101110_11010000_01111110_1;
      patterns[44755] = 25'b10101110_11010001_01111111_1;
      patterns[44756] = 25'b10101110_11010010_10000000_1;
      patterns[44757] = 25'b10101110_11010011_10000001_1;
      patterns[44758] = 25'b10101110_11010100_10000010_1;
      patterns[44759] = 25'b10101110_11010101_10000011_1;
      patterns[44760] = 25'b10101110_11010110_10000100_1;
      patterns[44761] = 25'b10101110_11010111_10000101_1;
      patterns[44762] = 25'b10101110_11011000_10000110_1;
      patterns[44763] = 25'b10101110_11011001_10000111_1;
      patterns[44764] = 25'b10101110_11011010_10001000_1;
      patterns[44765] = 25'b10101110_11011011_10001001_1;
      patterns[44766] = 25'b10101110_11011100_10001010_1;
      patterns[44767] = 25'b10101110_11011101_10001011_1;
      patterns[44768] = 25'b10101110_11011110_10001100_1;
      patterns[44769] = 25'b10101110_11011111_10001101_1;
      patterns[44770] = 25'b10101110_11100000_10001110_1;
      patterns[44771] = 25'b10101110_11100001_10001111_1;
      patterns[44772] = 25'b10101110_11100010_10010000_1;
      patterns[44773] = 25'b10101110_11100011_10010001_1;
      patterns[44774] = 25'b10101110_11100100_10010010_1;
      patterns[44775] = 25'b10101110_11100101_10010011_1;
      patterns[44776] = 25'b10101110_11100110_10010100_1;
      patterns[44777] = 25'b10101110_11100111_10010101_1;
      patterns[44778] = 25'b10101110_11101000_10010110_1;
      patterns[44779] = 25'b10101110_11101001_10010111_1;
      patterns[44780] = 25'b10101110_11101010_10011000_1;
      patterns[44781] = 25'b10101110_11101011_10011001_1;
      patterns[44782] = 25'b10101110_11101100_10011010_1;
      patterns[44783] = 25'b10101110_11101101_10011011_1;
      patterns[44784] = 25'b10101110_11101110_10011100_1;
      patterns[44785] = 25'b10101110_11101111_10011101_1;
      patterns[44786] = 25'b10101110_11110000_10011110_1;
      patterns[44787] = 25'b10101110_11110001_10011111_1;
      patterns[44788] = 25'b10101110_11110010_10100000_1;
      patterns[44789] = 25'b10101110_11110011_10100001_1;
      patterns[44790] = 25'b10101110_11110100_10100010_1;
      patterns[44791] = 25'b10101110_11110101_10100011_1;
      patterns[44792] = 25'b10101110_11110110_10100100_1;
      patterns[44793] = 25'b10101110_11110111_10100101_1;
      patterns[44794] = 25'b10101110_11111000_10100110_1;
      patterns[44795] = 25'b10101110_11111001_10100111_1;
      patterns[44796] = 25'b10101110_11111010_10101000_1;
      patterns[44797] = 25'b10101110_11111011_10101001_1;
      patterns[44798] = 25'b10101110_11111100_10101010_1;
      patterns[44799] = 25'b10101110_11111101_10101011_1;
      patterns[44800] = 25'b10101110_11111110_10101100_1;
      patterns[44801] = 25'b10101110_11111111_10101101_1;
      patterns[44802] = 25'b10101111_00000000_10101111_0;
      patterns[44803] = 25'b10101111_00000001_10110000_0;
      patterns[44804] = 25'b10101111_00000010_10110001_0;
      patterns[44805] = 25'b10101111_00000011_10110010_0;
      patterns[44806] = 25'b10101111_00000100_10110011_0;
      patterns[44807] = 25'b10101111_00000101_10110100_0;
      patterns[44808] = 25'b10101111_00000110_10110101_0;
      patterns[44809] = 25'b10101111_00000111_10110110_0;
      patterns[44810] = 25'b10101111_00001000_10110111_0;
      patterns[44811] = 25'b10101111_00001001_10111000_0;
      patterns[44812] = 25'b10101111_00001010_10111001_0;
      patterns[44813] = 25'b10101111_00001011_10111010_0;
      patterns[44814] = 25'b10101111_00001100_10111011_0;
      patterns[44815] = 25'b10101111_00001101_10111100_0;
      patterns[44816] = 25'b10101111_00001110_10111101_0;
      patterns[44817] = 25'b10101111_00001111_10111110_0;
      patterns[44818] = 25'b10101111_00010000_10111111_0;
      patterns[44819] = 25'b10101111_00010001_11000000_0;
      patterns[44820] = 25'b10101111_00010010_11000001_0;
      patterns[44821] = 25'b10101111_00010011_11000010_0;
      patterns[44822] = 25'b10101111_00010100_11000011_0;
      patterns[44823] = 25'b10101111_00010101_11000100_0;
      patterns[44824] = 25'b10101111_00010110_11000101_0;
      patterns[44825] = 25'b10101111_00010111_11000110_0;
      patterns[44826] = 25'b10101111_00011000_11000111_0;
      patterns[44827] = 25'b10101111_00011001_11001000_0;
      patterns[44828] = 25'b10101111_00011010_11001001_0;
      patterns[44829] = 25'b10101111_00011011_11001010_0;
      patterns[44830] = 25'b10101111_00011100_11001011_0;
      patterns[44831] = 25'b10101111_00011101_11001100_0;
      patterns[44832] = 25'b10101111_00011110_11001101_0;
      patterns[44833] = 25'b10101111_00011111_11001110_0;
      patterns[44834] = 25'b10101111_00100000_11001111_0;
      patterns[44835] = 25'b10101111_00100001_11010000_0;
      patterns[44836] = 25'b10101111_00100010_11010001_0;
      patterns[44837] = 25'b10101111_00100011_11010010_0;
      patterns[44838] = 25'b10101111_00100100_11010011_0;
      patterns[44839] = 25'b10101111_00100101_11010100_0;
      patterns[44840] = 25'b10101111_00100110_11010101_0;
      patterns[44841] = 25'b10101111_00100111_11010110_0;
      patterns[44842] = 25'b10101111_00101000_11010111_0;
      patterns[44843] = 25'b10101111_00101001_11011000_0;
      patterns[44844] = 25'b10101111_00101010_11011001_0;
      patterns[44845] = 25'b10101111_00101011_11011010_0;
      patterns[44846] = 25'b10101111_00101100_11011011_0;
      patterns[44847] = 25'b10101111_00101101_11011100_0;
      patterns[44848] = 25'b10101111_00101110_11011101_0;
      patterns[44849] = 25'b10101111_00101111_11011110_0;
      patterns[44850] = 25'b10101111_00110000_11011111_0;
      patterns[44851] = 25'b10101111_00110001_11100000_0;
      patterns[44852] = 25'b10101111_00110010_11100001_0;
      patterns[44853] = 25'b10101111_00110011_11100010_0;
      patterns[44854] = 25'b10101111_00110100_11100011_0;
      patterns[44855] = 25'b10101111_00110101_11100100_0;
      patterns[44856] = 25'b10101111_00110110_11100101_0;
      patterns[44857] = 25'b10101111_00110111_11100110_0;
      patterns[44858] = 25'b10101111_00111000_11100111_0;
      patterns[44859] = 25'b10101111_00111001_11101000_0;
      patterns[44860] = 25'b10101111_00111010_11101001_0;
      patterns[44861] = 25'b10101111_00111011_11101010_0;
      patterns[44862] = 25'b10101111_00111100_11101011_0;
      patterns[44863] = 25'b10101111_00111101_11101100_0;
      patterns[44864] = 25'b10101111_00111110_11101101_0;
      patterns[44865] = 25'b10101111_00111111_11101110_0;
      patterns[44866] = 25'b10101111_01000000_11101111_0;
      patterns[44867] = 25'b10101111_01000001_11110000_0;
      patterns[44868] = 25'b10101111_01000010_11110001_0;
      patterns[44869] = 25'b10101111_01000011_11110010_0;
      patterns[44870] = 25'b10101111_01000100_11110011_0;
      patterns[44871] = 25'b10101111_01000101_11110100_0;
      patterns[44872] = 25'b10101111_01000110_11110101_0;
      patterns[44873] = 25'b10101111_01000111_11110110_0;
      patterns[44874] = 25'b10101111_01001000_11110111_0;
      patterns[44875] = 25'b10101111_01001001_11111000_0;
      patterns[44876] = 25'b10101111_01001010_11111001_0;
      patterns[44877] = 25'b10101111_01001011_11111010_0;
      patterns[44878] = 25'b10101111_01001100_11111011_0;
      patterns[44879] = 25'b10101111_01001101_11111100_0;
      patterns[44880] = 25'b10101111_01001110_11111101_0;
      patterns[44881] = 25'b10101111_01001111_11111110_0;
      patterns[44882] = 25'b10101111_01010000_11111111_0;
      patterns[44883] = 25'b10101111_01010001_00000000_1;
      patterns[44884] = 25'b10101111_01010010_00000001_1;
      patterns[44885] = 25'b10101111_01010011_00000010_1;
      patterns[44886] = 25'b10101111_01010100_00000011_1;
      patterns[44887] = 25'b10101111_01010101_00000100_1;
      patterns[44888] = 25'b10101111_01010110_00000101_1;
      patterns[44889] = 25'b10101111_01010111_00000110_1;
      patterns[44890] = 25'b10101111_01011000_00000111_1;
      patterns[44891] = 25'b10101111_01011001_00001000_1;
      patterns[44892] = 25'b10101111_01011010_00001001_1;
      patterns[44893] = 25'b10101111_01011011_00001010_1;
      patterns[44894] = 25'b10101111_01011100_00001011_1;
      patterns[44895] = 25'b10101111_01011101_00001100_1;
      patterns[44896] = 25'b10101111_01011110_00001101_1;
      patterns[44897] = 25'b10101111_01011111_00001110_1;
      patterns[44898] = 25'b10101111_01100000_00001111_1;
      patterns[44899] = 25'b10101111_01100001_00010000_1;
      patterns[44900] = 25'b10101111_01100010_00010001_1;
      patterns[44901] = 25'b10101111_01100011_00010010_1;
      patterns[44902] = 25'b10101111_01100100_00010011_1;
      patterns[44903] = 25'b10101111_01100101_00010100_1;
      patterns[44904] = 25'b10101111_01100110_00010101_1;
      patterns[44905] = 25'b10101111_01100111_00010110_1;
      patterns[44906] = 25'b10101111_01101000_00010111_1;
      patterns[44907] = 25'b10101111_01101001_00011000_1;
      patterns[44908] = 25'b10101111_01101010_00011001_1;
      patterns[44909] = 25'b10101111_01101011_00011010_1;
      patterns[44910] = 25'b10101111_01101100_00011011_1;
      patterns[44911] = 25'b10101111_01101101_00011100_1;
      patterns[44912] = 25'b10101111_01101110_00011101_1;
      patterns[44913] = 25'b10101111_01101111_00011110_1;
      patterns[44914] = 25'b10101111_01110000_00011111_1;
      patterns[44915] = 25'b10101111_01110001_00100000_1;
      patterns[44916] = 25'b10101111_01110010_00100001_1;
      patterns[44917] = 25'b10101111_01110011_00100010_1;
      patterns[44918] = 25'b10101111_01110100_00100011_1;
      patterns[44919] = 25'b10101111_01110101_00100100_1;
      patterns[44920] = 25'b10101111_01110110_00100101_1;
      patterns[44921] = 25'b10101111_01110111_00100110_1;
      patterns[44922] = 25'b10101111_01111000_00100111_1;
      patterns[44923] = 25'b10101111_01111001_00101000_1;
      patterns[44924] = 25'b10101111_01111010_00101001_1;
      patterns[44925] = 25'b10101111_01111011_00101010_1;
      patterns[44926] = 25'b10101111_01111100_00101011_1;
      patterns[44927] = 25'b10101111_01111101_00101100_1;
      patterns[44928] = 25'b10101111_01111110_00101101_1;
      patterns[44929] = 25'b10101111_01111111_00101110_1;
      patterns[44930] = 25'b10101111_10000000_00101111_1;
      patterns[44931] = 25'b10101111_10000001_00110000_1;
      patterns[44932] = 25'b10101111_10000010_00110001_1;
      patterns[44933] = 25'b10101111_10000011_00110010_1;
      patterns[44934] = 25'b10101111_10000100_00110011_1;
      patterns[44935] = 25'b10101111_10000101_00110100_1;
      patterns[44936] = 25'b10101111_10000110_00110101_1;
      patterns[44937] = 25'b10101111_10000111_00110110_1;
      patterns[44938] = 25'b10101111_10001000_00110111_1;
      patterns[44939] = 25'b10101111_10001001_00111000_1;
      patterns[44940] = 25'b10101111_10001010_00111001_1;
      patterns[44941] = 25'b10101111_10001011_00111010_1;
      patterns[44942] = 25'b10101111_10001100_00111011_1;
      patterns[44943] = 25'b10101111_10001101_00111100_1;
      patterns[44944] = 25'b10101111_10001110_00111101_1;
      patterns[44945] = 25'b10101111_10001111_00111110_1;
      patterns[44946] = 25'b10101111_10010000_00111111_1;
      patterns[44947] = 25'b10101111_10010001_01000000_1;
      patterns[44948] = 25'b10101111_10010010_01000001_1;
      patterns[44949] = 25'b10101111_10010011_01000010_1;
      patterns[44950] = 25'b10101111_10010100_01000011_1;
      patterns[44951] = 25'b10101111_10010101_01000100_1;
      patterns[44952] = 25'b10101111_10010110_01000101_1;
      patterns[44953] = 25'b10101111_10010111_01000110_1;
      patterns[44954] = 25'b10101111_10011000_01000111_1;
      patterns[44955] = 25'b10101111_10011001_01001000_1;
      patterns[44956] = 25'b10101111_10011010_01001001_1;
      patterns[44957] = 25'b10101111_10011011_01001010_1;
      patterns[44958] = 25'b10101111_10011100_01001011_1;
      patterns[44959] = 25'b10101111_10011101_01001100_1;
      patterns[44960] = 25'b10101111_10011110_01001101_1;
      patterns[44961] = 25'b10101111_10011111_01001110_1;
      patterns[44962] = 25'b10101111_10100000_01001111_1;
      patterns[44963] = 25'b10101111_10100001_01010000_1;
      patterns[44964] = 25'b10101111_10100010_01010001_1;
      patterns[44965] = 25'b10101111_10100011_01010010_1;
      patterns[44966] = 25'b10101111_10100100_01010011_1;
      patterns[44967] = 25'b10101111_10100101_01010100_1;
      patterns[44968] = 25'b10101111_10100110_01010101_1;
      patterns[44969] = 25'b10101111_10100111_01010110_1;
      patterns[44970] = 25'b10101111_10101000_01010111_1;
      patterns[44971] = 25'b10101111_10101001_01011000_1;
      patterns[44972] = 25'b10101111_10101010_01011001_1;
      patterns[44973] = 25'b10101111_10101011_01011010_1;
      patterns[44974] = 25'b10101111_10101100_01011011_1;
      patterns[44975] = 25'b10101111_10101101_01011100_1;
      patterns[44976] = 25'b10101111_10101110_01011101_1;
      patterns[44977] = 25'b10101111_10101111_01011110_1;
      patterns[44978] = 25'b10101111_10110000_01011111_1;
      patterns[44979] = 25'b10101111_10110001_01100000_1;
      patterns[44980] = 25'b10101111_10110010_01100001_1;
      patterns[44981] = 25'b10101111_10110011_01100010_1;
      patterns[44982] = 25'b10101111_10110100_01100011_1;
      patterns[44983] = 25'b10101111_10110101_01100100_1;
      patterns[44984] = 25'b10101111_10110110_01100101_1;
      patterns[44985] = 25'b10101111_10110111_01100110_1;
      patterns[44986] = 25'b10101111_10111000_01100111_1;
      patterns[44987] = 25'b10101111_10111001_01101000_1;
      patterns[44988] = 25'b10101111_10111010_01101001_1;
      patterns[44989] = 25'b10101111_10111011_01101010_1;
      patterns[44990] = 25'b10101111_10111100_01101011_1;
      patterns[44991] = 25'b10101111_10111101_01101100_1;
      patterns[44992] = 25'b10101111_10111110_01101101_1;
      patterns[44993] = 25'b10101111_10111111_01101110_1;
      patterns[44994] = 25'b10101111_11000000_01101111_1;
      patterns[44995] = 25'b10101111_11000001_01110000_1;
      patterns[44996] = 25'b10101111_11000010_01110001_1;
      patterns[44997] = 25'b10101111_11000011_01110010_1;
      patterns[44998] = 25'b10101111_11000100_01110011_1;
      patterns[44999] = 25'b10101111_11000101_01110100_1;
      patterns[45000] = 25'b10101111_11000110_01110101_1;
      patterns[45001] = 25'b10101111_11000111_01110110_1;
      patterns[45002] = 25'b10101111_11001000_01110111_1;
      patterns[45003] = 25'b10101111_11001001_01111000_1;
      patterns[45004] = 25'b10101111_11001010_01111001_1;
      patterns[45005] = 25'b10101111_11001011_01111010_1;
      patterns[45006] = 25'b10101111_11001100_01111011_1;
      patterns[45007] = 25'b10101111_11001101_01111100_1;
      patterns[45008] = 25'b10101111_11001110_01111101_1;
      patterns[45009] = 25'b10101111_11001111_01111110_1;
      patterns[45010] = 25'b10101111_11010000_01111111_1;
      patterns[45011] = 25'b10101111_11010001_10000000_1;
      patterns[45012] = 25'b10101111_11010010_10000001_1;
      patterns[45013] = 25'b10101111_11010011_10000010_1;
      patterns[45014] = 25'b10101111_11010100_10000011_1;
      patterns[45015] = 25'b10101111_11010101_10000100_1;
      patterns[45016] = 25'b10101111_11010110_10000101_1;
      patterns[45017] = 25'b10101111_11010111_10000110_1;
      patterns[45018] = 25'b10101111_11011000_10000111_1;
      patterns[45019] = 25'b10101111_11011001_10001000_1;
      patterns[45020] = 25'b10101111_11011010_10001001_1;
      patterns[45021] = 25'b10101111_11011011_10001010_1;
      patterns[45022] = 25'b10101111_11011100_10001011_1;
      patterns[45023] = 25'b10101111_11011101_10001100_1;
      patterns[45024] = 25'b10101111_11011110_10001101_1;
      patterns[45025] = 25'b10101111_11011111_10001110_1;
      patterns[45026] = 25'b10101111_11100000_10001111_1;
      patterns[45027] = 25'b10101111_11100001_10010000_1;
      patterns[45028] = 25'b10101111_11100010_10010001_1;
      patterns[45029] = 25'b10101111_11100011_10010010_1;
      patterns[45030] = 25'b10101111_11100100_10010011_1;
      patterns[45031] = 25'b10101111_11100101_10010100_1;
      patterns[45032] = 25'b10101111_11100110_10010101_1;
      patterns[45033] = 25'b10101111_11100111_10010110_1;
      patterns[45034] = 25'b10101111_11101000_10010111_1;
      patterns[45035] = 25'b10101111_11101001_10011000_1;
      patterns[45036] = 25'b10101111_11101010_10011001_1;
      patterns[45037] = 25'b10101111_11101011_10011010_1;
      patterns[45038] = 25'b10101111_11101100_10011011_1;
      patterns[45039] = 25'b10101111_11101101_10011100_1;
      patterns[45040] = 25'b10101111_11101110_10011101_1;
      patterns[45041] = 25'b10101111_11101111_10011110_1;
      patterns[45042] = 25'b10101111_11110000_10011111_1;
      patterns[45043] = 25'b10101111_11110001_10100000_1;
      patterns[45044] = 25'b10101111_11110010_10100001_1;
      patterns[45045] = 25'b10101111_11110011_10100010_1;
      patterns[45046] = 25'b10101111_11110100_10100011_1;
      patterns[45047] = 25'b10101111_11110101_10100100_1;
      patterns[45048] = 25'b10101111_11110110_10100101_1;
      patterns[45049] = 25'b10101111_11110111_10100110_1;
      patterns[45050] = 25'b10101111_11111000_10100111_1;
      patterns[45051] = 25'b10101111_11111001_10101000_1;
      patterns[45052] = 25'b10101111_11111010_10101001_1;
      patterns[45053] = 25'b10101111_11111011_10101010_1;
      patterns[45054] = 25'b10101111_11111100_10101011_1;
      patterns[45055] = 25'b10101111_11111101_10101100_1;
      patterns[45056] = 25'b10101111_11111110_10101101_1;
      patterns[45057] = 25'b10101111_11111111_10101110_1;
      patterns[45058] = 25'b10110000_00000000_10110000_0;
      patterns[45059] = 25'b10110000_00000001_10110001_0;
      patterns[45060] = 25'b10110000_00000010_10110010_0;
      patterns[45061] = 25'b10110000_00000011_10110011_0;
      patterns[45062] = 25'b10110000_00000100_10110100_0;
      patterns[45063] = 25'b10110000_00000101_10110101_0;
      patterns[45064] = 25'b10110000_00000110_10110110_0;
      patterns[45065] = 25'b10110000_00000111_10110111_0;
      patterns[45066] = 25'b10110000_00001000_10111000_0;
      patterns[45067] = 25'b10110000_00001001_10111001_0;
      patterns[45068] = 25'b10110000_00001010_10111010_0;
      patterns[45069] = 25'b10110000_00001011_10111011_0;
      patterns[45070] = 25'b10110000_00001100_10111100_0;
      patterns[45071] = 25'b10110000_00001101_10111101_0;
      patterns[45072] = 25'b10110000_00001110_10111110_0;
      patterns[45073] = 25'b10110000_00001111_10111111_0;
      patterns[45074] = 25'b10110000_00010000_11000000_0;
      patterns[45075] = 25'b10110000_00010001_11000001_0;
      patterns[45076] = 25'b10110000_00010010_11000010_0;
      patterns[45077] = 25'b10110000_00010011_11000011_0;
      patterns[45078] = 25'b10110000_00010100_11000100_0;
      patterns[45079] = 25'b10110000_00010101_11000101_0;
      patterns[45080] = 25'b10110000_00010110_11000110_0;
      patterns[45081] = 25'b10110000_00010111_11000111_0;
      patterns[45082] = 25'b10110000_00011000_11001000_0;
      patterns[45083] = 25'b10110000_00011001_11001001_0;
      patterns[45084] = 25'b10110000_00011010_11001010_0;
      patterns[45085] = 25'b10110000_00011011_11001011_0;
      patterns[45086] = 25'b10110000_00011100_11001100_0;
      patterns[45087] = 25'b10110000_00011101_11001101_0;
      patterns[45088] = 25'b10110000_00011110_11001110_0;
      patterns[45089] = 25'b10110000_00011111_11001111_0;
      patterns[45090] = 25'b10110000_00100000_11010000_0;
      patterns[45091] = 25'b10110000_00100001_11010001_0;
      patterns[45092] = 25'b10110000_00100010_11010010_0;
      patterns[45093] = 25'b10110000_00100011_11010011_0;
      patterns[45094] = 25'b10110000_00100100_11010100_0;
      patterns[45095] = 25'b10110000_00100101_11010101_0;
      patterns[45096] = 25'b10110000_00100110_11010110_0;
      patterns[45097] = 25'b10110000_00100111_11010111_0;
      patterns[45098] = 25'b10110000_00101000_11011000_0;
      patterns[45099] = 25'b10110000_00101001_11011001_0;
      patterns[45100] = 25'b10110000_00101010_11011010_0;
      patterns[45101] = 25'b10110000_00101011_11011011_0;
      patterns[45102] = 25'b10110000_00101100_11011100_0;
      patterns[45103] = 25'b10110000_00101101_11011101_0;
      patterns[45104] = 25'b10110000_00101110_11011110_0;
      patterns[45105] = 25'b10110000_00101111_11011111_0;
      patterns[45106] = 25'b10110000_00110000_11100000_0;
      patterns[45107] = 25'b10110000_00110001_11100001_0;
      patterns[45108] = 25'b10110000_00110010_11100010_0;
      patterns[45109] = 25'b10110000_00110011_11100011_0;
      patterns[45110] = 25'b10110000_00110100_11100100_0;
      patterns[45111] = 25'b10110000_00110101_11100101_0;
      patterns[45112] = 25'b10110000_00110110_11100110_0;
      patterns[45113] = 25'b10110000_00110111_11100111_0;
      patterns[45114] = 25'b10110000_00111000_11101000_0;
      patterns[45115] = 25'b10110000_00111001_11101001_0;
      patterns[45116] = 25'b10110000_00111010_11101010_0;
      patterns[45117] = 25'b10110000_00111011_11101011_0;
      patterns[45118] = 25'b10110000_00111100_11101100_0;
      patterns[45119] = 25'b10110000_00111101_11101101_0;
      patterns[45120] = 25'b10110000_00111110_11101110_0;
      patterns[45121] = 25'b10110000_00111111_11101111_0;
      patterns[45122] = 25'b10110000_01000000_11110000_0;
      patterns[45123] = 25'b10110000_01000001_11110001_0;
      patterns[45124] = 25'b10110000_01000010_11110010_0;
      patterns[45125] = 25'b10110000_01000011_11110011_0;
      patterns[45126] = 25'b10110000_01000100_11110100_0;
      patterns[45127] = 25'b10110000_01000101_11110101_0;
      patterns[45128] = 25'b10110000_01000110_11110110_0;
      patterns[45129] = 25'b10110000_01000111_11110111_0;
      patterns[45130] = 25'b10110000_01001000_11111000_0;
      patterns[45131] = 25'b10110000_01001001_11111001_0;
      patterns[45132] = 25'b10110000_01001010_11111010_0;
      patterns[45133] = 25'b10110000_01001011_11111011_0;
      patterns[45134] = 25'b10110000_01001100_11111100_0;
      patterns[45135] = 25'b10110000_01001101_11111101_0;
      patterns[45136] = 25'b10110000_01001110_11111110_0;
      patterns[45137] = 25'b10110000_01001111_11111111_0;
      patterns[45138] = 25'b10110000_01010000_00000000_1;
      patterns[45139] = 25'b10110000_01010001_00000001_1;
      patterns[45140] = 25'b10110000_01010010_00000010_1;
      patterns[45141] = 25'b10110000_01010011_00000011_1;
      patterns[45142] = 25'b10110000_01010100_00000100_1;
      patterns[45143] = 25'b10110000_01010101_00000101_1;
      patterns[45144] = 25'b10110000_01010110_00000110_1;
      patterns[45145] = 25'b10110000_01010111_00000111_1;
      patterns[45146] = 25'b10110000_01011000_00001000_1;
      patterns[45147] = 25'b10110000_01011001_00001001_1;
      patterns[45148] = 25'b10110000_01011010_00001010_1;
      patterns[45149] = 25'b10110000_01011011_00001011_1;
      patterns[45150] = 25'b10110000_01011100_00001100_1;
      patterns[45151] = 25'b10110000_01011101_00001101_1;
      patterns[45152] = 25'b10110000_01011110_00001110_1;
      patterns[45153] = 25'b10110000_01011111_00001111_1;
      patterns[45154] = 25'b10110000_01100000_00010000_1;
      patterns[45155] = 25'b10110000_01100001_00010001_1;
      patterns[45156] = 25'b10110000_01100010_00010010_1;
      patterns[45157] = 25'b10110000_01100011_00010011_1;
      patterns[45158] = 25'b10110000_01100100_00010100_1;
      patterns[45159] = 25'b10110000_01100101_00010101_1;
      patterns[45160] = 25'b10110000_01100110_00010110_1;
      patterns[45161] = 25'b10110000_01100111_00010111_1;
      patterns[45162] = 25'b10110000_01101000_00011000_1;
      patterns[45163] = 25'b10110000_01101001_00011001_1;
      patterns[45164] = 25'b10110000_01101010_00011010_1;
      patterns[45165] = 25'b10110000_01101011_00011011_1;
      patterns[45166] = 25'b10110000_01101100_00011100_1;
      patterns[45167] = 25'b10110000_01101101_00011101_1;
      patterns[45168] = 25'b10110000_01101110_00011110_1;
      patterns[45169] = 25'b10110000_01101111_00011111_1;
      patterns[45170] = 25'b10110000_01110000_00100000_1;
      patterns[45171] = 25'b10110000_01110001_00100001_1;
      patterns[45172] = 25'b10110000_01110010_00100010_1;
      patterns[45173] = 25'b10110000_01110011_00100011_1;
      patterns[45174] = 25'b10110000_01110100_00100100_1;
      patterns[45175] = 25'b10110000_01110101_00100101_1;
      patterns[45176] = 25'b10110000_01110110_00100110_1;
      patterns[45177] = 25'b10110000_01110111_00100111_1;
      patterns[45178] = 25'b10110000_01111000_00101000_1;
      patterns[45179] = 25'b10110000_01111001_00101001_1;
      patterns[45180] = 25'b10110000_01111010_00101010_1;
      patterns[45181] = 25'b10110000_01111011_00101011_1;
      patterns[45182] = 25'b10110000_01111100_00101100_1;
      patterns[45183] = 25'b10110000_01111101_00101101_1;
      patterns[45184] = 25'b10110000_01111110_00101110_1;
      patterns[45185] = 25'b10110000_01111111_00101111_1;
      patterns[45186] = 25'b10110000_10000000_00110000_1;
      patterns[45187] = 25'b10110000_10000001_00110001_1;
      patterns[45188] = 25'b10110000_10000010_00110010_1;
      patterns[45189] = 25'b10110000_10000011_00110011_1;
      patterns[45190] = 25'b10110000_10000100_00110100_1;
      patterns[45191] = 25'b10110000_10000101_00110101_1;
      patterns[45192] = 25'b10110000_10000110_00110110_1;
      patterns[45193] = 25'b10110000_10000111_00110111_1;
      patterns[45194] = 25'b10110000_10001000_00111000_1;
      patterns[45195] = 25'b10110000_10001001_00111001_1;
      patterns[45196] = 25'b10110000_10001010_00111010_1;
      patterns[45197] = 25'b10110000_10001011_00111011_1;
      patterns[45198] = 25'b10110000_10001100_00111100_1;
      patterns[45199] = 25'b10110000_10001101_00111101_1;
      patterns[45200] = 25'b10110000_10001110_00111110_1;
      patterns[45201] = 25'b10110000_10001111_00111111_1;
      patterns[45202] = 25'b10110000_10010000_01000000_1;
      patterns[45203] = 25'b10110000_10010001_01000001_1;
      patterns[45204] = 25'b10110000_10010010_01000010_1;
      patterns[45205] = 25'b10110000_10010011_01000011_1;
      patterns[45206] = 25'b10110000_10010100_01000100_1;
      patterns[45207] = 25'b10110000_10010101_01000101_1;
      patterns[45208] = 25'b10110000_10010110_01000110_1;
      patterns[45209] = 25'b10110000_10010111_01000111_1;
      patterns[45210] = 25'b10110000_10011000_01001000_1;
      patterns[45211] = 25'b10110000_10011001_01001001_1;
      patterns[45212] = 25'b10110000_10011010_01001010_1;
      patterns[45213] = 25'b10110000_10011011_01001011_1;
      patterns[45214] = 25'b10110000_10011100_01001100_1;
      patterns[45215] = 25'b10110000_10011101_01001101_1;
      patterns[45216] = 25'b10110000_10011110_01001110_1;
      patterns[45217] = 25'b10110000_10011111_01001111_1;
      patterns[45218] = 25'b10110000_10100000_01010000_1;
      patterns[45219] = 25'b10110000_10100001_01010001_1;
      patterns[45220] = 25'b10110000_10100010_01010010_1;
      patterns[45221] = 25'b10110000_10100011_01010011_1;
      patterns[45222] = 25'b10110000_10100100_01010100_1;
      patterns[45223] = 25'b10110000_10100101_01010101_1;
      patterns[45224] = 25'b10110000_10100110_01010110_1;
      patterns[45225] = 25'b10110000_10100111_01010111_1;
      patterns[45226] = 25'b10110000_10101000_01011000_1;
      patterns[45227] = 25'b10110000_10101001_01011001_1;
      patterns[45228] = 25'b10110000_10101010_01011010_1;
      patterns[45229] = 25'b10110000_10101011_01011011_1;
      patterns[45230] = 25'b10110000_10101100_01011100_1;
      patterns[45231] = 25'b10110000_10101101_01011101_1;
      patterns[45232] = 25'b10110000_10101110_01011110_1;
      patterns[45233] = 25'b10110000_10101111_01011111_1;
      patterns[45234] = 25'b10110000_10110000_01100000_1;
      patterns[45235] = 25'b10110000_10110001_01100001_1;
      patterns[45236] = 25'b10110000_10110010_01100010_1;
      patterns[45237] = 25'b10110000_10110011_01100011_1;
      patterns[45238] = 25'b10110000_10110100_01100100_1;
      patterns[45239] = 25'b10110000_10110101_01100101_1;
      patterns[45240] = 25'b10110000_10110110_01100110_1;
      patterns[45241] = 25'b10110000_10110111_01100111_1;
      patterns[45242] = 25'b10110000_10111000_01101000_1;
      patterns[45243] = 25'b10110000_10111001_01101001_1;
      patterns[45244] = 25'b10110000_10111010_01101010_1;
      patterns[45245] = 25'b10110000_10111011_01101011_1;
      patterns[45246] = 25'b10110000_10111100_01101100_1;
      patterns[45247] = 25'b10110000_10111101_01101101_1;
      patterns[45248] = 25'b10110000_10111110_01101110_1;
      patterns[45249] = 25'b10110000_10111111_01101111_1;
      patterns[45250] = 25'b10110000_11000000_01110000_1;
      patterns[45251] = 25'b10110000_11000001_01110001_1;
      patterns[45252] = 25'b10110000_11000010_01110010_1;
      patterns[45253] = 25'b10110000_11000011_01110011_1;
      patterns[45254] = 25'b10110000_11000100_01110100_1;
      patterns[45255] = 25'b10110000_11000101_01110101_1;
      patterns[45256] = 25'b10110000_11000110_01110110_1;
      patterns[45257] = 25'b10110000_11000111_01110111_1;
      patterns[45258] = 25'b10110000_11001000_01111000_1;
      patterns[45259] = 25'b10110000_11001001_01111001_1;
      patterns[45260] = 25'b10110000_11001010_01111010_1;
      patterns[45261] = 25'b10110000_11001011_01111011_1;
      patterns[45262] = 25'b10110000_11001100_01111100_1;
      patterns[45263] = 25'b10110000_11001101_01111101_1;
      patterns[45264] = 25'b10110000_11001110_01111110_1;
      patterns[45265] = 25'b10110000_11001111_01111111_1;
      patterns[45266] = 25'b10110000_11010000_10000000_1;
      patterns[45267] = 25'b10110000_11010001_10000001_1;
      patterns[45268] = 25'b10110000_11010010_10000010_1;
      patterns[45269] = 25'b10110000_11010011_10000011_1;
      patterns[45270] = 25'b10110000_11010100_10000100_1;
      patterns[45271] = 25'b10110000_11010101_10000101_1;
      patterns[45272] = 25'b10110000_11010110_10000110_1;
      patterns[45273] = 25'b10110000_11010111_10000111_1;
      patterns[45274] = 25'b10110000_11011000_10001000_1;
      patterns[45275] = 25'b10110000_11011001_10001001_1;
      patterns[45276] = 25'b10110000_11011010_10001010_1;
      patterns[45277] = 25'b10110000_11011011_10001011_1;
      patterns[45278] = 25'b10110000_11011100_10001100_1;
      patterns[45279] = 25'b10110000_11011101_10001101_1;
      patterns[45280] = 25'b10110000_11011110_10001110_1;
      patterns[45281] = 25'b10110000_11011111_10001111_1;
      patterns[45282] = 25'b10110000_11100000_10010000_1;
      patterns[45283] = 25'b10110000_11100001_10010001_1;
      patterns[45284] = 25'b10110000_11100010_10010010_1;
      patterns[45285] = 25'b10110000_11100011_10010011_1;
      patterns[45286] = 25'b10110000_11100100_10010100_1;
      patterns[45287] = 25'b10110000_11100101_10010101_1;
      patterns[45288] = 25'b10110000_11100110_10010110_1;
      patterns[45289] = 25'b10110000_11100111_10010111_1;
      patterns[45290] = 25'b10110000_11101000_10011000_1;
      patterns[45291] = 25'b10110000_11101001_10011001_1;
      patterns[45292] = 25'b10110000_11101010_10011010_1;
      patterns[45293] = 25'b10110000_11101011_10011011_1;
      patterns[45294] = 25'b10110000_11101100_10011100_1;
      patterns[45295] = 25'b10110000_11101101_10011101_1;
      patterns[45296] = 25'b10110000_11101110_10011110_1;
      patterns[45297] = 25'b10110000_11101111_10011111_1;
      patterns[45298] = 25'b10110000_11110000_10100000_1;
      patterns[45299] = 25'b10110000_11110001_10100001_1;
      patterns[45300] = 25'b10110000_11110010_10100010_1;
      patterns[45301] = 25'b10110000_11110011_10100011_1;
      patterns[45302] = 25'b10110000_11110100_10100100_1;
      patterns[45303] = 25'b10110000_11110101_10100101_1;
      patterns[45304] = 25'b10110000_11110110_10100110_1;
      patterns[45305] = 25'b10110000_11110111_10100111_1;
      patterns[45306] = 25'b10110000_11111000_10101000_1;
      patterns[45307] = 25'b10110000_11111001_10101001_1;
      patterns[45308] = 25'b10110000_11111010_10101010_1;
      patterns[45309] = 25'b10110000_11111011_10101011_1;
      patterns[45310] = 25'b10110000_11111100_10101100_1;
      patterns[45311] = 25'b10110000_11111101_10101101_1;
      patterns[45312] = 25'b10110000_11111110_10101110_1;
      patterns[45313] = 25'b10110000_11111111_10101111_1;
      patterns[45314] = 25'b10110001_00000000_10110001_0;
      patterns[45315] = 25'b10110001_00000001_10110010_0;
      patterns[45316] = 25'b10110001_00000010_10110011_0;
      patterns[45317] = 25'b10110001_00000011_10110100_0;
      patterns[45318] = 25'b10110001_00000100_10110101_0;
      patterns[45319] = 25'b10110001_00000101_10110110_0;
      patterns[45320] = 25'b10110001_00000110_10110111_0;
      patterns[45321] = 25'b10110001_00000111_10111000_0;
      patterns[45322] = 25'b10110001_00001000_10111001_0;
      patterns[45323] = 25'b10110001_00001001_10111010_0;
      patterns[45324] = 25'b10110001_00001010_10111011_0;
      patterns[45325] = 25'b10110001_00001011_10111100_0;
      patterns[45326] = 25'b10110001_00001100_10111101_0;
      patterns[45327] = 25'b10110001_00001101_10111110_0;
      patterns[45328] = 25'b10110001_00001110_10111111_0;
      patterns[45329] = 25'b10110001_00001111_11000000_0;
      patterns[45330] = 25'b10110001_00010000_11000001_0;
      patterns[45331] = 25'b10110001_00010001_11000010_0;
      patterns[45332] = 25'b10110001_00010010_11000011_0;
      patterns[45333] = 25'b10110001_00010011_11000100_0;
      patterns[45334] = 25'b10110001_00010100_11000101_0;
      patterns[45335] = 25'b10110001_00010101_11000110_0;
      patterns[45336] = 25'b10110001_00010110_11000111_0;
      patterns[45337] = 25'b10110001_00010111_11001000_0;
      patterns[45338] = 25'b10110001_00011000_11001001_0;
      patterns[45339] = 25'b10110001_00011001_11001010_0;
      patterns[45340] = 25'b10110001_00011010_11001011_0;
      patterns[45341] = 25'b10110001_00011011_11001100_0;
      patterns[45342] = 25'b10110001_00011100_11001101_0;
      patterns[45343] = 25'b10110001_00011101_11001110_0;
      patterns[45344] = 25'b10110001_00011110_11001111_0;
      patterns[45345] = 25'b10110001_00011111_11010000_0;
      patterns[45346] = 25'b10110001_00100000_11010001_0;
      patterns[45347] = 25'b10110001_00100001_11010010_0;
      patterns[45348] = 25'b10110001_00100010_11010011_0;
      patterns[45349] = 25'b10110001_00100011_11010100_0;
      patterns[45350] = 25'b10110001_00100100_11010101_0;
      patterns[45351] = 25'b10110001_00100101_11010110_0;
      patterns[45352] = 25'b10110001_00100110_11010111_0;
      patterns[45353] = 25'b10110001_00100111_11011000_0;
      patterns[45354] = 25'b10110001_00101000_11011001_0;
      patterns[45355] = 25'b10110001_00101001_11011010_0;
      patterns[45356] = 25'b10110001_00101010_11011011_0;
      patterns[45357] = 25'b10110001_00101011_11011100_0;
      patterns[45358] = 25'b10110001_00101100_11011101_0;
      patterns[45359] = 25'b10110001_00101101_11011110_0;
      patterns[45360] = 25'b10110001_00101110_11011111_0;
      patterns[45361] = 25'b10110001_00101111_11100000_0;
      patterns[45362] = 25'b10110001_00110000_11100001_0;
      patterns[45363] = 25'b10110001_00110001_11100010_0;
      patterns[45364] = 25'b10110001_00110010_11100011_0;
      patterns[45365] = 25'b10110001_00110011_11100100_0;
      patterns[45366] = 25'b10110001_00110100_11100101_0;
      patterns[45367] = 25'b10110001_00110101_11100110_0;
      patterns[45368] = 25'b10110001_00110110_11100111_0;
      patterns[45369] = 25'b10110001_00110111_11101000_0;
      patterns[45370] = 25'b10110001_00111000_11101001_0;
      patterns[45371] = 25'b10110001_00111001_11101010_0;
      patterns[45372] = 25'b10110001_00111010_11101011_0;
      patterns[45373] = 25'b10110001_00111011_11101100_0;
      patterns[45374] = 25'b10110001_00111100_11101101_0;
      patterns[45375] = 25'b10110001_00111101_11101110_0;
      patterns[45376] = 25'b10110001_00111110_11101111_0;
      patterns[45377] = 25'b10110001_00111111_11110000_0;
      patterns[45378] = 25'b10110001_01000000_11110001_0;
      patterns[45379] = 25'b10110001_01000001_11110010_0;
      patterns[45380] = 25'b10110001_01000010_11110011_0;
      patterns[45381] = 25'b10110001_01000011_11110100_0;
      patterns[45382] = 25'b10110001_01000100_11110101_0;
      patterns[45383] = 25'b10110001_01000101_11110110_0;
      patterns[45384] = 25'b10110001_01000110_11110111_0;
      patterns[45385] = 25'b10110001_01000111_11111000_0;
      patterns[45386] = 25'b10110001_01001000_11111001_0;
      patterns[45387] = 25'b10110001_01001001_11111010_0;
      patterns[45388] = 25'b10110001_01001010_11111011_0;
      patterns[45389] = 25'b10110001_01001011_11111100_0;
      patterns[45390] = 25'b10110001_01001100_11111101_0;
      patterns[45391] = 25'b10110001_01001101_11111110_0;
      patterns[45392] = 25'b10110001_01001110_11111111_0;
      patterns[45393] = 25'b10110001_01001111_00000000_1;
      patterns[45394] = 25'b10110001_01010000_00000001_1;
      patterns[45395] = 25'b10110001_01010001_00000010_1;
      patterns[45396] = 25'b10110001_01010010_00000011_1;
      patterns[45397] = 25'b10110001_01010011_00000100_1;
      patterns[45398] = 25'b10110001_01010100_00000101_1;
      patterns[45399] = 25'b10110001_01010101_00000110_1;
      patterns[45400] = 25'b10110001_01010110_00000111_1;
      patterns[45401] = 25'b10110001_01010111_00001000_1;
      patterns[45402] = 25'b10110001_01011000_00001001_1;
      patterns[45403] = 25'b10110001_01011001_00001010_1;
      patterns[45404] = 25'b10110001_01011010_00001011_1;
      patterns[45405] = 25'b10110001_01011011_00001100_1;
      patterns[45406] = 25'b10110001_01011100_00001101_1;
      patterns[45407] = 25'b10110001_01011101_00001110_1;
      patterns[45408] = 25'b10110001_01011110_00001111_1;
      patterns[45409] = 25'b10110001_01011111_00010000_1;
      patterns[45410] = 25'b10110001_01100000_00010001_1;
      patterns[45411] = 25'b10110001_01100001_00010010_1;
      patterns[45412] = 25'b10110001_01100010_00010011_1;
      patterns[45413] = 25'b10110001_01100011_00010100_1;
      patterns[45414] = 25'b10110001_01100100_00010101_1;
      patterns[45415] = 25'b10110001_01100101_00010110_1;
      patterns[45416] = 25'b10110001_01100110_00010111_1;
      patterns[45417] = 25'b10110001_01100111_00011000_1;
      patterns[45418] = 25'b10110001_01101000_00011001_1;
      patterns[45419] = 25'b10110001_01101001_00011010_1;
      patterns[45420] = 25'b10110001_01101010_00011011_1;
      patterns[45421] = 25'b10110001_01101011_00011100_1;
      patterns[45422] = 25'b10110001_01101100_00011101_1;
      patterns[45423] = 25'b10110001_01101101_00011110_1;
      patterns[45424] = 25'b10110001_01101110_00011111_1;
      patterns[45425] = 25'b10110001_01101111_00100000_1;
      patterns[45426] = 25'b10110001_01110000_00100001_1;
      patterns[45427] = 25'b10110001_01110001_00100010_1;
      patterns[45428] = 25'b10110001_01110010_00100011_1;
      patterns[45429] = 25'b10110001_01110011_00100100_1;
      patterns[45430] = 25'b10110001_01110100_00100101_1;
      patterns[45431] = 25'b10110001_01110101_00100110_1;
      patterns[45432] = 25'b10110001_01110110_00100111_1;
      patterns[45433] = 25'b10110001_01110111_00101000_1;
      patterns[45434] = 25'b10110001_01111000_00101001_1;
      patterns[45435] = 25'b10110001_01111001_00101010_1;
      patterns[45436] = 25'b10110001_01111010_00101011_1;
      patterns[45437] = 25'b10110001_01111011_00101100_1;
      patterns[45438] = 25'b10110001_01111100_00101101_1;
      patterns[45439] = 25'b10110001_01111101_00101110_1;
      patterns[45440] = 25'b10110001_01111110_00101111_1;
      patterns[45441] = 25'b10110001_01111111_00110000_1;
      patterns[45442] = 25'b10110001_10000000_00110001_1;
      patterns[45443] = 25'b10110001_10000001_00110010_1;
      patterns[45444] = 25'b10110001_10000010_00110011_1;
      patterns[45445] = 25'b10110001_10000011_00110100_1;
      patterns[45446] = 25'b10110001_10000100_00110101_1;
      patterns[45447] = 25'b10110001_10000101_00110110_1;
      patterns[45448] = 25'b10110001_10000110_00110111_1;
      patterns[45449] = 25'b10110001_10000111_00111000_1;
      patterns[45450] = 25'b10110001_10001000_00111001_1;
      patterns[45451] = 25'b10110001_10001001_00111010_1;
      patterns[45452] = 25'b10110001_10001010_00111011_1;
      patterns[45453] = 25'b10110001_10001011_00111100_1;
      patterns[45454] = 25'b10110001_10001100_00111101_1;
      patterns[45455] = 25'b10110001_10001101_00111110_1;
      patterns[45456] = 25'b10110001_10001110_00111111_1;
      patterns[45457] = 25'b10110001_10001111_01000000_1;
      patterns[45458] = 25'b10110001_10010000_01000001_1;
      patterns[45459] = 25'b10110001_10010001_01000010_1;
      patterns[45460] = 25'b10110001_10010010_01000011_1;
      patterns[45461] = 25'b10110001_10010011_01000100_1;
      patterns[45462] = 25'b10110001_10010100_01000101_1;
      patterns[45463] = 25'b10110001_10010101_01000110_1;
      patterns[45464] = 25'b10110001_10010110_01000111_1;
      patterns[45465] = 25'b10110001_10010111_01001000_1;
      patterns[45466] = 25'b10110001_10011000_01001001_1;
      patterns[45467] = 25'b10110001_10011001_01001010_1;
      patterns[45468] = 25'b10110001_10011010_01001011_1;
      patterns[45469] = 25'b10110001_10011011_01001100_1;
      patterns[45470] = 25'b10110001_10011100_01001101_1;
      patterns[45471] = 25'b10110001_10011101_01001110_1;
      patterns[45472] = 25'b10110001_10011110_01001111_1;
      patterns[45473] = 25'b10110001_10011111_01010000_1;
      patterns[45474] = 25'b10110001_10100000_01010001_1;
      patterns[45475] = 25'b10110001_10100001_01010010_1;
      patterns[45476] = 25'b10110001_10100010_01010011_1;
      patterns[45477] = 25'b10110001_10100011_01010100_1;
      patterns[45478] = 25'b10110001_10100100_01010101_1;
      patterns[45479] = 25'b10110001_10100101_01010110_1;
      patterns[45480] = 25'b10110001_10100110_01010111_1;
      patterns[45481] = 25'b10110001_10100111_01011000_1;
      patterns[45482] = 25'b10110001_10101000_01011001_1;
      patterns[45483] = 25'b10110001_10101001_01011010_1;
      patterns[45484] = 25'b10110001_10101010_01011011_1;
      patterns[45485] = 25'b10110001_10101011_01011100_1;
      patterns[45486] = 25'b10110001_10101100_01011101_1;
      patterns[45487] = 25'b10110001_10101101_01011110_1;
      patterns[45488] = 25'b10110001_10101110_01011111_1;
      patterns[45489] = 25'b10110001_10101111_01100000_1;
      patterns[45490] = 25'b10110001_10110000_01100001_1;
      patterns[45491] = 25'b10110001_10110001_01100010_1;
      patterns[45492] = 25'b10110001_10110010_01100011_1;
      patterns[45493] = 25'b10110001_10110011_01100100_1;
      patterns[45494] = 25'b10110001_10110100_01100101_1;
      patterns[45495] = 25'b10110001_10110101_01100110_1;
      patterns[45496] = 25'b10110001_10110110_01100111_1;
      patterns[45497] = 25'b10110001_10110111_01101000_1;
      patterns[45498] = 25'b10110001_10111000_01101001_1;
      patterns[45499] = 25'b10110001_10111001_01101010_1;
      patterns[45500] = 25'b10110001_10111010_01101011_1;
      patterns[45501] = 25'b10110001_10111011_01101100_1;
      patterns[45502] = 25'b10110001_10111100_01101101_1;
      patterns[45503] = 25'b10110001_10111101_01101110_1;
      patterns[45504] = 25'b10110001_10111110_01101111_1;
      patterns[45505] = 25'b10110001_10111111_01110000_1;
      patterns[45506] = 25'b10110001_11000000_01110001_1;
      patterns[45507] = 25'b10110001_11000001_01110010_1;
      patterns[45508] = 25'b10110001_11000010_01110011_1;
      patterns[45509] = 25'b10110001_11000011_01110100_1;
      patterns[45510] = 25'b10110001_11000100_01110101_1;
      patterns[45511] = 25'b10110001_11000101_01110110_1;
      patterns[45512] = 25'b10110001_11000110_01110111_1;
      patterns[45513] = 25'b10110001_11000111_01111000_1;
      patterns[45514] = 25'b10110001_11001000_01111001_1;
      patterns[45515] = 25'b10110001_11001001_01111010_1;
      patterns[45516] = 25'b10110001_11001010_01111011_1;
      patterns[45517] = 25'b10110001_11001011_01111100_1;
      patterns[45518] = 25'b10110001_11001100_01111101_1;
      patterns[45519] = 25'b10110001_11001101_01111110_1;
      patterns[45520] = 25'b10110001_11001110_01111111_1;
      patterns[45521] = 25'b10110001_11001111_10000000_1;
      patterns[45522] = 25'b10110001_11010000_10000001_1;
      patterns[45523] = 25'b10110001_11010001_10000010_1;
      patterns[45524] = 25'b10110001_11010010_10000011_1;
      patterns[45525] = 25'b10110001_11010011_10000100_1;
      patterns[45526] = 25'b10110001_11010100_10000101_1;
      patterns[45527] = 25'b10110001_11010101_10000110_1;
      patterns[45528] = 25'b10110001_11010110_10000111_1;
      patterns[45529] = 25'b10110001_11010111_10001000_1;
      patterns[45530] = 25'b10110001_11011000_10001001_1;
      patterns[45531] = 25'b10110001_11011001_10001010_1;
      patterns[45532] = 25'b10110001_11011010_10001011_1;
      patterns[45533] = 25'b10110001_11011011_10001100_1;
      patterns[45534] = 25'b10110001_11011100_10001101_1;
      patterns[45535] = 25'b10110001_11011101_10001110_1;
      patterns[45536] = 25'b10110001_11011110_10001111_1;
      patterns[45537] = 25'b10110001_11011111_10010000_1;
      patterns[45538] = 25'b10110001_11100000_10010001_1;
      patterns[45539] = 25'b10110001_11100001_10010010_1;
      patterns[45540] = 25'b10110001_11100010_10010011_1;
      patterns[45541] = 25'b10110001_11100011_10010100_1;
      patterns[45542] = 25'b10110001_11100100_10010101_1;
      patterns[45543] = 25'b10110001_11100101_10010110_1;
      patterns[45544] = 25'b10110001_11100110_10010111_1;
      patterns[45545] = 25'b10110001_11100111_10011000_1;
      patterns[45546] = 25'b10110001_11101000_10011001_1;
      patterns[45547] = 25'b10110001_11101001_10011010_1;
      patterns[45548] = 25'b10110001_11101010_10011011_1;
      patterns[45549] = 25'b10110001_11101011_10011100_1;
      patterns[45550] = 25'b10110001_11101100_10011101_1;
      patterns[45551] = 25'b10110001_11101101_10011110_1;
      patterns[45552] = 25'b10110001_11101110_10011111_1;
      patterns[45553] = 25'b10110001_11101111_10100000_1;
      patterns[45554] = 25'b10110001_11110000_10100001_1;
      patterns[45555] = 25'b10110001_11110001_10100010_1;
      patterns[45556] = 25'b10110001_11110010_10100011_1;
      patterns[45557] = 25'b10110001_11110011_10100100_1;
      patterns[45558] = 25'b10110001_11110100_10100101_1;
      patterns[45559] = 25'b10110001_11110101_10100110_1;
      patterns[45560] = 25'b10110001_11110110_10100111_1;
      patterns[45561] = 25'b10110001_11110111_10101000_1;
      patterns[45562] = 25'b10110001_11111000_10101001_1;
      patterns[45563] = 25'b10110001_11111001_10101010_1;
      patterns[45564] = 25'b10110001_11111010_10101011_1;
      patterns[45565] = 25'b10110001_11111011_10101100_1;
      patterns[45566] = 25'b10110001_11111100_10101101_1;
      patterns[45567] = 25'b10110001_11111101_10101110_1;
      patterns[45568] = 25'b10110001_11111110_10101111_1;
      patterns[45569] = 25'b10110001_11111111_10110000_1;
      patterns[45570] = 25'b10110010_00000000_10110010_0;
      patterns[45571] = 25'b10110010_00000001_10110011_0;
      patterns[45572] = 25'b10110010_00000010_10110100_0;
      patterns[45573] = 25'b10110010_00000011_10110101_0;
      patterns[45574] = 25'b10110010_00000100_10110110_0;
      patterns[45575] = 25'b10110010_00000101_10110111_0;
      patterns[45576] = 25'b10110010_00000110_10111000_0;
      patterns[45577] = 25'b10110010_00000111_10111001_0;
      patterns[45578] = 25'b10110010_00001000_10111010_0;
      patterns[45579] = 25'b10110010_00001001_10111011_0;
      patterns[45580] = 25'b10110010_00001010_10111100_0;
      patterns[45581] = 25'b10110010_00001011_10111101_0;
      patterns[45582] = 25'b10110010_00001100_10111110_0;
      patterns[45583] = 25'b10110010_00001101_10111111_0;
      patterns[45584] = 25'b10110010_00001110_11000000_0;
      patterns[45585] = 25'b10110010_00001111_11000001_0;
      patterns[45586] = 25'b10110010_00010000_11000010_0;
      patterns[45587] = 25'b10110010_00010001_11000011_0;
      patterns[45588] = 25'b10110010_00010010_11000100_0;
      patterns[45589] = 25'b10110010_00010011_11000101_0;
      patterns[45590] = 25'b10110010_00010100_11000110_0;
      patterns[45591] = 25'b10110010_00010101_11000111_0;
      patterns[45592] = 25'b10110010_00010110_11001000_0;
      patterns[45593] = 25'b10110010_00010111_11001001_0;
      patterns[45594] = 25'b10110010_00011000_11001010_0;
      patterns[45595] = 25'b10110010_00011001_11001011_0;
      patterns[45596] = 25'b10110010_00011010_11001100_0;
      patterns[45597] = 25'b10110010_00011011_11001101_0;
      patterns[45598] = 25'b10110010_00011100_11001110_0;
      patterns[45599] = 25'b10110010_00011101_11001111_0;
      patterns[45600] = 25'b10110010_00011110_11010000_0;
      patterns[45601] = 25'b10110010_00011111_11010001_0;
      patterns[45602] = 25'b10110010_00100000_11010010_0;
      patterns[45603] = 25'b10110010_00100001_11010011_0;
      patterns[45604] = 25'b10110010_00100010_11010100_0;
      patterns[45605] = 25'b10110010_00100011_11010101_0;
      patterns[45606] = 25'b10110010_00100100_11010110_0;
      patterns[45607] = 25'b10110010_00100101_11010111_0;
      patterns[45608] = 25'b10110010_00100110_11011000_0;
      patterns[45609] = 25'b10110010_00100111_11011001_0;
      patterns[45610] = 25'b10110010_00101000_11011010_0;
      patterns[45611] = 25'b10110010_00101001_11011011_0;
      patterns[45612] = 25'b10110010_00101010_11011100_0;
      patterns[45613] = 25'b10110010_00101011_11011101_0;
      patterns[45614] = 25'b10110010_00101100_11011110_0;
      patterns[45615] = 25'b10110010_00101101_11011111_0;
      patterns[45616] = 25'b10110010_00101110_11100000_0;
      patterns[45617] = 25'b10110010_00101111_11100001_0;
      patterns[45618] = 25'b10110010_00110000_11100010_0;
      patterns[45619] = 25'b10110010_00110001_11100011_0;
      patterns[45620] = 25'b10110010_00110010_11100100_0;
      patterns[45621] = 25'b10110010_00110011_11100101_0;
      patterns[45622] = 25'b10110010_00110100_11100110_0;
      patterns[45623] = 25'b10110010_00110101_11100111_0;
      patterns[45624] = 25'b10110010_00110110_11101000_0;
      patterns[45625] = 25'b10110010_00110111_11101001_0;
      patterns[45626] = 25'b10110010_00111000_11101010_0;
      patterns[45627] = 25'b10110010_00111001_11101011_0;
      patterns[45628] = 25'b10110010_00111010_11101100_0;
      patterns[45629] = 25'b10110010_00111011_11101101_0;
      patterns[45630] = 25'b10110010_00111100_11101110_0;
      patterns[45631] = 25'b10110010_00111101_11101111_0;
      patterns[45632] = 25'b10110010_00111110_11110000_0;
      patterns[45633] = 25'b10110010_00111111_11110001_0;
      patterns[45634] = 25'b10110010_01000000_11110010_0;
      patterns[45635] = 25'b10110010_01000001_11110011_0;
      patterns[45636] = 25'b10110010_01000010_11110100_0;
      patterns[45637] = 25'b10110010_01000011_11110101_0;
      patterns[45638] = 25'b10110010_01000100_11110110_0;
      patterns[45639] = 25'b10110010_01000101_11110111_0;
      patterns[45640] = 25'b10110010_01000110_11111000_0;
      patterns[45641] = 25'b10110010_01000111_11111001_0;
      patterns[45642] = 25'b10110010_01001000_11111010_0;
      patterns[45643] = 25'b10110010_01001001_11111011_0;
      patterns[45644] = 25'b10110010_01001010_11111100_0;
      patterns[45645] = 25'b10110010_01001011_11111101_0;
      patterns[45646] = 25'b10110010_01001100_11111110_0;
      patterns[45647] = 25'b10110010_01001101_11111111_0;
      patterns[45648] = 25'b10110010_01001110_00000000_1;
      patterns[45649] = 25'b10110010_01001111_00000001_1;
      patterns[45650] = 25'b10110010_01010000_00000010_1;
      patterns[45651] = 25'b10110010_01010001_00000011_1;
      patterns[45652] = 25'b10110010_01010010_00000100_1;
      patterns[45653] = 25'b10110010_01010011_00000101_1;
      patterns[45654] = 25'b10110010_01010100_00000110_1;
      patterns[45655] = 25'b10110010_01010101_00000111_1;
      patterns[45656] = 25'b10110010_01010110_00001000_1;
      patterns[45657] = 25'b10110010_01010111_00001001_1;
      patterns[45658] = 25'b10110010_01011000_00001010_1;
      patterns[45659] = 25'b10110010_01011001_00001011_1;
      patterns[45660] = 25'b10110010_01011010_00001100_1;
      patterns[45661] = 25'b10110010_01011011_00001101_1;
      patterns[45662] = 25'b10110010_01011100_00001110_1;
      patterns[45663] = 25'b10110010_01011101_00001111_1;
      patterns[45664] = 25'b10110010_01011110_00010000_1;
      patterns[45665] = 25'b10110010_01011111_00010001_1;
      patterns[45666] = 25'b10110010_01100000_00010010_1;
      patterns[45667] = 25'b10110010_01100001_00010011_1;
      patterns[45668] = 25'b10110010_01100010_00010100_1;
      patterns[45669] = 25'b10110010_01100011_00010101_1;
      patterns[45670] = 25'b10110010_01100100_00010110_1;
      patterns[45671] = 25'b10110010_01100101_00010111_1;
      patterns[45672] = 25'b10110010_01100110_00011000_1;
      patterns[45673] = 25'b10110010_01100111_00011001_1;
      patterns[45674] = 25'b10110010_01101000_00011010_1;
      patterns[45675] = 25'b10110010_01101001_00011011_1;
      patterns[45676] = 25'b10110010_01101010_00011100_1;
      patterns[45677] = 25'b10110010_01101011_00011101_1;
      patterns[45678] = 25'b10110010_01101100_00011110_1;
      patterns[45679] = 25'b10110010_01101101_00011111_1;
      patterns[45680] = 25'b10110010_01101110_00100000_1;
      patterns[45681] = 25'b10110010_01101111_00100001_1;
      patterns[45682] = 25'b10110010_01110000_00100010_1;
      patterns[45683] = 25'b10110010_01110001_00100011_1;
      patterns[45684] = 25'b10110010_01110010_00100100_1;
      patterns[45685] = 25'b10110010_01110011_00100101_1;
      patterns[45686] = 25'b10110010_01110100_00100110_1;
      patterns[45687] = 25'b10110010_01110101_00100111_1;
      patterns[45688] = 25'b10110010_01110110_00101000_1;
      patterns[45689] = 25'b10110010_01110111_00101001_1;
      patterns[45690] = 25'b10110010_01111000_00101010_1;
      patterns[45691] = 25'b10110010_01111001_00101011_1;
      patterns[45692] = 25'b10110010_01111010_00101100_1;
      patterns[45693] = 25'b10110010_01111011_00101101_1;
      patterns[45694] = 25'b10110010_01111100_00101110_1;
      patterns[45695] = 25'b10110010_01111101_00101111_1;
      patterns[45696] = 25'b10110010_01111110_00110000_1;
      patterns[45697] = 25'b10110010_01111111_00110001_1;
      patterns[45698] = 25'b10110010_10000000_00110010_1;
      patterns[45699] = 25'b10110010_10000001_00110011_1;
      patterns[45700] = 25'b10110010_10000010_00110100_1;
      patterns[45701] = 25'b10110010_10000011_00110101_1;
      patterns[45702] = 25'b10110010_10000100_00110110_1;
      patterns[45703] = 25'b10110010_10000101_00110111_1;
      patterns[45704] = 25'b10110010_10000110_00111000_1;
      patterns[45705] = 25'b10110010_10000111_00111001_1;
      patterns[45706] = 25'b10110010_10001000_00111010_1;
      patterns[45707] = 25'b10110010_10001001_00111011_1;
      patterns[45708] = 25'b10110010_10001010_00111100_1;
      patterns[45709] = 25'b10110010_10001011_00111101_1;
      patterns[45710] = 25'b10110010_10001100_00111110_1;
      patterns[45711] = 25'b10110010_10001101_00111111_1;
      patterns[45712] = 25'b10110010_10001110_01000000_1;
      patterns[45713] = 25'b10110010_10001111_01000001_1;
      patterns[45714] = 25'b10110010_10010000_01000010_1;
      patterns[45715] = 25'b10110010_10010001_01000011_1;
      patterns[45716] = 25'b10110010_10010010_01000100_1;
      patterns[45717] = 25'b10110010_10010011_01000101_1;
      patterns[45718] = 25'b10110010_10010100_01000110_1;
      patterns[45719] = 25'b10110010_10010101_01000111_1;
      patterns[45720] = 25'b10110010_10010110_01001000_1;
      patterns[45721] = 25'b10110010_10010111_01001001_1;
      patterns[45722] = 25'b10110010_10011000_01001010_1;
      patterns[45723] = 25'b10110010_10011001_01001011_1;
      patterns[45724] = 25'b10110010_10011010_01001100_1;
      patterns[45725] = 25'b10110010_10011011_01001101_1;
      patterns[45726] = 25'b10110010_10011100_01001110_1;
      patterns[45727] = 25'b10110010_10011101_01001111_1;
      patterns[45728] = 25'b10110010_10011110_01010000_1;
      patterns[45729] = 25'b10110010_10011111_01010001_1;
      patterns[45730] = 25'b10110010_10100000_01010010_1;
      patterns[45731] = 25'b10110010_10100001_01010011_1;
      patterns[45732] = 25'b10110010_10100010_01010100_1;
      patterns[45733] = 25'b10110010_10100011_01010101_1;
      patterns[45734] = 25'b10110010_10100100_01010110_1;
      patterns[45735] = 25'b10110010_10100101_01010111_1;
      patterns[45736] = 25'b10110010_10100110_01011000_1;
      patterns[45737] = 25'b10110010_10100111_01011001_1;
      patterns[45738] = 25'b10110010_10101000_01011010_1;
      patterns[45739] = 25'b10110010_10101001_01011011_1;
      patterns[45740] = 25'b10110010_10101010_01011100_1;
      patterns[45741] = 25'b10110010_10101011_01011101_1;
      patterns[45742] = 25'b10110010_10101100_01011110_1;
      patterns[45743] = 25'b10110010_10101101_01011111_1;
      patterns[45744] = 25'b10110010_10101110_01100000_1;
      patterns[45745] = 25'b10110010_10101111_01100001_1;
      patterns[45746] = 25'b10110010_10110000_01100010_1;
      patterns[45747] = 25'b10110010_10110001_01100011_1;
      patterns[45748] = 25'b10110010_10110010_01100100_1;
      patterns[45749] = 25'b10110010_10110011_01100101_1;
      patterns[45750] = 25'b10110010_10110100_01100110_1;
      patterns[45751] = 25'b10110010_10110101_01100111_1;
      patterns[45752] = 25'b10110010_10110110_01101000_1;
      patterns[45753] = 25'b10110010_10110111_01101001_1;
      patterns[45754] = 25'b10110010_10111000_01101010_1;
      patterns[45755] = 25'b10110010_10111001_01101011_1;
      patterns[45756] = 25'b10110010_10111010_01101100_1;
      patterns[45757] = 25'b10110010_10111011_01101101_1;
      patterns[45758] = 25'b10110010_10111100_01101110_1;
      patterns[45759] = 25'b10110010_10111101_01101111_1;
      patterns[45760] = 25'b10110010_10111110_01110000_1;
      patterns[45761] = 25'b10110010_10111111_01110001_1;
      patterns[45762] = 25'b10110010_11000000_01110010_1;
      patterns[45763] = 25'b10110010_11000001_01110011_1;
      patterns[45764] = 25'b10110010_11000010_01110100_1;
      patterns[45765] = 25'b10110010_11000011_01110101_1;
      patterns[45766] = 25'b10110010_11000100_01110110_1;
      patterns[45767] = 25'b10110010_11000101_01110111_1;
      patterns[45768] = 25'b10110010_11000110_01111000_1;
      patterns[45769] = 25'b10110010_11000111_01111001_1;
      patterns[45770] = 25'b10110010_11001000_01111010_1;
      patterns[45771] = 25'b10110010_11001001_01111011_1;
      patterns[45772] = 25'b10110010_11001010_01111100_1;
      patterns[45773] = 25'b10110010_11001011_01111101_1;
      patterns[45774] = 25'b10110010_11001100_01111110_1;
      patterns[45775] = 25'b10110010_11001101_01111111_1;
      patterns[45776] = 25'b10110010_11001110_10000000_1;
      patterns[45777] = 25'b10110010_11001111_10000001_1;
      patterns[45778] = 25'b10110010_11010000_10000010_1;
      patterns[45779] = 25'b10110010_11010001_10000011_1;
      patterns[45780] = 25'b10110010_11010010_10000100_1;
      patterns[45781] = 25'b10110010_11010011_10000101_1;
      patterns[45782] = 25'b10110010_11010100_10000110_1;
      patterns[45783] = 25'b10110010_11010101_10000111_1;
      patterns[45784] = 25'b10110010_11010110_10001000_1;
      patterns[45785] = 25'b10110010_11010111_10001001_1;
      patterns[45786] = 25'b10110010_11011000_10001010_1;
      patterns[45787] = 25'b10110010_11011001_10001011_1;
      patterns[45788] = 25'b10110010_11011010_10001100_1;
      patterns[45789] = 25'b10110010_11011011_10001101_1;
      patterns[45790] = 25'b10110010_11011100_10001110_1;
      patterns[45791] = 25'b10110010_11011101_10001111_1;
      patterns[45792] = 25'b10110010_11011110_10010000_1;
      patterns[45793] = 25'b10110010_11011111_10010001_1;
      patterns[45794] = 25'b10110010_11100000_10010010_1;
      patterns[45795] = 25'b10110010_11100001_10010011_1;
      patterns[45796] = 25'b10110010_11100010_10010100_1;
      patterns[45797] = 25'b10110010_11100011_10010101_1;
      patterns[45798] = 25'b10110010_11100100_10010110_1;
      patterns[45799] = 25'b10110010_11100101_10010111_1;
      patterns[45800] = 25'b10110010_11100110_10011000_1;
      patterns[45801] = 25'b10110010_11100111_10011001_1;
      patterns[45802] = 25'b10110010_11101000_10011010_1;
      patterns[45803] = 25'b10110010_11101001_10011011_1;
      patterns[45804] = 25'b10110010_11101010_10011100_1;
      patterns[45805] = 25'b10110010_11101011_10011101_1;
      patterns[45806] = 25'b10110010_11101100_10011110_1;
      patterns[45807] = 25'b10110010_11101101_10011111_1;
      patterns[45808] = 25'b10110010_11101110_10100000_1;
      patterns[45809] = 25'b10110010_11101111_10100001_1;
      patterns[45810] = 25'b10110010_11110000_10100010_1;
      patterns[45811] = 25'b10110010_11110001_10100011_1;
      patterns[45812] = 25'b10110010_11110010_10100100_1;
      patterns[45813] = 25'b10110010_11110011_10100101_1;
      patterns[45814] = 25'b10110010_11110100_10100110_1;
      patterns[45815] = 25'b10110010_11110101_10100111_1;
      patterns[45816] = 25'b10110010_11110110_10101000_1;
      patterns[45817] = 25'b10110010_11110111_10101001_1;
      patterns[45818] = 25'b10110010_11111000_10101010_1;
      patterns[45819] = 25'b10110010_11111001_10101011_1;
      patterns[45820] = 25'b10110010_11111010_10101100_1;
      patterns[45821] = 25'b10110010_11111011_10101101_1;
      patterns[45822] = 25'b10110010_11111100_10101110_1;
      patterns[45823] = 25'b10110010_11111101_10101111_1;
      patterns[45824] = 25'b10110010_11111110_10110000_1;
      patterns[45825] = 25'b10110010_11111111_10110001_1;
      patterns[45826] = 25'b10110011_00000000_10110011_0;
      patterns[45827] = 25'b10110011_00000001_10110100_0;
      patterns[45828] = 25'b10110011_00000010_10110101_0;
      patterns[45829] = 25'b10110011_00000011_10110110_0;
      patterns[45830] = 25'b10110011_00000100_10110111_0;
      patterns[45831] = 25'b10110011_00000101_10111000_0;
      patterns[45832] = 25'b10110011_00000110_10111001_0;
      patterns[45833] = 25'b10110011_00000111_10111010_0;
      patterns[45834] = 25'b10110011_00001000_10111011_0;
      patterns[45835] = 25'b10110011_00001001_10111100_0;
      patterns[45836] = 25'b10110011_00001010_10111101_0;
      patterns[45837] = 25'b10110011_00001011_10111110_0;
      patterns[45838] = 25'b10110011_00001100_10111111_0;
      patterns[45839] = 25'b10110011_00001101_11000000_0;
      patterns[45840] = 25'b10110011_00001110_11000001_0;
      patterns[45841] = 25'b10110011_00001111_11000010_0;
      patterns[45842] = 25'b10110011_00010000_11000011_0;
      patterns[45843] = 25'b10110011_00010001_11000100_0;
      patterns[45844] = 25'b10110011_00010010_11000101_0;
      patterns[45845] = 25'b10110011_00010011_11000110_0;
      patterns[45846] = 25'b10110011_00010100_11000111_0;
      patterns[45847] = 25'b10110011_00010101_11001000_0;
      patterns[45848] = 25'b10110011_00010110_11001001_0;
      patterns[45849] = 25'b10110011_00010111_11001010_0;
      patterns[45850] = 25'b10110011_00011000_11001011_0;
      patterns[45851] = 25'b10110011_00011001_11001100_0;
      patterns[45852] = 25'b10110011_00011010_11001101_0;
      patterns[45853] = 25'b10110011_00011011_11001110_0;
      patterns[45854] = 25'b10110011_00011100_11001111_0;
      patterns[45855] = 25'b10110011_00011101_11010000_0;
      patterns[45856] = 25'b10110011_00011110_11010001_0;
      patterns[45857] = 25'b10110011_00011111_11010010_0;
      patterns[45858] = 25'b10110011_00100000_11010011_0;
      patterns[45859] = 25'b10110011_00100001_11010100_0;
      patterns[45860] = 25'b10110011_00100010_11010101_0;
      patterns[45861] = 25'b10110011_00100011_11010110_0;
      patterns[45862] = 25'b10110011_00100100_11010111_0;
      patterns[45863] = 25'b10110011_00100101_11011000_0;
      patterns[45864] = 25'b10110011_00100110_11011001_0;
      patterns[45865] = 25'b10110011_00100111_11011010_0;
      patterns[45866] = 25'b10110011_00101000_11011011_0;
      patterns[45867] = 25'b10110011_00101001_11011100_0;
      patterns[45868] = 25'b10110011_00101010_11011101_0;
      patterns[45869] = 25'b10110011_00101011_11011110_0;
      patterns[45870] = 25'b10110011_00101100_11011111_0;
      patterns[45871] = 25'b10110011_00101101_11100000_0;
      patterns[45872] = 25'b10110011_00101110_11100001_0;
      patterns[45873] = 25'b10110011_00101111_11100010_0;
      patterns[45874] = 25'b10110011_00110000_11100011_0;
      patterns[45875] = 25'b10110011_00110001_11100100_0;
      patterns[45876] = 25'b10110011_00110010_11100101_0;
      patterns[45877] = 25'b10110011_00110011_11100110_0;
      patterns[45878] = 25'b10110011_00110100_11100111_0;
      patterns[45879] = 25'b10110011_00110101_11101000_0;
      patterns[45880] = 25'b10110011_00110110_11101001_0;
      patterns[45881] = 25'b10110011_00110111_11101010_0;
      patterns[45882] = 25'b10110011_00111000_11101011_0;
      patterns[45883] = 25'b10110011_00111001_11101100_0;
      patterns[45884] = 25'b10110011_00111010_11101101_0;
      patterns[45885] = 25'b10110011_00111011_11101110_0;
      patterns[45886] = 25'b10110011_00111100_11101111_0;
      patterns[45887] = 25'b10110011_00111101_11110000_0;
      patterns[45888] = 25'b10110011_00111110_11110001_0;
      patterns[45889] = 25'b10110011_00111111_11110010_0;
      patterns[45890] = 25'b10110011_01000000_11110011_0;
      patterns[45891] = 25'b10110011_01000001_11110100_0;
      patterns[45892] = 25'b10110011_01000010_11110101_0;
      patterns[45893] = 25'b10110011_01000011_11110110_0;
      patterns[45894] = 25'b10110011_01000100_11110111_0;
      patterns[45895] = 25'b10110011_01000101_11111000_0;
      patterns[45896] = 25'b10110011_01000110_11111001_0;
      patterns[45897] = 25'b10110011_01000111_11111010_0;
      patterns[45898] = 25'b10110011_01001000_11111011_0;
      patterns[45899] = 25'b10110011_01001001_11111100_0;
      patterns[45900] = 25'b10110011_01001010_11111101_0;
      patterns[45901] = 25'b10110011_01001011_11111110_0;
      patterns[45902] = 25'b10110011_01001100_11111111_0;
      patterns[45903] = 25'b10110011_01001101_00000000_1;
      patterns[45904] = 25'b10110011_01001110_00000001_1;
      patterns[45905] = 25'b10110011_01001111_00000010_1;
      patterns[45906] = 25'b10110011_01010000_00000011_1;
      patterns[45907] = 25'b10110011_01010001_00000100_1;
      patterns[45908] = 25'b10110011_01010010_00000101_1;
      patterns[45909] = 25'b10110011_01010011_00000110_1;
      patterns[45910] = 25'b10110011_01010100_00000111_1;
      patterns[45911] = 25'b10110011_01010101_00001000_1;
      patterns[45912] = 25'b10110011_01010110_00001001_1;
      patterns[45913] = 25'b10110011_01010111_00001010_1;
      patterns[45914] = 25'b10110011_01011000_00001011_1;
      patterns[45915] = 25'b10110011_01011001_00001100_1;
      patterns[45916] = 25'b10110011_01011010_00001101_1;
      patterns[45917] = 25'b10110011_01011011_00001110_1;
      patterns[45918] = 25'b10110011_01011100_00001111_1;
      patterns[45919] = 25'b10110011_01011101_00010000_1;
      patterns[45920] = 25'b10110011_01011110_00010001_1;
      patterns[45921] = 25'b10110011_01011111_00010010_1;
      patterns[45922] = 25'b10110011_01100000_00010011_1;
      patterns[45923] = 25'b10110011_01100001_00010100_1;
      patterns[45924] = 25'b10110011_01100010_00010101_1;
      patterns[45925] = 25'b10110011_01100011_00010110_1;
      patterns[45926] = 25'b10110011_01100100_00010111_1;
      patterns[45927] = 25'b10110011_01100101_00011000_1;
      patterns[45928] = 25'b10110011_01100110_00011001_1;
      patterns[45929] = 25'b10110011_01100111_00011010_1;
      patterns[45930] = 25'b10110011_01101000_00011011_1;
      patterns[45931] = 25'b10110011_01101001_00011100_1;
      patterns[45932] = 25'b10110011_01101010_00011101_1;
      patterns[45933] = 25'b10110011_01101011_00011110_1;
      patterns[45934] = 25'b10110011_01101100_00011111_1;
      patterns[45935] = 25'b10110011_01101101_00100000_1;
      patterns[45936] = 25'b10110011_01101110_00100001_1;
      patterns[45937] = 25'b10110011_01101111_00100010_1;
      patterns[45938] = 25'b10110011_01110000_00100011_1;
      patterns[45939] = 25'b10110011_01110001_00100100_1;
      patterns[45940] = 25'b10110011_01110010_00100101_1;
      patterns[45941] = 25'b10110011_01110011_00100110_1;
      patterns[45942] = 25'b10110011_01110100_00100111_1;
      patterns[45943] = 25'b10110011_01110101_00101000_1;
      patterns[45944] = 25'b10110011_01110110_00101001_1;
      patterns[45945] = 25'b10110011_01110111_00101010_1;
      patterns[45946] = 25'b10110011_01111000_00101011_1;
      patterns[45947] = 25'b10110011_01111001_00101100_1;
      patterns[45948] = 25'b10110011_01111010_00101101_1;
      patterns[45949] = 25'b10110011_01111011_00101110_1;
      patterns[45950] = 25'b10110011_01111100_00101111_1;
      patterns[45951] = 25'b10110011_01111101_00110000_1;
      patterns[45952] = 25'b10110011_01111110_00110001_1;
      patterns[45953] = 25'b10110011_01111111_00110010_1;
      patterns[45954] = 25'b10110011_10000000_00110011_1;
      patterns[45955] = 25'b10110011_10000001_00110100_1;
      patterns[45956] = 25'b10110011_10000010_00110101_1;
      patterns[45957] = 25'b10110011_10000011_00110110_1;
      patterns[45958] = 25'b10110011_10000100_00110111_1;
      patterns[45959] = 25'b10110011_10000101_00111000_1;
      patterns[45960] = 25'b10110011_10000110_00111001_1;
      patterns[45961] = 25'b10110011_10000111_00111010_1;
      patterns[45962] = 25'b10110011_10001000_00111011_1;
      patterns[45963] = 25'b10110011_10001001_00111100_1;
      patterns[45964] = 25'b10110011_10001010_00111101_1;
      patterns[45965] = 25'b10110011_10001011_00111110_1;
      patterns[45966] = 25'b10110011_10001100_00111111_1;
      patterns[45967] = 25'b10110011_10001101_01000000_1;
      patterns[45968] = 25'b10110011_10001110_01000001_1;
      patterns[45969] = 25'b10110011_10001111_01000010_1;
      patterns[45970] = 25'b10110011_10010000_01000011_1;
      patterns[45971] = 25'b10110011_10010001_01000100_1;
      patterns[45972] = 25'b10110011_10010010_01000101_1;
      patterns[45973] = 25'b10110011_10010011_01000110_1;
      patterns[45974] = 25'b10110011_10010100_01000111_1;
      patterns[45975] = 25'b10110011_10010101_01001000_1;
      patterns[45976] = 25'b10110011_10010110_01001001_1;
      patterns[45977] = 25'b10110011_10010111_01001010_1;
      patterns[45978] = 25'b10110011_10011000_01001011_1;
      patterns[45979] = 25'b10110011_10011001_01001100_1;
      patterns[45980] = 25'b10110011_10011010_01001101_1;
      patterns[45981] = 25'b10110011_10011011_01001110_1;
      patterns[45982] = 25'b10110011_10011100_01001111_1;
      patterns[45983] = 25'b10110011_10011101_01010000_1;
      patterns[45984] = 25'b10110011_10011110_01010001_1;
      patterns[45985] = 25'b10110011_10011111_01010010_1;
      patterns[45986] = 25'b10110011_10100000_01010011_1;
      patterns[45987] = 25'b10110011_10100001_01010100_1;
      patterns[45988] = 25'b10110011_10100010_01010101_1;
      patterns[45989] = 25'b10110011_10100011_01010110_1;
      patterns[45990] = 25'b10110011_10100100_01010111_1;
      patterns[45991] = 25'b10110011_10100101_01011000_1;
      patterns[45992] = 25'b10110011_10100110_01011001_1;
      patterns[45993] = 25'b10110011_10100111_01011010_1;
      patterns[45994] = 25'b10110011_10101000_01011011_1;
      patterns[45995] = 25'b10110011_10101001_01011100_1;
      patterns[45996] = 25'b10110011_10101010_01011101_1;
      patterns[45997] = 25'b10110011_10101011_01011110_1;
      patterns[45998] = 25'b10110011_10101100_01011111_1;
      patterns[45999] = 25'b10110011_10101101_01100000_1;
      patterns[46000] = 25'b10110011_10101110_01100001_1;
      patterns[46001] = 25'b10110011_10101111_01100010_1;
      patterns[46002] = 25'b10110011_10110000_01100011_1;
      patterns[46003] = 25'b10110011_10110001_01100100_1;
      patterns[46004] = 25'b10110011_10110010_01100101_1;
      patterns[46005] = 25'b10110011_10110011_01100110_1;
      patterns[46006] = 25'b10110011_10110100_01100111_1;
      patterns[46007] = 25'b10110011_10110101_01101000_1;
      patterns[46008] = 25'b10110011_10110110_01101001_1;
      patterns[46009] = 25'b10110011_10110111_01101010_1;
      patterns[46010] = 25'b10110011_10111000_01101011_1;
      patterns[46011] = 25'b10110011_10111001_01101100_1;
      patterns[46012] = 25'b10110011_10111010_01101101_1;
      patterns[46013] = 25'b10110011_10111011_01101110_1;
      patterns[46014] = 25'b10110011_10111100_01101111_1;
      patterns[46015] = 25'b10110011_10111101_01110000_1;
      patterns[46016] = 25'b10110011_10111110_01110001_1;
      patterns[46017] = 25'b10110011_10111111_01110010_1;
      patterns[46018] = 25'b10110011_11000000_01110011_1;
      patterns[46019] = 25'b10110011_11000001_01110100_1;
      patterns[46020] = 25'b10110011_11000010_01110101_1;
      patterns[46021] = 25'b10110011_11000011_01110110_1;
      patterns[46022] = 25'b10110011_11000100_01110111_1;
      patterns[46023] = 25'b10110011_11000101_01111000_1;
      patterns[46024] = 25'b10110011_11000110_01111001_1;
      patterns[46025] = 25'b10110011_11000111_01111010_1;
      patterns[46026] = 25'b10110011_11001000_01111011_1;
      patterns[46027] = 25'b10110011_11001001_01111100_1;
      patterns[46028] = 25'b10110011_11001010_01111101_1;
      patterns[46029] = 25'b10110011_11001011_01111110_1;
      patterns[46030] = 25'b10110011_11001100_01111111_1;
      patterns[46031] = 25'b10110011_11001101_10000000_1;
      patterns[46032] = 25'b10110011_11001110_10000001_1;
      patterns[46033] = 25'b10110011_11001111_10000010_1;
      patterns[46034] = 25'b10110011_11010000_10000011_1;
      patterns[46035] = 25'b10110011_11010001_10000100_1;
      patterns[46036] = 25'b10110011_11010010_10000101_1;
      patterns[46037] = 25'b10110011_11010011_10000110_1;
      patterns[46038] = 25'b10110011_11010100_10000111_1;
      patterns[46039] = 25'b10110011_11010101_10001000_1;
      patterns[46040] = 25'b10110011_11010110_10001001_1;
      patterns[46041] = 25'b10110011_11010111_10001010_1;
      patterns[46042] = 25'b10110011_11011000_10001011_1;
      patterns[46043] = 25'b10110011_11011001_10001100_1;
      patterns[46044] = 25'b10110011_11011010_10001101_1;
      patterns[46045] = 25'b10110011_11011011_10001110_1;
      patterns[46046] = 25'b10110011_11011100_10001111_1;
      patterns[46047] = 25'b10110011_11011101_10010000_1;
      patterns[46048] = 25'b10110011_11011110_10010001_1;
      patterns[46049] = 25'b10110011_11011111_10010010_1;
      patterns[46050] = 25'b10110011_11100000_10010011_1;
      patterns[46051] = 25'b10110011_11100001_10010100_1;
      patterns[46052] = 25'b10110011_11100010_10010101_1;
      patterns[46053] = 25'b10110011_11100011_10010110_1;
      patterns[46054] = 25'b10110011_11100100_10010111_1;
      patterns[46055] = 25'b10110011_11100101_10011000_1;
      patterns[46056] = 25'b10110011_11100110_10011001_1;
      patterns[46057] = 25'b10110011_11100111_10011010_1;
      patterns[46058] = 25'b10110011_11101000_10011011_1;
      patterns[46059] = 25'b10110011_11101001_10011100_1;
      patterns[46060] = 25'b10110011_11101010_10011101_1;
      patterns[46061] = 25'b10110011_11101011_10011110_1;
      patterns[46062] = 25'b10110011_11101100_10011111_1;
      patterns[46063] = 25'b10110011_11101101_10100000_1;
      patterns[46064] = 25'b10110011_11101110_10100001_1;
      patterns[46065] = 25'b10110011_11101111_10100010_1;
      patterns[46066] = 25'b10110011_11110000_10100011_1;
      patterns[46067] = 25'b10110011_11110001_10100100_1;
      patterns[46068] = 25'b10110011_11110010_10100101_1;
      patterns[46069] = 25'b10110011_11110011_10100110_1;
      patterns[46070] = 25'b10110011_11110100_10100111_1;
      patterns[46071] = 25'b10110011_11110101_10101000_1;
      patterns[46072] = 25'b10110011_11110110_10101001_1;
      patterns[46073] = 25'b10110011_11110111_10101010_1;
      patterns[46074] = 25'b10110011_11111000_10101011_1;
      patterns[46075] = 25'b10110011_11111001_10101100_1;
      patterns[46076] = 25'b10110011_11111010_10101101_1;
      patterns[46077] = 25'b10110011_11111011_10101110_1;
      patterns[46078] = 25'b10110011_11111100_10101111_1;
      patterns[46079] = 25'b10110011_11111101_10110000_1;
      patterns[46080] = 25'b10110011_11111110_10110001_1;
      patterns[46081] = 25'b10110011_11111111_10110010_1;
      patterns[46082] = 25'b10110100_00000000_10110100_0;
      patterns[46083] = 25'b10110100_00000001_10110101_0;
      patterns[46084] = 25'b10110100_00000010_10110110_0;
      patterns[46085] = 25'b10110100_00000011_10110111_0;
      patterns[46086] = 25'b10110100_00000100_10111000_0;
      patterns[46087] = 25'b10110100_00000101_10111001_0;
      patterns[46088] = 25'b10110100_00000110_10111010_0;
      patterns[46089] = 25'b10110100_00000111_10111011_0;
      patterns[46090] = 25'b10110100_00001000_10111100_0;
      patterns[46091] = 25'b10110100_00001001_10111101_0;
      patterns[46092] = 25'b10110100_00001010_10111110_0;
      patterns[46093] = 25'b10110100_00001011_10111111_0;
      patterns[46094] = 25'b10110100_00001100_11000000_0;
      patterns[46095] = 25'b10110100_00001101_11000001_0;
      patterns[46096] = 25'b10110100_00001110_11000010_0;
      patterns[46097] = 25'b10110100_00001111_11000011_0;
      patterns[46098] = 25'b10110100_00010000_11000100_0;
      patterns[46099] = 25'b10110100_00010001_11000101_0;
      patterns[46100] = 25'b10110100_00010010_11000110_0;
      patterns[46101] = 25'b10110100_00010011_11000111_0;
      patterns[46102] = 25'b10110100_00010100_11001000_0;
      patterns[46103] = 25'b10110100_00010101_11001001_0;
      patterns[46104] = 25'b10110100_00010110_11001010_0;
      patterns[46105] = 25'b10110100_00010111_11001011_0;
      patterns[46106] = 25'b10110100_00011000_11001100_0;
      patterns[46107] = 25'b10110100_00011001_11001101_0;
      patterns[46108] = 25'b10110100_00011010_11001110_0;
      patterns[46109] = 25'b10110100_00011011_11001111_0;
      patterns[46110] = 25'b10110100_00011100_11010000_0;
      patterns[46111] = 25'b10110100_00011101_11010001_0;
      patterns[46112] = 25'b10110100_00011110_11010010_0;
      patterns[46113] = 25'b10110100_00011111_11010011_0;
      patterns[46114] = 25'b10110100_00100000_11010100_0;
      patterns[46115] = 25'b10110100_00100001_11010101_0;
      patterns[46116] = 25'b10110100_00100010_11010110_0;
      patterns[46117] = 25'b10110100_00100011_11010111_0;
      patterns[46118] = 25'b10110100_00100100_11011000_0;
      patterns[46119] = 25'b10110100_00100101_11011001_0;
      patterns[46120] = 25'b10110100_00100110_11011010_0;
      patterns[46121] = 25'b10110100_00100111_11011011_0;
      patterns[46122] = 25'b10110100_00101000_11011100_0;
      patterns[46123] = 25'b10110100_00101001_11011101_0;
      patterns[46124] = 25'b10110100_00101010_11011110_0;
      patterns[46125] = 25'b10110100_00101011_11011111_0;
      patterns[46126] = 25'b10110100_00101100_11100000_0;
      patterns[46127] = 25'b10110100_00101101_11100001_0;
      patterns[46128] = 25'b10110100_00101110_11100010_0;
      patterns[46129] = 25'b10110100_00101111_11100011_0;
      patterns[46130] = 25'b10110100_00110000_11100100_0;
      patterns[46131] = 25'b10110100_00110001_11100101_0;
      patterns[46132] = 25'b10110100_00110010_11100110_0;
      patterns[46133] = 25'b10110100_00110011_11100111_0;
      patterns[46134] = 25'b10110100_00110100_11101000_0;
      patterns[46135] = 25'b10110100_00110101_11101001_0;
      patterns[46136] = 25'b10110100_00110110_11101010_0;
      patterns[46137] = 25'b10110100_00110111_11101011_0;
      patterns[46138] = 25'b10110100_00111000_11101100_0;
      patterns[46139] = 25'b10110100_00111001_11101101_0;
      patterns[46140] = 25'b10110100_00111010_11101110_0;
      patterns[46141] = 25'b10110100_00111011_11101111_0;
      patterns[46142] = 25'b10110100_00111100_11110000_0;
      patterns[46143] = 25'b10110100_00111101_11110001_0;
      patterns[46144] = 25'b10110100_00111110_11110010_0;
      patterns[46145] = 25'b10110100_00111111_11110011_0;
      patterns[46146] = 25'b10110100_01000000_11110100_0;
      patterns[46147] = 25'b10110100_01000001_11110101_0;
      patterns[46148] = 25'b10110100_01000010_11110110_0;
      patterns[46149] = 25'b10110100_01000011_11110111_0;
      patterns[46150] = 25'b10110100_01000100_11111000_0;
      patterns[46151] = 25'b10110100_01000101_11111001_0;
      patterns[46152] = 25'b10110100_01000110_11111010_0;
      patterns[46153] = 25'b10110100_01000111_11111011_0;
      patterns[46154] = 25'b10110100_01001000_11111100_0;
      patterns[46155] = 25'b10110100_01001001_11111101_0;
      patterns[46156] = 25'b10110100_01001010_11111110_0;
      patterns[46157] = 25'b10110100_01001011_11111111_0;
      patterns[46158] = 25'b10110100_01001100_00000000_1;
      patterns[46159] = 25'b10110100_01001101_00000001_1;
      patterns[46160] = 25'b10110100_01001110_00000010_1;
      patterns[46161] = 25'b10110100_01001111_00000011_1;
      patterns[46162] = 25'b10110100_01010000_00000100_1;
      patterns[46163] = 25'b10110100_01010001_00000101_1;
      patterns[46164] = 25'b10110100_01010010_00000110_1;
      patterns[46165] = 25'b10110100_01010011_00000111_1;
      patterns[46166] = 25'b10110100_01010100_00001000_1;
      patterns[46167] = 25'b10110100_01010101_00001001_1;
      patterns[46168] = 25'b10110100_01010110_00001010_1;
      patterns[46169] = 25'b10110100_01010111_00001011_1;
      patterns[46170] = 25'b10110100_01011000_00001100_1;
      patterns[46171] = 25'b10110100_01011001_00001101_1;
      patterns[46172] = 25'b10110100_01011010_00001110_1;
      patterns[46173] = 25'b10110100_01011011_00001111_1;
      patterns[46174] = 25'b10110100_01011100_00010000_1;
      patterns[46175] = 25'b10110100_01011101_00010001_1;
      patterns[46176] = 25'b10110100_01011110_00010010_1;
      patterns[46177] = 25'b10110100_01011111_00010011_1;
      patterns[46178] = 25'b10110100_01100000_00010100_1;
      patterns[46179] = 25'b10110100_01100001_00010101_1;
      patterns[46180] = 25'b10110100_01100010_00010110_1;
      patterns[46181] = 25'b10110100_01100011_00010111_1;
      patterns[46182] = 25'b10110100_01100100_00011000_1;
      patterns[46183] = 25'b10110100_01100101_00011001_1;
      patterns[46184] = 25'b10110100_01100110_00011010_1;
      patterns[46185] = 25'b10110100_01100111_00011011_1;
      patterns[46186] = 25'b10110100_01101000_00011100_1;
      patterns[46187] = 25'b10110100_01101001_00011101_1;
      patterns[46188] = 25'b10110100_01101010_00011110_1;
      patterns[46189] = 25'b10110100_01101011_00011111_1;
      patterns[46190] = 25'b10110100_01101100_00100000_1;
      patterns[46191] = 25'b10110100_01101101_00100001_1;
      patterns[46192] = 25'b10110100_01101110_00100010_1;
      patterns[46193] = 25'b10110100_01101111_00100011_1;
      patterns[46194] = 25'b10110100_01110000_00100100_1;
      patterns[46195] = 25'b10110100_01110001_00100101_1;
      patterns[46196] = 25'b10110100_01110010_00100110_1;
      patterns[46197] = 25'b10110100_01110011_00100111_1;
      patterns[46198] = 25'b10110100_01110100_00101000_1;
      patterns[46199] = 25'b10110100_01110101_00101001_1;
      patterns[46200] = 25'b10110100_01110110_00101010_1;
      patterns[46201] = 25'b10110100_01110111_00101011_1;
      patterns[46202] = 25'b10110100_01111000_00101100_1;
      patterns[46203] = 25'b10110100_01111001_00101101_1;
      patterns[46204] = 25'b10110100_01111010_00101110_1;
      patterns[46205] = 25'b10110100_01111011_00101111_1;
      patterns[46206] = 25'b10110100_01111100_00110000_1;
      patterns[46207] = 25'b10110100_01111101_00110001_1;
      patterns[46208] = 25'b10110100_01111110_00110010_1;
      patterns[46209] = 25'b10110100_01111111_00110011_1;
      patterns[46210] = 25'b10110100_10000000_00110100_1;
      patterns[46211] = 25'b10110100_10000001_00110101_1;
      patterns[46212] = 25'b10110100_10000010_00110110_1;
      patterns[46213] = 25'b10110100_10000011_00110111_1;
      patterns[46214] = 25'b10110100_10000100_00111000_1;
      patterns[46215] = 25'b10110100_10000101_00111001_1;
      patterns[46216] = 25'b10110100_10000110_00111010_1;
      patterns[46217] = 25'b10110100_10000111_00111011_1;
      patterns[46218] = 25'b10110100_10001000_00111100_1;
      patterns[46219] = 25'b10110100_10001001_00111101_1;
      patterns[46220] = 25'b10110100_10001010_00111110_1;
      patterns[46221] = 25'b10110100_10001011_00111111_1;
      patterns[46222] = 25'b10110100_10001100_01000000_1;
      patterns[46223] = 25'b10110100_10001101_01000001_1;
      patterns[46224] = 25'b10110100_10001110_01000010_1;
      patterns[46225] = 25'b10110100_10001111_01000011_1;
      patterns[46226] = 25'b10110100_10010000_01000100_1;
      patterns[46227] = 25'b10110100_10010001_01000101_1;
      patterns[46228] = 25'b10110100_10010010_01000110_1;
      patterns[46229] = 25'b10110100_10010011_01000111_1;
      patterns[46230] = 25'b10110100_10010100_01001000_1;
      patterns[46231] = 25'b10110100_10010101_01001001_1;
      patterns[46232] = 25'b10110100_10010110_01001010_1;
      patterns[46233] = 25'b10110100_10010111_01001011_1;
      patterns[46234] = 25'b10110100_10011000_01001100_1;
      patterns[46235] = 25'b10110100_10011001_01001101_1;
      patterns[46236] = 25'b10110100_10011010_01001110_1;
      patterns[46237] = 25'b10110100_10011011_01001111_1;
      patterns[46238] = 25'b10110100_10011100_01010000_1;
      patterns[46239] = 25'b10110100_10011101_01010001_1;
      patterns[46240] = 25'b10110100_10011110_01010010_1;
      patterns[46241] = 25'b10110100_10011111_01010011_1;
      patterns[46242] = 25'b10110100_10100000_01010100_1;
      patterns[46243] = 25'b10110100_10100001_01010101_1;
      patterns[46244] = 25'b10110100_10100010_01010110_1;
      patterns[46245] = 25'b10110100_10100011_01010111_1;
      patterns[46246] = 25'b10110100_10100100_01011000_1;
      patterns[46247] = 25'b10110100_10100101_01011001_1;
      patterns[46248] = 25'b10110100_10100110_01011010_1;
      patterns[46249] = 25'b10110100_10100111_01011011_1;
      patterns[46250] = 25'b10110100_10101000_01011100_1;
      patterns[46251] = 25'b10110100_10101001_01011101_1;
      patterns[46252] = 25'b10110100_10101010_01011110_1;
      patterns[46253] = 25'b10110100_10101011_01011111_1;
      patterns[46254] = 25'b10110100_10101100_01100000_1;
      patterns[46255] = 25'b10110100_10101101_01100001_1;
      patterns[46256] = 25'b10110100_10101110_01100010_1;
      patterns[46257] = 25'b10110100_10101111_01100011_1;
      patterns[46258] = 25'b10110100_10110000_01100100_1;
      patterns[46259] = 25'b10110100_10110001_01100101_1;
      patterns[46260] = 25'b10110100_10110010_01100110_1;
      patterns[46261] = 25'b10110100_10110011_01100111_1;
      patterns[46262] = 25'b10110100_10110100_01101000_1;
      patterns[46263] = 25'b10110100_10110101_01101001_1;
      patterns[46264] = 25'b10110100_10110110_01101010_1;
      patterns[46265] = 25'b10110100_10110111_01101011_1;
      patterns[46266] = 25'b10110100_10111000_01101100_1;
      patterns[46267] = 25'b10110100_10111001_01101101_1;
      patterns[46268] = 25'b10110100_10111010_01101110_1;
      patterns[46269] = 25'b10110100_10111011_01101111_1;
      patterns[46270] = 25'b10110100_10111100_01110000_1;
      patterns[46271] = 25'b10110100_10111101_01110001_1;
      patterns[46272] = 25'b10110100_10111110_01110010_1;
      patterns[46273] = 25'b10110100_10111111_01110011_1;
      patterns[46274] = 25'b10110100_11000000_01110100_1;
      patterns[46275] = 25'b10110100_11000001_01110101_1;
      patterns[46276] = 25'b10110100_11000010_01110110_1;
      patterns[46277] = 25'b10110100_11000011_01110111_1;
      patterns[46278] = 25'b10110100_11000100_01111000_1;
      patterns[46279] = 25'b10110100_11000101_01111001_1;
      patterns[46280] = 25'b10110100_11000110_01111010_1;
      patterns[46281] = 25'b10110100_11000111_01111011_1;
      patterns[46282] = 25'b10110100_11001000_01111100_1;
      patterns[46283] = 25'b10110100_11001001_01111101_1;
      patterns[46284] = 25'b10110100_11001010_01111110_1;
      patterns[46285] = 25'b10110100_11001011_01111111_1;
      patterns[46286] = 25'b10110100_11001100_10000000_1;
      patterns[46287] = 25'b10110100_11001101_10000001_1;
      patterns[46288] = 25'b10110100_11001110_10000010_1;
      patterns[46289] = 25'b10110100_11001111_10000011_1;
      patterns[46290] = 25'b10110100_11010000_10000100_1;
      patterns[46291] = 25'b10110100_11010001_10000101_1;
      patterns[46292] = 25'b10110100_11010010_10000110_1;
      patterns[46293] = 25'b10110100_11010011_10000111_1;
      patterns[46294] = 25'b10110100_11010100_10001000_1;
      patterns[46295] = 25'b10110100_11010101_10001001_1;
      patterns[46296] = 25'b10110100_11010110_10001010_1;
      patterns[46297] = 25'b10110100_11010111_10001011_1;
      patterns[46298] = 25'b10110100_11011000_10001100_1;
      patterns[46299] = 25'b10110100_11011001_10001101_1;
      patterns[46300] = 25'b10110100_11011010_10001110_1;
      patterns[46301] = 25'b10110100_11011011_10001111_1;
      patterns[46302] = 25'b10110100_11011100_10010000_1;
      patterns[46303] = 25'b10110100_11011101_10010001_1;
      patterns[46304] = 25'b10110100_11011110_10010010_1;
      patterns[46305] = 25'b10110100_11011111_10010011_1;
      patterns[46306] = 25'b10110100_11100000_10010100_1;
      patterns[46307] = 25'b10110100_11100001_10010101_1;
      patterns[46308] = 25'b10110100_11100010_10010110_1;
      patterns[46309] = 25'b10110100_11100011_10010111_1;
      patterns[46310] = 25'b10110100_11100100_10011000_1;
      patterns[46311] = 25'b10110100_11100101_10011001_1;
      patterns[46312] = 25'b10110100_11100110_10011010_1;
      patterns[46313] = 25'b10110100_11100111_10011011_1;
      patterns[46314] = 25'b10110100_11101000_10011100_1;
      patterns[46315] = 25'b10110100_11101001_10011101_1;
      patterns[46316] = 25'b10110100_11101010_10011110_1;
      patterns[46317] = 25'b10110100_11101011_10011111_1;
      patterns[46318] = 25'b10110100_11101100_10100000_1;
      patterns[46319] = 25'b10110100_11101101_10100001_1;
      patterns[46320] = 25'b10110100_11101110_10100010_1;
      patterns[46321] = 25'b10110100_11101111_10100011_1;
      patterns[46322] = 25'b10110100_11110000_10100100_1;
      patterns[46323] = 25'b10110100_11110001_10100101_1;
      patterns[46324] = 25'b10110100_11110010_10100110_1;
      patterns[46325] = 25'b10110100_11110011_10100111_1;
      patterns[46326] = 25'b10110100_11110100_10101000_1;
      patterns[46327] = 25'b10110100_11110101_10101001_1;
      patterns[46328] = 25'b10110100_11110110_10101010_1;
      patterns[46329] = 25'b10110100_11110111_10101011_1;
      patterns[46330] = 25'b10110100_11111000_10101100_1;
      patterns[46331] = 25'b10110100_11111001_10101101_1;
      patterns[46332] = 25'b10110100_11111010_10101110_1;
      patterns[46333] = 25'b10110100_11111011_10101111_1;
      patterns[46334] = 25'b10110100_11111100_10110000_1;
      patterns[46335] = 25'b10110100_11111101_10110001_1;
      patterns[46336] = 25'b10110100_11111110_10110010_1;
      patterns[46337] = 25'b10110100_11111111_10110011_1;
      patterns[46338] = 25'b10110101_00000000_10110101_0;
      patterns[46339] = 25'b10110101_00000001_10110110_0;
      patterns[46340] = 25'b10110101_00000010_10110111_0;
      patterns[46341] = 25'b10110101_00000011_10111000_0;
      patterns[46342] = 25'b10110101_00000100_10111001_0;
      patterns[46343] = 25'b10110101_00000101_10111010_0;
      patterns[46344] = 25'b10110101_00000110_10111011_0;
      patterns[46345] = 25'b10110101_00000111_10111100_0;
      patterns[46346] = 25'b10110101_00001000_10111101_0;
      patterns[46347] = 25'b10110101_00001001_10111110_0;
      patterns[46348] = 25'b10110101_00001010_10111111_0;
      patterns[46349] = 25'b10110101_00001011_11000000_0;
      patterns[46350] = 25'b10110101_00001100_11000001_0;
      patterns[46351] = 25'b10110101_00001101_11000010_0;
      patterns[46352] = 25'b10110101_00001110_11000011_0;
      patterns[46353] = 25'b10110101_00001111_11000100_0;
      patterns[46354] = 25'b10110101_00010000_11000101_0;
      patterns[46355] = 25'b10110101_00010001_11000110_0;
      patterns[46356] = 25'b10110101_00010010_11000111_0;
      patterns[46357] = 25'b10110101_00010011_11001000_0;
      patterns[46358] = 25'b10110101_00010100_11001001_0;
      patterns[46359] = 25'b10110101_00010101_11001010_0;
      patterns[46360] = 25'b10110101_00010110_11001011_0;
      patterns[46361] = 25'b10110101_00010111_11001100_0;
      patterns[46362] = 25'b10110101_00011000_11001101_0;
      patterns[46363] = 25'b10110101_00011001_11001110_0;
      patterns[46364] = 25'b10110101_00011010_11001111_0;
      patterns[46365] = 25'b10110101_00011011_11010000_0;
      patterns[46366] = 25'b10110101_00011100_11010001_0;
      patterns[46367] = 25'b10110101_00011101_11010010_0;
      patterns[46368] = 25'b10110101_00011110_11010011_0;
      patterns[46369] = 25'b10110101_00011111_11010100_0;
      patterns[46370] = 25'b10110101_00100000_11010101_0;
      patterns[46371] = 25'b10110101_00100001_11010110_0;
      patterns[46372] = 25'b10110101_00100010_11010111_0;
      patterns[46373] = 25'b10110101_00100011_11011000_0;
      patterns[46374] = 25'b10110101_00100100_11011001_0;
      patterns[46375] = 25'b10110101_00100101_11011010_0;
      patterns[46376] = 25'b10110101_00100110_11011011_0;
      patterns[46377] = 25'b10110101_00100111_11011100_0;
      patterns[46378] = 25'b10110101_00101000_11011101_0;
      patterns[46379] = 25'b10110101_00101001_11011110_0;
      patterns[46380] = 25'b10110101_00101010_11011111_0;
      patterns[46381] = 25'b10110101_00101011_11100000_0;
      patterns[46382] = 25'b10110101_00101100_11100001_0;
      patterns[46383] = 25'b10110101_00101101_11100010_0;
      patterns[46384] = 25'b10110101_00101110_11100011_0;
      patterns[46385] = 25'b10110101_00101111_11100100_0;
      patterns[46386] = 25'b10110101_00110000_11100101_0;
      patterns[46387] = 25'b10110101_00110001_11100110_0;
      patterns[46388] = 25'b10110101_00110010_11100111_0;
      patterns[46389] = 25'b10110101_00110011_11101000_0;
      patterns[46390] = 25'b10110101_00110100_11101001_0;
      patterns[46391] = 25'b10110101_00110101_11101010_0;
      patterns[46392] = 25'b10110101_00110110_11101011_0;
      patterns[46393] = 25'b10110101_00110111_11101100_0;
      patterns[46394] = 25'b10110101_00111000_11101101_0;
      patterns[46395] = 25'b10110101_00111001_11101110_0;
      patterns[46396] = 25'b10110101_00111010_11101111_0;
      patterns[46397] = 25'b10110101_00111011_11110000_0;
      patterns[46398] = 25'b10110101_00111100_11110001_0;
      patterns[46399] = 25'b10110101_00111101_11110010_0;
      patterns[46400] = 25'b10110101_00111110_11110011_0;
      patterns[46401] = 25'b10110101_00111111_11110100_0;
      patterns[46402] = 25'b10110101_01000000_11110101_0;
      patterns[46403] = 25'b10110101_01000001_11110110_0;
      patterns[46404] = 25'b10110101_01000010_11110111_0;
      patterns[46405] = 25'b10110101_01000011_11111000_0;
      patterns[46406] = 25'b10110101_01000100_11111001_0;
      patterns[46407] = 25'b10110101_01000101_11111010_0;
      patterns[46408] = 25'b10110101_01000110_11111011_0;
      patterns[46409] = 25'b10110101_01000111_11111100_0;
      patterns[46410] = 25'b10110101_01001000_11111101_0;
      patterns[46411] = 25'b10110101_01001001_11111110_0;
      patterns[46412] = 25'b10110101_01001010_11111111_0;
      patterns[46413] = 25'b10110101_01001011_00000000_1;
      patterns[46414] = 25'b10110101_01001100_00000001_1;
      patterns[46415] = 25'b10110101_01001101_00000010_1;
      patterns[46416] = 25'b10110101_01001110_00000011_1;
      patterns[46417] = 25'b10110101_01001111_00000100_1;
      patterns[46418] = 25'b10110101_01010000_00000101_1;
      patterns[46419] = 25'b10110101_01010001_00000110_1;
      patterns[46420] = 25'b10110101_01010010_00000111_1;
      patterns[46421] = 25'b10110101_01010011_00001000_1;
      patterns[46422] = 25'b10110101_01010100_00001001_1;
      patterns[46423] = 25'b10110101_01010101_00001010_1;
      patterns[46424] = 25'b10110101_01010110_00001011_1;
      patterns[46425] = 25'b10110101_01010111_00001100_1;
      patterns[46426] = 25'b10110101_01011000_00001101_1;
      patterns[46427] = 25'b10110101_01011001_00001110_1;
      patterns[46428] = 25'b10110101_01011010_00001111_1;
      patterns[46429] = 25'b10110101_01011011_00010000_1;
      patterns[46430] = 25'b10110101_01011100_00010001_1;
      patterns[46431] = 25'b10110101_01011101_00010010_1;
      patterns[46432] = 25'b10110101_01011110_00010011_1;
      patterns[46433] = 25'b10110101_01011111_00010100_1;
      patterns[46434] = 25'b10110101_01100000_00010101_1;
      patterns[46435] = 25'b10110101_01100001_00010110_1;
      patterns[46436] = 25'b10110101_01100010_00010111_1;
      patterns[46437] = 25'b10110101_01100011_00011000_1;
      patterns[46438] = 25'b10110101_01100100_00011001_1;
      patterns[46439] = 25'b10110101_01100101_00011010_1;
      patterns[46440] = 25'b10110101_01100110_00011011_1;
      patterns[46441] = 25'b10110101_01100111_00011100_1;
      patterns[46442] = 25'b10110101_01101000_00011101_1;
      patterns[46443] = 25'b10110101_01101001_00011110_1;
      patterns[46444] = 25'b10110101_01101010_00011111_1;
      patterns[46445] = 25'b10110101_01101011_00100000_1;
      patterns[46446] = 25'b10110101_01101100_00100001_1;
      patterns[46447] = 25'b10110101_01101101_00100010_1;
      patterns[46448] = 25'b10110101_01101110_00100011_1;
      patterns[46449] = 25'b10110101_01101111_00100100_1;
      patterns[46450] = 25'b10110101_01110000_00100101_1;
      patterns[46451] = 25'b10110101_01110001_00100110_1;
      patterns[46452] = 25'b10110101_01110010_00100111_1;
      patterns[46453] = 25'b10110101_01110011_00101000_1;
      patterns[46454] = 25'b10110101_01110100_00101001_1;
      patterns[46455] = 25'b10110101_01110101_00101010_1;
      patterns[46456] = 25'b10110101_01110110_00101011_1;
      patterns[46457] = 25'b10110101_01110111_00101100_1;
      patterns[46458] = 25'b10110101_01111000_00101101_1;
      patterns[46459] = 25'b10110101_01111001_00101110_1;
      patterns[46460] = 25'b10110101_01111010_00101111_1;
      patterns[46461] = 25'b10110101_01111011_00110000_1;
      patterns[46462] = 25'b10110101_01111100_00110001_1;
      patterns[46463] = 25'b10110101_01111101_00110010_1;
      patterns[46464] = 25'b10110101_01111110_00110011_1;
      patterns[46465] = 25'b10110101_01111111_00110100_1;
      patterns[46466] = 25'b10110101_10000000_00110101_1;
      patterns[46467] = 25'b10110101_10000001_00110110_1;
      patterns[46468] = 25'b10110101_10000010_00110111_1;
      patterns[46469] = 25'b10110101_10000011_00111000_1;
      patterns[46470] = 25'b10110101_10000100_00111001_1;
      patterns[46471] = 25'b10110101_10000101_00111010_1;
      patterns[46472] = 25'b10110101_10000110_00111011_1;
      patterns[46473] = 25'b10110101_10000111_00111100_1;
      patterns[46474] = 25'b10110101_10001000_00111101_1;
      patterns[46475] = 25'b10110101_10001001_00111110_1;
      patterns[46476] = 25'b10110101_10001010_00111111_1;
      patterns[46477] = 25'b10110101_10001011_01000000_1;
      patterns[46478] = 25'b10110101_10001100_01000001_1;
      patterns[46479] = 25'b10110101_10001101_01000010_1;
      patterns[46480] = 25'b10110101_10001110_01000011_1;
      patterns[46481] = 25'b10110101_10001111_01000100_1;
      patterns[46482] = 25'b10110101_10010000_01000101_1;
      patterns[46483] = 25'b10110101_10010001_01000110_1;
      patterns[46484] = 25'b10110101_10010010_01000111_1;
      patterns[46485] = 25'b10110101_10010011_01001000_1;
      patterns[46486] = 25'b10110101_10010100_01001001_1;
      patterns[46487] = 25'b10110101_10010101_01001010_1;
      patterns[46488] = 25'b10110101_10010110_01001011_1;
      patterns[46489] = 25'b10110101_10010111_01001100_1;
      patterns[46490] = 25'b10110101_10011000_01001101_1;
      patterns[46491] = 25'b10110101_10011001_01001110_1;
      patterns[46492] = 25'b10110101_10011010_01001111_1;
      patterns[46493] = 25'b10110101_10011011_01010000_1;
      patterns[46494] = 25'b10110101_10011100_01010001_1;
      patterns[46495] = 25'b10110101_10011101_01010010_1;
      patterns[46496] = 25'b10110101_10011110_01010011_1;
      patterns[46497] = 25'b10110101_10011111_01010100_1;
      patterns[46498] = 25'b10110101_10100000_01010101_1;
      patterns[46499] = 25'b10110101_10100001_01010110_1;
      patterns[46500] = 25'b10110101_10100010_01010111_1;
      patterns[46501] = 25'b10110101_10100011_01011000_1;
      patterns[46502] = 25'b10110101_10100100_01011001_1;
      patterns[46503] = 25'b10110101_10100101_01011010_1;
      patterns[46504] = 25'b10110101_10100110_01011011_1;
      patterns[46505] = 25'b10110101_10100111_01011100_1;
      patterns[46506] = 25'b10110101_10101000_01011101_1;
      patterns[46507] = 25'b10110101_10101001_01011110_1;
      patterns[46508] = 25'b10110101_10101010_01011111_1;
      patterns[46509] = 25'b10110101_10101011_01100000_1;
      patterns[46510] = 25'b10110101_10101100_01100001_1;
      patterns[46511] = 25'b10110101_10101101_01100010_1;
      patterns[46512] = 25'b10110101_10101110_01100011_1;
      patterns[46513] = 25'b10110101_10101111_01100100_1;
      patterns[46514] = 25'b10110101_10110000_01100101_1;
      patterns[46515] = 25'b10110101_10110001_01100110_1;
      patterns[46516] = 25'b10110101_10110010_01100111_1;
      patterns[46517] = 25'b10110101_10110011_01101000_1;
      patterns[46518] = 25'b10110101_10110100_01101001_1;
      patterns[46519] = 25'b10110101_10110101_01101010_1;
      patterns[46520] = 25'b10110101_10110110_01101011_1;
      patterns[46521] = 25'b10110101_10110111_01101100_1;
      patterns[46522] = 25'b10110101_10111000_01101101_1;
      patterns[46523] = 25'b10110101_10111001_01101110_1;
      patterns[46524] = 25'b10110101_10111010_01101111_1;
      patterns[46525] = 25'b10110101_10111011_01110000_1;
      patterns[46526] = 25'b10110101_10111100_01110001_1;
      patterns[46527] = 25'b10110101_10111101_01110010_1;
      patterns[46528] = 25'b10110101_10111110_01110011_1;
      patterns[46529] = 25'b10110101_10111111_01110100_1;
      patterns[46530] = 25'b10110101_11000000_01110101_1;
      patterns[46531] = 25'b10110101_11000001_01110110_1;
      patterns[46532] = 25'b10110101_11000010_01110111_1;
      patterns[46533] = 25'b10110101_11000011_01111000_1;
      patterns[46534] = 25'b10110101_11000100_01111001_1;
      patterns[46535] = 25'b10110101_11000101_01111010_1;
      patterns[46536] = 25'b10110101_11000110_01111011_1;
      patterns[46537] = 25'b10110101_11000111_01111100_1;
      patterns[46538] = 25'b10110101_11001000_01111101_1;
      patterns[46539] = 25'b10110101_11001001_01111110_1;
      patterns[46540] = 25'b10110101_11001010_01111111_1;
      patterns[46541] = 25'b10110101_11001011_10000000_1;
      patterns[46542] = 25'b10110101_11001100_10000001_1;
      patterns[46543] = 25'b10110101_11001101_10000010_1;
      patterns[46544] = 25'b10110101_11001110_10000011_1;
      patterns[46545] = 25'b10110101_11001111_10000100_1;
      patterns[46546] = 25'b10110101_11010000_10000101_1;
      patterns[46547] = 25'b10110101_11010001_10000110_1;
      patterns[46548] = 25'b10110101_11010010_10000111_1;
      patterns[46549] = 25'b10110101_11010011_10001000_1;
      patterns[46550] = 25'b10110101_11010100_10001001_1;
      patterns[46551] = 25'b10110101_11010101_10001010_1;
      patterns[46552] = 25'b10110101_11010110_10001011_1;
      patterns[46553] = 25'b10110101_11010111_10001100_1;
      patterns[46554] = 25'b10110101_11011000_10001101_1;
      patterns[46555] = 25'b10110101_11011001_10001110_1;
      patterns[46556] = 25'b10110101_11011010_10001111_1;
      patterns[46557] = 25'b10110101_11011011_10010000_1;
      patterns[46558] = 25'b10110101_11011100_10010001_1;
      patterns[46559] = 25'b10110101_11011101_10010010_1;
      patterns[46560] = 25'b10110101_11011110_10010011_1;
      patterns[46561] = 25'b10110101_11011111_10010100_1;
      patterns[46562] = 25'b10110101_11100000_10010101_1;
      patterns[46563] = 25'b10110101_11100001_10010110_1;
      patterns[46564] = 25'b10110101_11100010_10010111_1;
      patterns[46565] = 25'b10110101_11100011_10011000_1;
      patterns[46566] = 25'b10110101_11100100_10011001_1;
      patterns[46567] = 25'b10110101_11100101_10011010_1;
      patterns[46568] = 25'b10110101_11100110_10011011_1;
      patterns[46569] = 25'b10110101_11100111_10011100_1;
      patterns[46570] = 25'b10110101_11101000_10011101_1;
      patterns[46571] = 25'b10110101_11101001_10011110_1;
      patterns[46572] = 25'b10110101_11101010_10011111_1;
      patterns[46573] = 25'b10110101_11101011_10100000_1;
      patterns[46574] = 25'b10110101_11101100_10100001_1;
      patterns[46575] = 25'b10110101_11101101_10100010_1;
      patterns[46576] = 25'b10110101_11101110_10100011_1;
      patterns[46577] = 25'b10110101_11101111_10100100_1;
      patterns[46578] = 25'b10110101_11110000_10100101_1;
      patterns[46579] = 25'b10110101_11110001_10100110_1;
      patterns[46580] = 25'b10110101_11110010_10100111_1;
      patterns[46581] = 25'b10110101_11110011_10101000_1;
      patterns[46582] = 25'b10110101_11110100_10101001_1;
      patterns[46583] = 25'b10110101_11110101_10101010_1;
      patterns[46584] = 25'b10110101_11110110_10101011_1;
      patterns[46585] = 25'b10110101_11110111_10101100_1;
      patterns[46586] = 25'b10110101_11111000_10101101_1;
      patterns[46587] = 25'b10110101_11111001_10101110_1;
      patterns[46588] = 25'b10110101_11111010_10101111_1;
      patterns[46589] = 25'b10110101_11111011_10110000_1;
      patterns[46590] = 25'b10110101_11111100_10110001_1;
      patterns[46591] = 25'b10110101_11111101_10110010_1;
      patterns[46592] = 25'b10110101_11111110_10110011_1;
      patterns[46593] = 25'b10110101_11111111_10110100_1;
      patterns[46594] = 25'b10110110_00000000_10110110_0;
      patterns[46595] = 25'b10110110_00000001_10110111_0;
      patterns[46596] = 25'b10110110_00000010_10111000_0;
      patterns[46597] = 25'b10110110_00000011_10111001_0;
      patterns[46598] = 25'b10110110_00000100_10111010_0;
      patterns[46599] = 25'b10110110_00000101_10111011_0;
      patterns[46600] = 25'b10110110_00000110_10111100_0;
      patterns[46601] = 25'b10110110_00000111_10111101_0;
      patterns[46602] = 25'b10110110_00001000_10111110_0;
      patterns[46603] = 25'b10110110_00001001_10111111_0;
      patterns[46604] = 25'b10110110_00001010_11000000_0;
      patterns[46605] = 25'b10110110_00001011_11000001_0;
      patterns[46606] = 25'b10110110_00001100_11000010_0;
      patterns[46607] = 25'b10110110_00001101_11000011_0;
      patterns[46608] = 25'b10110110_00001110_11000100_0;
      patterns[46609] = 25'b10110110_00001111_11000101_0;
      patterns[46610] = 25'b10110110_00010000_11000110_0;
      patterns[46611] = 25'b10110110_00010001_11000111_0;
      patterns[46612] = 25'b10110110_00010010_11001000_0;
      patterns[46613] = 25'b10110110_00010011_11001001_0;
      patterns[46614] = 25'b10110110_00010100_11001010_0;
      patterns[46615] = 25'b10110110_00010101_11001011_0;
      patterns[46616] = 25'b10110110_00010110_11001100_0;
      patterns[46617] = 25'b10110110_00010111_11001101_0;
      patterns[46618] = 25'b10110110_00011000_11001110_0;
      patterns[46619] = 25'b10110110_00011001_11001111_0;
      patterns[46620] = 25'b10110110_00011010_11010000_0;
      patterns[46621] = 25'b10110110_00011011_11010001_0;
      patterns[46622] = 25'b10110110_00011100_11010010_0;
      patterns[46623] = 25'b10110110_00011101_11010011_0;
      patterns[46624] = 25'b10110110_00011110_11010100_0;
      patterns[46625] = 25'b10110110_00011111_11010101_0;
      patterns[46626] = 25'b10110110_00100000_11010110_0;
      patterns[46627] = 25'b10110110_00100001_11010111_0;
      patterns[46628] = 25'b10110110_00100010_11011000_0;
      patterns[46629] = 25'b10110110_00100011_11011001_0;
      patterns[46630] = 25'b10110110_00100100_11011010_0;
      patterns[46631] = 25'b10110110_00100101_11011011_0;
      patterns[46632] = 25'b10110110_00100110_11011100_0;
      patterns[46633] = 25'b10110110_00100111_11011101_0;
      patterns[46634] = 25'b10110110_00101000_11011110_0;
      patterns[46635] = 25'b10110110_00101001_11011111_0;
      patterns[46636] = 25'b10110110_00101010_11100000_0;
      patterns[46637] = 25'b10110110_00101011_11100001_0;
      patterns[46638] = 25'b10110110_00101100_11100010_0;
      patterns[46639] = 25'b10110110_00101101_11100011_0;
      patterns[46640] = 25'b10110110_00101110_11100100_0;
      patterns[46641] = 25'b10110110_00101111_11100101_0;
      patterns[46642] = 25'b10110110_00110000_11100110_0;
      patterns[46643] = 25'b10110110_00110001_11100111_0;
      patterns[46644] = 25'b10110110_00110010_11101000_0;
      patterns[46645] = 25'b10110110_00110011_11101001_0;
      patterns[46646] = 25'b10110110_00110100_11101010_0;
      patterns[46647] = 25'b10110110_00110101_11101011_0;
      patterns[46648] = 25'b10110110_00110110_11101100_0;
      patterns[46649] = 25'b10110110_00110111_11101101_0;
      patterns[46650] = 25'b10110110_00111000_11101110_0;
      patterns[46651] = 25'b10110110_00111001_11101111_0;
      patterns[46652] = 25'b10110110_00111010_11110000_0;
      patterns[46653] = 25'b10110110_00111011_11110001_0;
      patterns[46654] = 25'b10110110_00111100_11110010_0;
      patterns[46655] = 25'b10110110_00111101_11110011_0;
      patterns[46656] = 25'b10110110_00111110_11110100_0;
      patterns[46657] = 25'b10110110_00111111_11110101_0;
      patterns[46658] = 25'b10110110_01000000_11110110_0;
      patterns[46659] = 25'b10110110_01000001_11110111_0;
      patterns[46660] = 25'b10110110_01000010_11111000_0;
      patterns[46661] = 25'b10110110_01000011_11111001_0;
      patterns[46662] = 25'b10110110_01000100_11111010_0;
      patterns[46663] = 25'b10110110_01000101_11111011_0;
      patterns[46664] = 25'b10110110_01000110_11111100_0;
      patterns[46665] = 25'b10110110_01000111_11111101_0;
      patterns[46666] = 25'b10110110_01001000_11111110_0;
      patterns[46667] = 25'b10110110_01001001_11111111_0;
      patterns[46668] = 25'b10110110_01001010_00000000_1;
      patterns[46669] = 25'b10110110_01001011_00000001_1;
      patterns[46670] = 25'b10110110_01001100_00000010_1;
      patterns[46671] = 25'b10110110_01001101_00000011_1;
      patterns[46672] = 25'b10110110_01001110_00000100_1;
      patterns[46673] = 25'b10110110_01001111_00000101_1;
      patterns[46674] = 25'b10110110_01010000_00000110_1;
      patterns[46675] = 25'b10110110_01010001_00000111_1;
      patterns[46676] = 25'b10110110_01010010_00001000_1;
      patterns[46677] = 25'b10110110_01010011_00001001_1;
      patterns[46678] = 25'b10110110_01010100_00001010_1;
      patterns[46679] = 25'b10110110_01010101_00001011_1;
      patterns[46680] = 25'b10110110_01010110_00001100_1;
      patterns[46681] = 25'b10110110_01010111_00001101_1;
      patterns[46682] = 25'b10110110_01011000_00001110_1;
      patterns[46683] = 25'b10110110_01011001_00001111_1;
      patterns[46684] = 25'b10110110_01011010_00010000_1;
      patterns[46685] = 25'b10110110_01011011_00010001_1;
      patterns[46686] = 25'b10110110_01011100_00010010_1;
      patterns[46687] = 25'b10110110_01011101_00010011_1;
      patterns[46688] = 25'b10110110_01011110_00010100_1;
      patterns[46689] = 25'b10110110_01011111_00010101_1;
      patterns[46690] = 25'b10110110_01100000_00010110_1;
      patterns[46691] = 25'b10110110_01100001_00010111_1;
      patterns[46692] = 25'b10110110_01100010_00011000_1;
      patterns[46693] = 25'b10110110_01100011_00011001_1;
      patterns[46694] = 25'b10110110_01100100_00011010_1;
      patterns[46695] = 25'b10110110_01100101_00011011_1;
      patterns[46696] = 25'b10110110_01100110_00011100_1;
      patterns[46697] = 25'b10110110_01100111_00011101_1;
      patterns[46698] = 25'b10110110_01101000_00011110_1;
      patterns[46699] = 25'b10110110_01101001_00011111_1;
      patterns[46700] = 25'b10110110_01101010_00100000_1;
      patterns[46701] = 25'b10110110_01101011_00100001_1;
      patterns[46702] = 25'b10110110_01101100_00100010_1;
      patterns[46703] = 25'b10110110_01101101_00100011_1;
      patterns[46704] = 25'b10110110_01101110_00100100_1;
      patterns[46705] = 25'b10110110_01101111_00100101_1;
      patterns[46706] = 25'b10110110_01110000_00100110_1;
      patterns[46707] = 25'b10110110_01110001_00100111_1;
      patterns[46708] = 25'b10110110_01110010_00101000_1;
      patterns[46709] = 25'b10110110_01110011_00101001_1;
      patterns[46710] = 25'b10110110_01110100_00101010_1;
      patterns[46711] = 25'b10110110_01110101_00101011_1;
      patterns[46712] = 25'b10110110_01110110_00101100_1;
      patterns[46713] = 25'b10110110_01110111_00101101_1;
      patterns[46714] = 25'b10110110_01111000_00101110_1;
      patterns[46715] = 25'b10110110_01111001_00101111_1;
      patterns[46716] = 25'b10110110_01111010_00110000_1;
      patterns[46717] = 25'b10110110_01111011_00110001_1;
      patterns[46718] = 25'b10110110_01111100_00110010_1;
      patterns[46719] = 25'b10110110_01111101_00110011_1;
      patterns[46720] = 25'b10110110_01111110_00110100_1;
      patterns[46721] = 25'b10110110_01111111_00110101_1;
      patterns[46722] = 25'b10110110_10000000_00110110_1;
      patterns[46723] = 25'b10110110_10000001_00110111_1;
      patterns[46724] = 25'b10110110_10000010_00111000_1;
      patterns[46725] = 25'b10110110_10000011_00111001_1;
      patterns[46726] = 25'b10110110_10000100_00111010_1;
      patterns[46727] = 25'b10110110_10000101_00111011_1;
      patterns[46728] = 25'b10110110_10000110_00111100_1;
      patterns[46729] = 25'b10110110_10000111_00111101_1;
      patterns[46730] = 25'b10110110_10001000_00111110_1;
      patterns[46731] = 25'b10110110_10001001_00111111_1;
      patterns[46732] = 25'b10110110_10001010_01000000_1;
      patterns[46733] = 25'b10110110_10001011_01000001_1;
      patterns[46734] = 25'b10110110_10001100_01000010_1;
      patterns[46735] = 25'b10110110_10001101_01000011_1;
      patterns[46736] = 25'b10110110_10001110_01000100_1;
      patterns[46737] = 25'b10110110_10001111_01000101_1;
      patterns[46738] = 25'b10110110_10010000_01000110_1;
      patterns[46739] = 25'b10110110_10010001_01000111_1;
      patterns[46740] = 25'b10110110_10010010_01001000_1;
      patterns[46741] = 25'b10110110_10010011_01001001_1;
      patterns[46742] = 25'b10110110_10010100_01001010_1;
      patterns[46743] = 25'b10110110_10010101_01001011_1;
      patterns[46744] = 25'b10110110_10010110_01001100_1;
      patterns[46745] = 25'b10110110_10010111_01001101_1;
      patterns[46746] = 25'b10110110_10011000_01001110_1;
      patterns[46747] = 25'b10110110_10011001_01001111_1;
      patterns[46748] = 25'b10110110_10011010_01010000_1;
      patterns[46749] = 25'b10110110_10011011_01010001_1;
      patterns[46750] = 25'b10110110_10011100_01010010_1;
      patterns[46751] = 25'b10110110_10011101_01010011_1;
      patterns[46752] = 25'b10110110_10011110_01010100_1;
      patterns[46753] = 25'b10110110_10011111_01010101_1;
      patterns[46754] = 25'b10110110_10100000_01010110_1;
      patterns[46755] = 25'b10110110_10100001_01010111_1;
      patterns[46756] = 25'b10110110_10100010_01011000_1;
      patterns[46757] = 25'b10110110_10100011_01011001_1;
      patterns[46758] = 25'b10110110_10100100_01011010_1;
      patterns[46759] = 25'b10110110_10100101_01011011_1;
      patterns[46760] = 25'b10110110_10100110_01011100_1;
      patterns[46761] = 25'b10110110_10100111_01011101_1;
      patterns[46762] = 25'b10110110_10101000_01011110_1;
      patterns[46763] = 25'b10110110_10101001_01011111_1;
      patterns[46764] = 25'b10110110_10101010_01100000_1;
      patterns[46765] = 25'b10110110_10101011_01100001_1;
      patterns[46766] = 25'b10110110_10101100_01100010_1;
      patterns[46767] = 25'b10110110_10101101_01100011_1;
      patterns[46768] = 25'b10110110_10101110_01100100_1;
      patterns[46769] = 25'b10110110_10101111_01100101_1;
      patterns[46770] = 25'b10110110_10110000_01100110_1;
      patterns[46771] = 25'b10110110_10110001_01100111_1;
      patterns[46772] = 25'b10110110_10110010_01101000_1;
      patterns[46773] = 25'b10110110_10110011_01101001_1;
      patterns[46774] = 25'b10110110_10110100_01101010_1;
      patterns[46775] = 25'b10110110_10110101_01101011_1;
      patterns[46776] = 25'b10110110_10110110_01101100_1;
      patterns[46777] = 25'b10110110_10110111_01101101_1;
      patterns[46778] = 25'b10110110_10111000_01101110_1;
      patterns[46779] = 25'b10110110_10111001_01101111_1;
      patterns[46780] = 25'b10110110_10111010_01110000_1;
      patterns[46781] = 25'b10110110_10111011_01110001_1;
      patterns[46782] = 25'b10110110_10111100_01110010_1;
      patterns[46783] = 25'b10110110_10111101_01110011_1;
      patterns[46784] = 25'b10110110_10111110_01110100_1;
      patterns[46785] = 25'b10110110_10111111_01110101_1;
      patterns[46786] = 25'b10110110_11000000_01110110_1;
      patterns[46787] = 25'b10110110_11000001_01110111_1;
      patterns[46788] = 25'b10110110_11000010_01111000_1;
      patterns[46789] = 25'b10110110_11000011_01111001_1;
      patterns[46790] = 25'b10110110_11000100_01111010_1;
      patterns[46791] = 25'b10110110_11000101_01111011_1;
      patterns[46792] = 25'b10110110_11000110_01111100_1;
      patterns[46793] = 25'b10110110_11000111_01111101_1;
      patterns[46794] = 25'b10110110_11001000_01111110_1;
      patterns[46795] = 25'b10110110_11001001_01111111_1;
      patterns[46796] = 25'b10110110_11001010_10000000_1;
      patterns[46797] = 25'b10110110_11001011_10000001_1;
      patterns[46798] = 25'b10110110_11001100_10000010_1;
      patterns[46799] = 25'b10110110_11001101_10000011_1;
      patterns[46800] = 25'b10110110_11001110_10000100_1;
      patterns[46801] = 25'b10110110_11001111_10000101_1;
      patterns[46802] = 25'b10110110_11010000_10000110_1;
      patterns[46803] = 25'b10110110_11010001_10000111_1;
      patterns[46804] = 25'b10110110_11010010_10001000_1;
      patterns[46805] = 25'b10110110_11010011_10001001_1;
      patterns[46806] = 25'b10110110_11010100_10001010_1;
      patterns[46807] = 25'b10110110_11010101_10001011_1;
      patterns[46808] = 25'b10110110_11010110_10001100_1;
      patterns[46809] = 25'b10110110_11010111_10001101_1;
      patterns[46810] = 25'b10110110_11011000_10001110_1;
      patterns[46811] = 25'b10110110_11011001_10001111_1;
      patterns[46812] = 25'b10110110_11011010_10010000_1;
      patterns[46813] = 25'b10110110_11011011_10010001_1;
      patterns[46814] = 25'b10110110_11011100_10010010_1;
      patterns[46815] = 25'b10110110_11011101_10010011_1;
      patterns[46816] = 25'b10110110_11011110_10010100_1;
      patterns[46817] = 25'b10110110_11011111_10010101_1;
      patterns[46818] = 25'b10110110_11100000_10010110_1;
      patterns[46819] = 25'b10110110_11100001_10010111_1;
      patterns[46820] = 25'b10110110_11100010_10011000_1;
      patterns[46821] = 25'b10110110_11100011_10011001_1;
      patterns[46822] = 25'b10110110_11100100_10011010_1;
      patterns[46823] = 25'b10110110_11100101_10011011_1;
      patterns[46824] = 25'b10110110_11100110_10011100_1;
      patterns[46825] = 25'b10110110_11100111_10011101_1;
      patterns[46826] = 25'b10110110_11101000_10011110_1;
      patterns[46827] = 25'b10110110_11101001_10011111_1;
      patterns[46828] = 25'b10110110_11101010_10100000_1;
      patterns[46829] = 25'b10110110_11101011_10100001_1;
      patterns[46830] = 25'b10110110_11101100_10100010_1;
      patterns[46831] = 25'b10110110_11101101_10100011_1;
      patterns[46832] = 25'b10110110_11101110_10100100_1;
      patterns[46833] = 25'b10110110_11101111_10100101_1;
      patterns[46834] = 25'b10110110_11110000_10100110_1;
      patterns[46835] = 25'b10110110_11110001_10100111_1;
      patterns[46836] = 25'b10110110_11110010_10101000_1;
      patterns[46837] = 25'b10110110_11110011_10101001_1;
      patterns[46838] = 25'b10110110_11110100_10101010_1;
      patterns[46839] = 25'b10110110_11110101_10101011_1;
      patterns[46840] = 25'b10110110_11110110_10101100_1;
      patterns[46841] = 25'b10110110_11110111_10101101_1;
      patterns[46842] = 25'b10110110_11111000_10101110_1;
      patterns[46843] = 25'b10110110_11111001_10101111_1;
      patterns[46844] = 25'b10110110_11111010_10110000_1;
      patterns[46845] = 25'b10110110_11111011_10110001_1;
      patterns[46846] = 25'b10110110_11111100_10110010_1;
      patterns[46847] = 25'b10110110_11111101_10110011_1;
      patterns[46848] = 25'b10110110_11111110_10110100_1;
      patterns[46849] = 25'b10110110_11111111_10110101_1;
      patterns[46850] = 25'b10110111_00000000_10110111_0;
      patterns[46851] = 25'b10110111_00000001_10111000_0;
      patterns[46852] = 25'b10110111_00000010_10111001_0;
      patterns[46853] = 25'b10110111_00000011_10111010_0;
      patterns[46854] = 25'b10110111_00000100_10111011_0;
      patterns[46855] = 25'b10110111_00000101_10111100_0;
      patterns[46856] = 25'b10110111_00000110_10111101_0;
      patterns[46857] = 25'b10110111_00000111_10111110_0;
      patterns[46858] = 25'b10110111_00001000_10111111_0;
      patterns[46859] = 25'b10110111_00001001_11000000_0;
      patterns[46860] = 25'b10110111_00001010_11000001_0;
      patterns[46861] = 25'b10110111_00001011_11000010_0;
      patterns[46862] = 25'b10110111_00001100_11000011_0;
      patterns[46863] = 25'b10110111_00001101_11000100_0;
      patterns[46864] = 25'b10110111_00001110_11000101_0;
      patterns[46865] = 25'b10110111_00001111_11000110_0;
      patterns[46866] = 25'b10110111_00010000_11000111_0;
      patterns[46867] = 25'b10110111_00010001_11001000_0;
      patterns[46868] = 25'b10110111_00010010_11001001_0;
      patterns[46869] = 25'b10110111_00010011_11001010_0;
      patterns[46870] = 25'b10110111_00010100_11001011_0;
      patterns[46871] = 25'b10110111_00010101_11001100_0;
      patterns[46872] = 25'b10110111_00010110_11001101_0;
      patterns[46873] = 25'b10110111_00010111_11001110_0;
      patterns[46874] = 25'b10110111_00011000_11001111_0;
      patterns[46875] = 25'b10110111_00011001_11010000_0;
      patterns[46876] = 25'b10110111_00011010_11010001_0;
      patterns[46877] = 25'b10110111_00011011_11010010_0;
      patterns[46878] = 25'b10110111_00011100_11010011_0;
      patterns[46879] = 25'b10110111_00011101_11010100_0;
      patterns[46880] = 25'b10110111_00011110_11010101_0;
      patterns[46881] = 25'b10110111_00011111_11010110_0;
      patterns[46882] = 25'b10110111_00100000_11010111_0;
      patterns[46883] = 25'b10110111_00100001_11011000_0;
      patterns[46884] = 25'b10110111_00100010_11011001_0;
      patterns[46885] = 25'b10110111_00100011_11011010_0;
      patterns[46886] = 25'b10110111_00100100_11011011_0;
      patterns[46887] = 25'b10110111_00100101_11011100_0;
      patterns[46888] = 25'b10110111_00100110_11011101_0;
      patterns[46889] = 25'b10110111_00100111_11011110_0;
      patterns[46890] = 25'b10110111_00101000_11011111_0;
      patterns[46891] = 25'b10110111_00101001_11100000_0;
      patterns[46892] = 25'b10110111_00101010_11100001_0;
      patterns[46893] = 25'b10110111_00101011_11100010_0;
      patterns[46894] = 25'b10110111_00101100_11100011_0;
      patterns[46895] = 25'b10110111_00101101_11100100_0;
      patterns[46896] = 25'b10110111_00101110_11100101_0;
      patterns[46897] = 25'b10110111_00101111_11100110_0;
      patterns[46898] = 25'b10110111_00110000_11100111_0;
      patterns[46899] = 25'b10110111_00110001_11101000_0;
      patterns[46900] = 25'b10110111_00110010_11101001_0;
      patterns[46901] = 25'b10110111_00110011_11101010_0;
      patterns[46902] = 25'b10110111_00110100_11101011_0;
      patterns[46903] = 25'b10110111_00110101_11101100_0;
      patterns[46904] = 25'b10110111_00110110_11101101_0;
      patterns[46905] = 25'b10110111_00110111_11101110_0;
      patterns[46906] = 25'b10110111_00111000_11101111_0;
      patterns[46907] = 25'b10110111_00111001_11110000_0;
      patterns[46908] = 25'b10110111_00111010_11110001_0;
      patterns[46909] = 25'b10110111_00111011_11110010_0;
      patterns[46910] = 25'b10110111_00111100_11110011_0;
      patterns[46911] = 25'b10110111_00111101_11110100_0;
      patterns[46912] = 25'b10110111_00111110_11110101_0;
      patterns[46913] = 25'b10110111_00111111_11110110_0;
      patterns[46914] = 25'b10110111_01000000_11110111_0;
      patterns[46915] = 25'b10110111_01000001_11111000_0;
      patterns[46916] = 25'b10110111_01000010_11111001_0;
      patterns[46917] = 25'b10110111_01000011_11111010_0;
      patterns[46918] = 25'b10110111_01000100_11111011_0;
      patterns[46919] = 25'b10110111_01000101_11111100_0;
      patterns[46920] = 25'b10110111_01000110_11111101_0;
      patterns[46921] = 25'b10110111_01000111_11111110_0;
      patterns[46922] = 25'b10110111_01001000_11111111_0;
      patterns[46923] = 25'b10110111_01001001_00000000_1;
      patterns[46924] = 25'b10110111_01001010_00000001_1;
      patterns[46925] = 25'b10110111_01001011_00000010_1;
      patterns[46926] = 25'b10110111_01001100_00000011_1;
      patterns[46927] = 25'b10110111_01001101_00000100_1;
      patterns[46928] = 25'b10110111_01001110_00000101_1;
      patterns[46929] = 25'b10110111_01001111_00000110_1;
      patterns[46930] = 25'b10110111_01010000_00000111_1;
      patterns[46931] = 25'b10110111_01010001_00001000_1;
      patterns[46932] = 25'b10110111_01010010_00001001_1;
      patterns[46933] = 25'b10110111_01010011_00001010_1;
      patterns[46934] = 25'b10110111_01010100_00001011_1;
      patterns[46935] = 25'b10110111_01010101_00001100_1;
      patterns[46936] = 25'b10110111_01010110_00001101_1;
      patterns[46937] = 25'b10110111_01010111_00001110_1;
      patterns[46938] = 25'b10110111_01011000_00001111_1;
      patterns[46939] = 25'b10110111_01011001_00010000_1;
      patterns[46940] = 25'b10110111_01011010_00010001_1;
      patterns[46941] = 25'b10110111_01011011_00010010_1;
      patterns[46942] = 25'b10110111_01011100_00010011_1;
      patterns[46943] = 25'b10110111_01011101_00010100_1;
      patterns[46944] = 25'b10110111_01011110_00010101_1;
      patterns[46945] = 25'b10110111_01011111_00010110_1;
      patterns[46946] = 25'b10110111_01100000_00010111_1;
      patterns[46947] = 25'b10110111_01100001_00011000_1;
      patterns[46948] = 25'b10110111_01100010_00011001_1;
      patterns[46949] = 25'b10110111_01100011_00011010_1;
      patterns[46950] = 25'b10110111_01100100_00011011_1;
      patterns[46951] = 25'b10110111_01100101_00011100_1;
      patterns[46952] = 25'b10110111_01100110_00011101_1;
      patterns[46953] = 25'b10110111_01100111_00011110_1;
      patterns[46954] = 25'b10110111_01101000_00011111_1;
      patterns[46955] = 25'b10110111_01101001_00100000_1;
      patterns[46956] = 25'b10110111_01101010_00100001_1;
      patterns[46957] = 25'b10110111_01101011_00100010_1;
      patterns[46958] = 25'b10110111_01101100_00100011_1;
      patterns[46959] = 25'b10110111_01101101_00100100_1;
      patterns[46960] = 25'b10110111_01101110_00100101_1;
      patterns[46961] = 25'b10110111_01101111_00100110_1;
      patterns[46962] = 25'b10110111_01110000_00100111_1;
      patterns[46963] = 25'b10110111_01110001_00101000_1;
      patterns[46964] = 25'b10110111_01110010_00101001_1;
      patterns[46965] = 25'b10110111_01110011_00101010_1;
      patterns[46966] = 25'b10110111_01110100_00101011_1;
      patterns[46967] = 25'b10110111_01110101_00101100_1;
      patterns[46968] = 25'b10110111_01110110_00101101_1;
      patterns[46969] = 25'b10110111_01110111_00101110_1;
      patterns[46970] = 25'b10110111_01111000_00101111_1;
      patterns[46971] = 25'b10110111_01111001_00110000_1;
      patterns[46972] = 25'b10110111_01111010_00110001_1;
      patterns[46973] = 25'b10110111_01111011_00110010_1;
      patterns[46974] = 25'b10110111_01111100_00110011_1;
      patterns[46975] = 25'b10110111_01111101_00110100_1;
      patterns[46976] = 25'b10110111_01111110_00110101_1;
      patterns[46977] = 25'b10110111_01111111_00110110_1;
      patterns[46978] = 25'b10110111_10000000_00110111_1;
      patterns[46979] = 25'b10110111_10000001_00111000_1;
      patterns[46980] = 25'b10110111_10000010_00111001_1;
      patterns[46981] = 25'b10110111_10000011_00111010_1;
      patterns[46982] = 25'b10110111_10000100_00111011_1;
      patterns[46983] = 25'b10110111_10000101_00111100_1;
      patterns[46984] = 25'b10110111_10000110_00111101_1;
      patterns[46985] = 25'b10110111_10000111_00111110_1;
      patterns[46986] = 25'b10110111_10001000_00111111_1;
      patterns[46987] = 25'b10110111_10001001_01000000_1;
      patterns[46988] = 25'b10110111_10001010_01000001_1;
      patterns[46989] = 25'b10110111_10001011_01000010_1;
      patterns[46990] = 25'b10110111_10001100_01000011_1;
      patterns[46991] = 25'b10110111_10001101_01000100_1;
      patterns[46992] = 25'b10110111_10001110_01000101_1;
      patterns[46993] = 25'b10110111_10001111_01000110_1;
      patterns[46994] = 25'b10110111_10010000_01000111_1;
      patterns[46995] = 25'b10110111_10010001_01001000_1;
      patterns[46996] = 25'b10110111_10010010_01001001_1;
      patterns[46997] = 25'b10110111_10010011_01001010_1;
      patterns[46998] = 25'b10110111_10010100_01001011_1;
      patterns[46999] = 25'b10110111_10010101_01001100_1;
      patterns[47000] = 25'b10110111_10010110_01001101_1;
      patterns[47001] = 25'b10110111_10010111_01001110_1;
      patterns[47002] = 25'b10110111_10011000_01001111_1;
      patterns[47003] = 25'b10110111_10011001_01010000_1;
      patterns[47004] = 25'b10110111_10011010_01010001_1;
      patterns[47005] = 25'b10110111_10011011_01010010_1;
      patterns[47006] = 25'b10110111_10011100_01010011_1;
      patterns[47007] = 25'b10110111_10011101_01010100_1;
      patterns[47008] = 25'b10110111_10011110_01010101_1;
      patterns[47009] = 25'b10110111_10011111_01010110_1;
      patterns[47010] = 25'b10110111_10100000_01010111_1;
      patterns[47011] = 25'b10110111_10100001_01011000_1;
      patterns[47012] = 25'b10110111_10100010_01011001_1;
      patterns[47013] = 25'b10110111_10100011_01011010_1;
      patterns[47014] = 25'b10110111_10100100_01011011_1;
      patterns[47015] = 25'b10110111_10100101_01011100_1;
      patterns[47016] = 25'b10110111_10100110_01011101_1;
      patterns[47017] = 25'b10110111_10100111_01011110_1;
      patterns[47018] = 25'b10110111_10101000_01011111_1;
      patterns[47019] = 25'b10110111_10101001_01100000_1;
      patterns[47020] = 25'b10110111_10101010_01100001_1;
      patterns[47021] = 25'b10110111_10101011_01100010_1;
      patterns[47022] = 25'b10110111_10101100_01100011_1;
      patterns[47023] = 25'b10110111_10101101_01100100_1;
      patterns[47024] = 25'b10110111_10101110_01100101_1;
      patterns[47025] = 25'b10110111_10101111_01100110_1;
      patterns[47026] = 25'b10110111_10110000_01100111_1;
      patterns[47027] = 25'b10110111_10110001_01101000_1;
      patterns[47028] = 25'b10110111_10110010_01101001_1;
      patterns[47029] = 25'b10110111_10110011_01101010_1;
      patterns[47030] = 25'b10110111_10110100_01101011_1;
      patterns[47031] = 25'b10110111_10110101_01101100_1;
      patterns[47032] = 25'b10110111_10110110_01101101_1;
      patterns[47033] = 25'b10110111_10110111_01101110_1;
      patterns[47034] = 25'b10110111_10111000_01101111_1;
      patterns[47035] = 25'b10110111_10111001_01110000_1;
      patterns[47036] = 25'b10110111_10111010_01110001_1;
      patterns[47037] = 25'b10110111_10111011_01110010_1;
      patterns[47038] = 25'b10110111_10111100_01110011_1;
      patterns[47039] = 25'b10110111_10111101_01110100_1;
      patterns[47040] = 25'b10110111_10111110_01110101_1;
      patterns[47041] = 25'b10110111_10111111_01110110_1;
      patterns[47042] = 25'b10110111_11000000_01110111_1;
      patterns[47043] = 25'b10110111_11000001_01111000_1;
      patterns[47044] = 25'b10110111_11000010_01111001_1;
      patterns[47045] = 25'b10110111_11000011_01111010_1;
      patterns[47046] = 25'b10110111_11000100_01111011_1;
      patterns[47047] = 25'b10110111_11000101_01111100_1;
      patterns[47048] = 25'b10110111_11000110_01111101_1;
      patterns[47049] = 25'b10110111_11000111_01111110_1;
      patterns[47050] = 25'b10110111_11001000_01111111_1;
      patterns[47051] = 25'b10110111_11001001_10000000_1;
      patterns[47052] = 25'b10110111_11001010_10000001_1;
      patterns[47053] = 25'b10110111_11001011_10000010_1;
      patterns[47054] = 25'b10110111_11001100_10000011_1;
      patterns[47055] = 25'b10110111_11001101_10000100_1;
      patterns[47056] = 25'b10110111_11001110_10000101_1;
      patterns[47057] = 25'b10110111_11001111_10000110_1;
      patterns[47058] = 25'b10110111_11010000_10000111_1;
      patterns[47059] = 25'b10110111_11010001_10001000_1;
      patterns[47060] = 25'b10110111_11010010_10001001_1;
      patterns[47061] = 25'b10110111_11010011_10001010_1;
      patterns[47062] = 25'b10110111_11010100_10001011_1;
      patterns[47063] = 25'b10110111_11010101_10001100_1;
      patterns[47064] = 25'b10110111_11010110_10001101_1;
      patterns[47065] = 25'b10110111_11010111_10001110_1;
      patterns[47066] = 25'b10110111_11011000_10001111_1;
      patterns[47067] = 25'b10110111_11011001_10010000_1;
      patterns[47068] = 25'b10110111_11011010_10010001_1;
      patterns[47069] = 25'b10110111_11011011_10010010_1;
      patterns[47070] = 25'b10110111_11011100_10010011_1;
      patterns[47071] = 25'b10110111_11011101_10010100_1;
      patterns[47072] = 25'b10110111_11011110_10010101_1;
      patterns[47073] = 25'b10110111_11011111_10010110_1;
      patterns[47074] = 25'b10110111_11100000_10010111_1;
      patterns[47075] = 25'b10110111_11100001_10011000_1;
      patterns[47076] = 25'b10110111_11100010_10011001_1;
      patterns[47077] = 25'b10110111_11100011_10011010_1;
      patterns[47078] = 25'b10110111_11100100_10011011_1;
      patterns[47079] = 25'b10110111_11100101_10011100_1;
      patterns[47080] = 25'b10110111_11100110_10011101_1;
      patterns[47081] = 25'b10110111_11100111_10011110_1;
      patterns[47082] = 25'b10110111_11101000_10011111_1;
      patterns[47083] = 25'b10110111_11101001_10100000_1;
      patterns[47084] = 25'b10110111_11101010_10100001_1;
      patterns[47085] = 25'b10110111_11101011_10100010_1;
      patterns[47086] = 25'b10110111_11101100_10100011_1;
      patterns[47087] = 25'b10110111_11101101_10100100_1;
      patterns[47088] = 25'b10110111_11101110_10100101_1;
      patterns[47089] = 25'b10110111_11101111_10100110_1;
      patterns[47090] = 25'b10110111_11110000_10100111_1;
      patterns[47091] = 25'b10110111_11110001_10101000_1;
      patterns[47092] = 25'b10110111_11110010_10101001_1;
      patterns[47093] = 25'b10110111_11110011_10101010_1;
      patterns[47094] = 25'b10110111_11110100_10101011_1;
      patterns[47095] = 25'b10110111_11110101_10101100_1;
      patterns[47096] = 25'b10110111_11110110_10101101_1;
      patterns[47097] = 25'b10110111_11110111_10101110_1;
      patterns[47098] = 25'b10110111_11111000_10101111_1;
      patterns[47099] = 25'b10110111_11111001_10110000_1;
      patterns[47100] = 25'b10110111_11111010_10110001_1;
      patterns[47101] = 25'b10110111_11111011_10110010_1;
      patterns[47102] = 25'b10110111_11111100_10110011_1;
      patterns[47103] = 25'b10110111_11111101_10110100_1;
      patterns[47104] = 25'b10110111_11111110_10110101_1;
      patterns[47105] = 25'b10110111_11111111_10110110_1;
      patterns[47106] = 25'b10111000_00000000_10111000_0;
      patterns[47107] = 25'b10111000_00000001_10111001_0;
      patterns[47108] = 25'b10111000_00000010_10111010_0;
      patterns[47109] = 25'b10111000_00000011_10111011_0;
      patterns[47110] = 25'b10111000_00000100_10111100_0;
      patterns[47111] = 25'b10111000_00000101_10111101_0;
      patterns[47112] = 25'b10111000_00000110_10111110_0;
      patterns[47113] = 25'b10111000_00000111_10111111_0;
      patterns[47114] = 25'b10111000_00001000_11000000_0;
      patterns[47115] = 25'b10111000_00001001_11000001_0;
      patterns[47116] = 25'b10111000_00001010_11000010_0;
      patterns[47117] = 25'b10111000_00001011_11000011_0;
      patterns[47118] = 25'b10111000_00001100_11000100_0;
      patterns[47119] = 25'b10111000_00001101_11000101_0;
      patterns[47120] = 25'b10111000_00001110_11000110_0;
      patterns[47121] = 25'b10111000_00001111_11000111_0;
      patterns[47122] = 25'b10111000_00010000_11001000_0;
      patterns[47123] = 25'b10111000_00010001_11001001_0;
      patterns[47124] = 25'b10111000_00010010_11001010_0;
      patterns[47125] = 25'b10111000_00010011_11001011_0;
      patterns[47126] = 25'b10111000_00010100_11001100_0;
      patterns[47127] = 25'b10111000_00010101_11001101_0;
      patterns[47128] = 25'b10111000_00010110_11001110_0;
      patterns[47129] = 25'b10111000_00010111_11001111_0;
      patterns[47130] = 25'b10111000_00011000_11010000_0;
      patterns[47131] = 25'b10111000_00011001_11010001_0;
      patterns[47132] = 25'b10111000_00011010_11010010_0;
      patterns[47133] = 25'b10111000_00011011_11010011_0;
      patterns[47134] = 25'b10111000_00011100_11010100_0;
      patterns[47135] = 25'b10111000_00011101_11010101_0;
      patterns[47136] = 25'b10111000_00011110_11010110_0;
      patterns[47137] = 25'b10111000_00011111_11010111_0;
      patterns[47138] = 25'b10111000_00100000_11011000_0;
      patterns[47139] = 25'b10111000_00100001_11011001_0;
      patterns[47140] = 25'b10111000_00100010_11011010_0;
      patterns[47141] = 25'b10111000_00100011_11011011_0;
      patterns[47142] = 25'b10111000_00100100_11011100_0;
      patterns[47143] = 25'b10111000_00100101_11011101_0;
      patterns[47144] = 25'b10111000_00100110_11011110_0;
      patterns[47145] = 25'b10111000_00100111_11011111_0;
      patterns[47146] = 25'b10111000_00101000_11100000_0;
      patterns[47147] = 25'b10111000_00101001_11100001_0;
      patterns[47148] = 25'b10111000_00101010_11100010_0;
      patterns[47149] = 25'b10111000_00101011_11100011_0;
      patterns[47150] = 25'b10111000_00101100_11100100_0;
      patterns[47151] = 25'b10111000_00101101_11100101_0;
      patterns[47152] = 25'b10111000_00101110_11100110_0;
      patterns[47153] = 25'b10111000_00101111_11100111_0;
      patterns[47154] = 25'b10111000_00110000_11101000_0;
      patterns[47155] = 25'b10111000_00110001_11101001_0;
      patterns[47156] = 25'b10111000_00110010_11101010_0;
      patterns[47157] = 25'b10111000_00110011_11101011_0;
      patterns[47158] = 25'b10111000_00110100_11101100_0;
      patterns[47159] = 25'b10111000_00110101_11101101_0;
      patterns[47160] = 25'b10111000_00110110_11101110_0;
      patterns[47161] = 25'b10111000_00110111_11101111_0;
      patterns[47162] = 25'b10111000_00111000_11110000_0;
      patterns[47163] = 25'b10111000_00111001_11110001_0;
      patterns[47164] = 25'b10111000_00111010_11110010_0;
      patterns[47165] = 25'b10111000_00111011_11110011_0;
      patterns[47166] = 25'b10111000_00111100_11110100_0;
      patterns[47167] = 25'b10111000_00111101_11110101_0;
      patterns[47168] = 25'b10111000_00111110_11110110_0;
      patterns[47169] = 25'b10111000_00111111_11110111_0;
      patterns[47170] = 25'b10111000_01000000_11111000_0;
      patterns[47171] = 25'b10111000_01000001_11111001_0;
      patterns[47172] = 25'b10111000_01000010_11111010_0;
      patterns[47173] = 25'b10111000_01000011_11111011_0;
      patterns[47174] = 25'b10111000_01000100_11111100_0;
      patterns[47175] = 25'b10111000_01000101_11111101_0;
      patterns[47176] = 25'b10111000_01000110_11111110_0;
      patterns[47177] = 25'b10111000_01000111_11111111_0;
      patterns[47178] = 25'b10111000_01001000_00000000_1;
      patterns[47179] = 25'b10111000_01001001_00000001_1;
      patterns[47180] = 25'b10111000_01001010_00000010_1;
      patterns[47181] = 25'b10111000_01001011_00000011_1;
      patterns[47182] = 25'b10111000_01001100_00000100_1;
      patterns[47183] = 25'b10111000_01001101_00000101_1;
      patterns[47184] = 25'b10111000_01001110_00000110_1;
      patterns[47185] = 25'b10111000_01001111_00000111_1;
      patterns[47186] = 25'b10111000_01010000_00001000_1;
      patterns[47187] = 25'b10111000_01010001_00001001_1;
      patterns[47188] = 25'b10111000_01010010_00001010_1;
      patterns[47189] = 25'b10111000_01010011_00001011_1;
      patterns[47190] = 25'b10111000_01010100_00001100_1;
      patterns[47191] = 25'b10111000_01010101_00001101_1;
      patterns[47192] = 25'b10111000_01010110_00001110_1;
      patterns[47193] = 25'b10111000_01010111_00001111_1;
      patterns[47194] = 25'b10111000_01011000_00010000_1;
      patterns[47195] = 25'b10111000_01011001_00010001_1;
      patterns[47196] = 25'b10111000_01011010_00010010_1;
      patterns[47197] = 25'b10111000_01011011_00010011_1;
      patterns[47198] = 25'b10111000_01011100_00010100_1;
      patterns[47199] = 25'b10111000_01011101_00010101_1;
      patterns[47200] = 25'b10111000_01011110_00010110_1;
      patterns[47201] = 25'b10111000_01011111_00010111_1;
      patterns[47202] = 25'b10111000_01100000_00011000_1;
      patterns[47203] = 25'b10111000_01100001_00011001_1;
      patterns[47204] = 25'b10111000_01100010_00011010_1;
      patterns[47205] = 25'b10111000_01100011_00011011_1;
      patterns[47206] = 25'b10111000_01100100_00011100_1;
      patterns[47207] = 25'b10111000_01100101_00011101_1;
      patterns[47208] = 25'b10111000_01100110_00011110_1;
      patterns[47209] = 25'b10111000_01100111_00011111_1;
      patterns[47210] = 25'b10111000_01101000_00100000_1;
      patterns[47211] = 25'b10111000_01101001_00100001_1;
      patterns[47212] = 25'b10111000_01101010_00100010_1;
      patterns[47213] = 25'b10111000_01101011_00100011_1;
      patterns[47214] = 25'b10111000_01101100_00100100_1;
      patterns[47215] = 25'b10111000_01101101_00100101_1;
      patterns[47216] = 25'b10111000_01101110_00100110_1;
      patterns[47217] = 25'b10111000_01101111_00100111_1;
      patterns[47218] = 25'b10111000_01110000_00101000_1;
      patterns[47219] = 25'b10111000_01110001_00101001_1;
      patterns[47220] = 25'b10111000_01110010_00101010_1;
      patterns[47221] = 25'b10111000_01110011_00101011_1;
      patterns[47222] = 25'b10111000_01110100_00101100_1;
      patterns[47223] = 25'b10111000_01110101_00101101_1;
      patterns[47224] = 25'b10111000_01110110_00101110_1;
      patterns[47225] = 25'b10111000_01110111_00101111_1;
      patterns[47226] = 25'b10111000_01111000_00110000_1;
      patterns[47227] = 25'b10111000_01111001_00110001_1;
      patterns[47228] = 25'b10111000_01111010_00110010_1;
      patterns[47229] = 25'b10111000_01111011_00110011_1;
      patterns[47230] = 25'b10111000_01111100_00110100_1;
      patterns[47231] = 25'b10111000_01111101_00110101_1;
      patterns[47232] = 25'b10111000_01111110_00110110_1;
      patterns[47233] = 25'b10111000_01111111_00110111_1;
      patterns[47234] = 25'b10111000_10000000_00111000_1;
      patterns[47235] = 25'b10111000_10000001_00111001_1;
      patterns[47236] = 25'b10111000_10000010_00111010_1;
      patterns[47237] = 25'b10111000_10000011_00111011_1;
      patterns[47238] = 25'b10111000_10000100_00111100_1;
      patterns[47239] = 25'b10111000_10000101_00111101_1;
      patterns[47240] = 25'b10111000_10000110_00111110_1;
      patterns[47241] = 25'b10111000_10000111_00111111_1;
      patterns[47242] = 25'b10111000_10001000_01000000_1;
      patterns[47243] = 25'b10111000_10001001_01000001_1;
      patterns[47244] = 25'b10111000_10001010_01000010_1;
      patterns[47245] = 25'b10111000_10001011_01000011_1;
      patterns[47246] = 25'b10111000_10001100_01000100_1;
      patterns[47247] = 25'b10111000_10001101_01000101_1;
      patterns[47248] = 25'b10111000_10001110_01000110_1;
      patterns[47249] = 25'b10111000_10001111_01000111_1;
      patterns[47250] = 25'b10111000_10010000_01001000_1;
      patterns[47251] = 25'b10111000_10010001_01001001_1;
      patterns[47252] = 25'b10111000_10010010_01001010_1;
      patterns[47253] = 25'b10111000_10010011_01001011_1;
      patterns[47254] = 25'b10111000_10010100_01001100_1;
      patterns[47255] = 25'b10111000_10010101_01001101_1;
      patterns[47256] = 25'b10111000_10010110_01001110_1;
      patterns[47257] = 25'b10111000_10010111_01001111_1;
      patterns[47258] = 25'b10111000_10011000_01010000_1;
      patterns[47259] = 25'b10111000_10011001_01010001_1;
      patterns[47260] = 25'b10111000_10011010_01010010_1;
      patterns[47261] = 25'b10111000_10011011_01010011_1;
      patterns[47262] = 25'b10111000_10011100_01010100_1;
      patterns[47263] = 25'b10111000_10011101_01010101_1;
      patterns[47264] = 25'b10111000_10011110_01010110_1;
      patterns[47265] = 25'b10111000_10011111_01010111_1;
      patterns[47266] = 25'b10111000_10100000_01011000_1;
      patterns[47267] = 25'b10111000_10100001_01011001_1;
      patterns[47268] = 25'b10111000_10100010_01011010_1;
      patterns[47269] = 25'b10111000_10100011_01011011_1;
      patterns[47270] = 25'b10111000_10100100_01011100_1;
      patterns[47271] = 25'b10111000_10100101_01011101_1;
      patterns[47272] = 25'b10111000_10100110_01011110_1;
      patterns[47273] = 25'b10111000_10100111_01011111_1;
      patterns[47274] = 25'b10111000_10101000_01100000_1;
      patterns[47275] = 25'b10111000_10101001_01100001_1;
      patterns[47276] = 25'b10111000_10101010_01100010_1;
      patterns[47277] = 25'b10111000_10101011_01100011_1;
      patterns[47278] = 25'b10111000_10101100_01100100_1;
      patterns[47279] = 25'b10111000_10101101_01100101_1;
      patterns[47280] = 25'b10111000_10101110_01100110_1;
      patterns[47281] = 25'b10111000_10101111_01100111_1;
      patterns[47282] = 25'b10111000_10110000_01101000_1;
      patterns[47283] = 25'b10111000_10110001_01101001_1;
      patterns[47284] = 25'b10111000_10110010_01101010_1;
      patterns[47285] = 25'b10111000_10110011_01101011_1;
      patterns[47286] = 25'b10111000_10110100_01101100_1;
      patterns[47287] = 25'b10111000_10110101_01101101_1;
      patterns[47288] = 25'b10111000_10110110_01101110_1;
      patterns[47289] = 25'b10111000_10110111_01101111_1;
      patterns[47290] = 25'b10111000_10111000_01110000_1;
      patterns[47291] = 25'b10111000_10111001_01110001_1;
      patterns[47292] = 25'b10111000_10111010_01110010_1;
      patterns[47293] = 25'b10111000_10111011_01110011_1;
      patterns[47294] = 25'b10111000_10111100_01110100_1;
      patterns[47295] = 25'b10111000_10111101_01110101_1;
      patterns[47296] = 25'b10111000_10111110_01110110_1;
      patterns[47297] = 25'b10111000_10111111_01110111_1;
      patterns[47298] = 25'b10111000_11000000_01111000_1;
      patterns[47299] = 25'b10111000_11000001_01111001_1;
      patterns[47300] = 25'b10111000_11000010_01111010_1;
      patterns[47301] = 25'b10111000_11000011_01111011_1;
      patterns[47302] = 25'b10111000_11000100_01111100_1;
      patterns[47303] = 25'b10111000_11000101_01111101_1;
      patterns[47304] = 25'b10111000_11000110_01111110_1;
      patterns[47305] = 25'b10111000_11000111_01111111_1;
      patterns[47306] = 25'b10111000_11001000_10000000_1;
      patterns[47307] = 25'b10111000_11001001_10000001_1;
      patterns[47308] = 25'b10111000_11001010_10000010_1;
      patterns[47309] = 25'b10111000_11001011_10000011_1;
      patterns[47310] = 25'b10111000_11001100_10000100_1;
      patterns[47311] = 25'b10111000_11001101_10000101_1;
      patterns[47312] = 25'b10111000_11001110_10000110_1;
      patterns[47313] = 25'b10111000_11001111_10000111_1;
      patterns[47314] = 25'b10111000_11010000_10001000_1;
      patterns[47315] = 25'b10111000_11010001_10001001_1;
      patterns[47316] = 25'b10111000_11010010_10001010_1;
      patterns[47317] = 25'b10111000_11010011_10001011_1;
      patterns[47318] = 25'b10111000_11010100_10001100_1;
      patterns[47319] = 25'b10111000_11010101_10001101_1;
      patterns[47320] = 25'b10111000_11010110_10001110_1;
      patterns[47321] = 25'b10111000_11010111_10001111_1;
      patterns[47322] = 25'b10111000_11011000_10010000_1;
      patterns[47323] = 25'b10111000_11011001_10010001_1;
      patterns[47324] = 25'b10111000_11011010_10010010_1;
      patterns[47325] = 25'b10111000_11011011_10010011_1;
      patterns[47326] = 25'b10111000_11011100_10010100_1;
      patterns[47327] = 25'b10111000_11011101_10010101_1;
      patterns[47328] = 25'b10111000_11011110_10010110_1;
      patterns[47329] = 25'b10111000_11011111_10010111_1;
      patterns[47330] = 25'b10111000_11100000_10011000_1;
      patterns[47331] = 25'b10111000_11100001_10011001_1;
      patterns[47332] = 25'b10111000_11100010_10011010_1;
      patterns[47333] = 25'b10111000_11100011_10011011_1;
      patterns[47334] = 25'b10111000_11100100_10011100_1;
      patterns[47335] = 25'b10111000_11100101_10011101_1;
      patterns[47336] = 25'b10111000_11100110_10011110_1;
      patterns[47337] = 25'b10111000_11100111_10011111_1;
      patterns[47338] = 25'b10111000_11101000_10100000_1;
      patterns[47339] = 25'b10111000_11101001_10100001_1;
      patterns[47340] = 25'b10111000_11101010_10100010_1;
      patterns[47341] = 25'b10111000_11101011_10100011_1;
      patterns[47342] = 25'b10111000_11101100_10100100_1;
      patterns[47343] = 25'b10111000_11101101_10100101_1;
      patterns[47344] = 25'b10111000_11101110_10100110_1;
      patterns[47345] = 25'b10111000_11101111_10100111_1;
      patterns[47346] = 25'b10111000_11110000_10101000_1;
      patterns[47347] = 25'b10111000_11110001_10101001_1;
      patterns[47348] = 25'b10111000_11110010_10101010_1;
      patterns[47349] = 25'b10111000_11110011_10101011_1;
      patterns[47350] = 25'b10111000_11110100_10101100_1;
      patterns[47351] = 25'b10111000_11110101_10101101_1;
      patterns[47352] = 25'b10111000_11110110_10101110_1;
      patterns[47353] = 25'b10111000_11110111_10101111_1;
      patterns[47354] = 25'b10111000_11111000_10110000_1;
      patterns[47355] = 25'b10111000_11111001_10110001_1;
      patterns[47356] = 25'b10111000_11111010_10110010_1;
      patterns[47357] = 25'b10111000_11111011_10110011_1;
      patterns[47358] = 25'b10111000_11111100_10110100_1;
      patterns[47359] = 25'b10111000_11111101_10110101_1;
      patterns[47360] = 25'b10111000_11111110_10110110_1;
      patterns[47361] = 25'b10111000_11111111_10110111_1;
      patterns[47362] = 25'b10111001_00000000_10111001_0;
      patterns[47363] = 25'b10111001_00000001_10111010_0;
      patterns[47364] = 25'b10111001_00000010_10111011_0;
      patterns[47365] = 25'b10111001_00000011_10111100_0;
      patterns[47366] = 25'b10111001_00000100_10111101_0;
      patterns[47367] = 25'b10111001_00000101_10111110_0;
      patterns[47368] = 25'b10111001_00000110_10111111_0;
      patterns[47369] = 25'b10111001_00000111_11000000_0;
      patterns[47370] = 25'b10111001_00001000_11000001_0;
      patterns[47371] = 25'b10111001_00001001_11000010_0;
      patterns[47372] = 25'b10111001_00001010_11000011_0;
      patterns[47373] = 25'b10111001_00001011_11000100_0;
      patterns[47374] = 25'b10111001_00001100_11000101_0;
      patterns[47375] = 25'b10111001_00001101_11000110_0;
      patterns[47376] = 25'b10111001_00001110_11000111_0;
      patterns[47377] = 25'b10111001_00001111_11001000_0;
      patterns[47378] = 25'b10111001_00010000_11001001_0;
      patterns[47379] = 25'b10111001_00010001_11001010_0;
      patterns[47380] = 25'b10111001_00010010_11001011_0;
      patterns[47381] = 25'b10111001_00010011_11001100_0;
      patterns[47382] = 25'b10111001_00010100_11001101_0;
      patterns[47383] = 25'b10111001_00010101_11001110_0;
      patterns[47384] = 25'b10111001_00010110_11001111_0;
      patterns[47385] = 25'b10111001_00010111_11010000_0;
      patterns[47386] = 25'b10111001_00011000_11010001_0;
      patterns[47387] = 25'b10111001_00011001_11010010_0;
      patterns[47388] = 25'b10111001_00011010_11010011_0;
      patterns[47389] = 25'b10111001_00011011_11010100_0;
      patterns[47390] = 25'b10111001_00011100_11010101_0;
      patterns[47391] = 25'b10111001_00011101_11010110_0;
      patterns[47392] = 25'b10111001_00011110_11010111_0;
      patterns[47393] = 25'b10111001_00011111_11011000_0;
      patterns[47394] = 25'b10111001_00100000_11011001_0;
      patterns[47395] = 25'b10111001_00100001_11011010_0;
      patterns[47396] = 25'b10111001_00100010_11011011_0;
      patterns[47397] = 25'b10111001_00100011_11011100_0;
      patterns[47398] = 25'b10111001_00100100_11011101_0;
      patterns[47399] = 25'b10111001_00100101_11011110_0;
      patterns[47400] = 25'b10111001_00100110_11011111_0;
      patterns[47401] = 25'b10111001_00100111_11100000_0;
      patterns[47402] = 25'b10111001_00101000_11100001_0;
      patterns[47403] = 25'b10111001_00101001_11100010_0;
      patterns[47404] = 25'b10111001_00101010_11100011_0;
      patterns[47405] = 25'b10111001_00101011_11100100_0;
      patterns[47406] = 25'b10111001_00101100_11100101_0;
      patterns[47407] = 25'b10111001_00101101_11100110_0;
      patterns[47408] = 25'b10111001_00101110_11100111_0;
      patterns[47409] = 25'b10111001_00101111_11101000_0;
      patterns[47410] = 25'b10111001_00110000_11101001_0;
      patterns[47411] = 25'b10111001_00110001_11101010_0;
      patterns[47412] = 25'b10111001_00110010_11101011_0;
      patterns[47413] = 25'b10111001_00110011_11101100_0;
      patterns[47414] = 25'b10111001_00110100_11101101_0;
      patterns[47415] = 25'b10111001_00110101_11101110_0;
      patterns[47416] = 25'b10111001_00110110_11101111_0;
      patterns[47417] = 25'b10111001_00110111_11110000_0;
      patterns[47418] = 25'b10111001_00111000_11110001_0;
      patterns[47419] = 25'b10111001_00111001_11110010_0;
      patterns[47420] = 25'b10111001_00111010_11110011_0;
      patterns[47421] = 25'b10111001_00111011_11110100_0;
      patterns[47422] = 25'b10111001_00111100_11110101_0;
      patterns[47423] = 25'b10111001_00111101_11110110_0;
      patterns[47424] = 25'b10111001_00111110_11110111_0;
      patterns[47425] = 25'b10111001_00111111_11111000_0;
      patterns[47426] = 25'b10111001_01000000_11111001_0;
      patterns[47427] = 25'b10111001_01000001_11111010_0;
      patterns[47428] = 25'b10111001_01000010_11111011_0;
      patterns[47429] = 25'b10111001_01000011_11111100_0;
      patterns[47430] = 25'b10111001_01000100_11111101_0;
      patterns[47431] = 25'b10111001_01000101_11111110_0;
      patterns[47432] = 25'b10111001_01000110_11111111_0;
      patterns[47433] = 25'b10111001_01000111_00000000_1;
      patterns[47434] = 25'b10111001_01001000_00000001_1;
      patterns[47435] = 25'b10111001_01001001_00000010_1;
      patterns[47436] = 25'b10111001_01001010_00000011_1;
      patterns[47437] = 25'b10111001_01001011_00000100_1;
      patterns[47438] = 25'b10111001_01001100_00000101_1;
      patterns[47439] = 25'b10111001_01001101_00000110_1;
      patterns[47440] = 25'b10111001_01001110_00000111_1;
      patterns[47441] = 25'b10111001_01001111_00001000_1;
      patterns[47442] = 25'b10111001_01010000_00001001_1;
      patterns[47443] = 25'b10111001_01010001_00001010_1;
      patterns[47444] = 25'b10111001_01010010_00001011_1;
      patterns[47445] = 25'b10111001_01010011_00001100_1;
      patterns[47446] = 25'b10111001_01010100_00001101_1;
      patterns[47447] = 25'b10111001_01010101_00001110_1;
      patterns[47448] = 25'b10111001_01010110_00001111_1;
      patterns[47449] = 25'b10111001_01010111_00010000_1;
      patterns[47450] = 25'b10111001_01011000_00010001_1;
      patterns[47451] = 25'b10111001_01011001_00010010_1;
      patterns[47452] = 25'b10111001_01011010_00010011_1;
      patterns[47453] = 25'b10111001_01011011_00010100_1;
      patterns[47454] = 25'b10111001_01011100_00010101_1;
      patterns[47455] = 25'b10111001_01011101_00010110_1;
      patterns[47456] = 25'b10111001_01011110_00010111_1;
      patterns[47457] = 25'b10111001_01011111_00011000_1;
      patterns[47458] = 25'b10111001_01100000_00011001_1;
      patterns[47459] = 25'b10111001_01100001_00011010_1;
      patterns[47460] = 25'b10111001_01100010_00011011_1;
      patterns[47461] = 25'b10111001_01100011_00011100_1;
      patterns[47462] = 25'b10111001_01100100_00011101_1;
      patterns[47463] = 25'b10111001_01100101_00011110_1;
      patterns[47464] = 25'b10111001_01100110_00011111_1;
      patterns[47465] = 25'b10111001_01100111_00100000_1;
      patterns[47466] = 25'b10111001_01101000_00100001_1;
      patterns[47467] = 25'b10111001_01101001_00100010_1;
      patterns[47468] = 25'b10111001_01101010_00100011_1;
      patterns[47469] = 25'b10111001_01101011_00100100_1;
      patterns[47470] = 25'b10111001_01101100_00100101_1;
      patterns[47471] = 25'b10111001_01101101_00100110_1;
      patterns[47472] = 25'b10111001_01101110_00100111_1;
      patterns[47473] = 25'b10111001_01101111_00101000_1;
      patterns[47474] = 25'b10111001_01110000_00101001_1;
      patterns[47475] = 25'b10111001_01110001_00101010_1;
      patterns[47476] = 25'b10111001_01110010_00101011_1;
      patterns[47477] = 25'b10111001_01110011_00101100_1;
      patterns[47478] = 25'b10111001_01110100_00101101_1;
      patterns[47479] = 25'b10111001_01110101_00101110_1;
      patterns[47480] = 25'b10111001_01110110_00101111_1;
      patterns[47481] = 25'b10111001_01110111_00110000_1;
      patterns[47482] = 25'b10111001_01111000_00110001_1;
      patterns[47483] = 25'b10111001_01111001_00110010_1;
      patterns[47484] = 25'b10111001_01111010_00110011_1;
      patterns[47485] = 25'b10111001_01111011_00110100_1;
      patterns[47486] = 25'b10111001_01111100_00110101_1;
      patterns[47487] = 25'b10111001_01111101_00110110_1;
      patterns[47488] = 25'b10111001_01111110_00110111_1;
      patterns[47489] = 25'b10111001_01111111_00111000_1;
      patterns[47490] = 25'b10111001_10000000_00111001_1;
      patterns[47491] = 25'b10111001_10000001_00111010_1;
      patterns[47492] = 25'b10111001_10000010_00111011_1;
      patterns[47493] = 25'b10111001_10000011_00111100_1;
      patterns[47494] = 25'b10111001_10000100_00111101_1;
      patterns[47495] = 25'b10111001_10000101_00111110_1;
      patterns[47496] = 25'b10111001_10000110_00111111_1;
      patterns[47497] = 25'b10111001_10000111_01000000_1;
      patterns[47498] = 25'b10111001_10001000_01000001_1;
      patterns[47499] = 25'b10111001_10001001_01000010_1;
      patterns[47500] = 25'b10111001_10001010_01000011_1;
      patterns[47501] = 25'b10111001_10001011_01000100_1;
      patterns[47502] = 25'b10111001_10001100_01000101_1;
      patterns[47503] = 25'b10111001_10001101_01000110_1;
      patterns[47504] = 25'b10111001_10001110_01000111_1;
      patterns[47505] = 25'b10111001_10001111_01001000_1;
      patterns[47506] = 25'b10111001_10010000_01001001_1;
      patterns[47507] = 25'b10111001_10010001_01001010_1;
      patterns[47508] = 25'b10111001_10010010_01001011_1;
      patterns[47509] = 25'b10111001_10010011_01001100_1;
      patterns[47510] = 25'b10111001_10010100_01001101_1;
      patterns[47511] = 25'b10111001_10010101_01001110_1;
      patterns[47512] = 25'b10111001_10010110_01001111_1;
      patterns[47513] = 25'b10111001_10010111_01010000_1;
      patterns[47514] = 25'b10111001_10011000_01010001_1;
      patterns[47515] = 25'b10111001_10011001_01010010_1;
      patterns[47516] = 25'b10111001_10011010_01010011_1;
      patterns[47517] = 25'b10111001_10011011_01010100_1;
      patterns[47518] = 25'b10111001_10011100_01010101_1;
      patterns[47519] = 25'b10111001_10011101_01010110_1;
      patterns[47520] = 25'b10111001_10011110_01010111_1;
      patterns[47521] = 25'b10111001_10011111_01011000_1;
      patterns[47522] = 25'b10111001_10100000_01011001_1;
      patterns[47523] = 25'b10111001_10100001_01011010_1;
      patterns[47524] = 25'b10111001_10100010_01011011_1;
      patterns[47525] = 25'b10111001_10100011_01011100_1;
      patterns[47526] = 25'b10111001_10100100_01011101_1;
      patterns[47527] = 25'b10111001_10100101_01011110_1;
      patterns[47528] = 25'b10111001_10100110_01011111_1;
      patterns[47529] = 25'b10111001_10100111_01100000_1;
      patterns[47530] = 25'b10111001_10101000_01100001_1;
      patterns[47531] = 25'b10111001_10101001_01100010_1;
      patterns[47532] = 25'b10111001_10101010_01100011_1;
      patterns[47533] = 25'b10111001_10101011_01100100_1;
      patterns[47534] = 25'b10111001_10101100_01100101_1;
      patterns[47535] = 25'b10111001_10101101_01100110_1;
      patterns[47536] = 25'b10111001_10101110_01100111_1;
      patterns[47537] = 25'b10111001_10101111_01101000_1;
      patterns[47538] = 25'b10111001_10110000_01101001_1;
      patterns[47539] = 25'b10111001_10110001_01101010_1;
      patterns[47540] = 25'b10111001_10110010_01101011_1;
      patterns[47541] = 25'b10111001_10110011_01101100_1;
      patterns[47542] = 25'b10111001_10110100_01101101_1;
      patterns[47543] = 25'b10111001_10110101_01101110_1;
      patterns[47544] = 25'b10111001_10110110_01101111_1;
      patterns[47545] = 25'b10111001_10110111_01110000_1;
      patterns[47546] = 25'b10111001_10111000_01110001_1;
      patterns[47547] = 25'b10111001_10111001_01110010_1;
      patterns[47548] = 25'b10111001_10111010_01110011_1;
      patterns[47549] = 25'b10111001_10111011_01110100_1;
      patterns[47550] = 25'b10111001_10111100_01110101_1;
      patterns[47551] = 25'b10111001_10111101_01110110_1;
      patterns[47552] = 25'b10111001_10111110_01110111_1;
      patterns[47553] = 25'b10111001_10111111_01111000_1;
      patterns[47554] = 25'b10111001_11000000_01111001_1;
      patterns[47555] = 25'b10111001_11000001_01111010_1;
      patterns[47556] = 25'b10111001_11000010_01111011_1;
      patterns[47557] = 25'b10111001_11000011_01111100_1;
      patterns[47558] = 25'b10111001_11000100_01111101_1;
      patterns[47559] = 25'b10111001_11000101_01111110_1;
      patterns[47560] = 25'b10111001_11000110_01111111_1;
      patterns[47561] = 25'b10111001_11000111_10000000_1;
      patterns[47562] = 25'b10111001_11001000_10000001_1;
      patterns[47563] = 25'b10111001_11001001_10000010_1;
      patterns[47564] = 25'b10111001_11001010_10000011_1;
      patterns[47565] = 25'b10111001_11001011_10000100_1;
      patterns[47566] = 25'b10111001_11001100_10000101_1;
      patterns[47567] = 25'b10111001_11001101_10000110_1;
      patterns[47568] = 25'b10111001_11001110_10000111_1;
      patterns[47569] = 25'b10111001_11001111_10001000_1;
      patterns[47570] = 25'b10111001_11010000_10001001_1;
      patterns[47571] = 25'b10111001_11010001_10001010_1;
      patterns[47572] = 25'b10111001_11010010_10001011_1;
      patterns[47573] = 25'b10111001_11010011_10001100_1;
      patterns[47574] = 25'b10111001_11010100_10001101_1;
      patterns[47575] = 25'b10111001_11010101_10001110_1;
      patterns[47576] = 25'b10111001_11010110_10001111_1;
      patterns[47577] = 25'b10111001_11010111_10010000_1;
      patterns[47578] = 25'b10111001_11011000_10010001_1;
      patterns[47579] = 25'b10111001_11011001_10010010_1;
      patterns[47580] = 25'b10111001_11011010_10010011_1;
      patterns[47581] = 25'b10111001_11011011_10010100_1;
      patterns[47582] = 25'b10111001_11011100_10010101_1;
      patterns[47583] = 25'b10111001_11011101_10010110_1;
      patterns[47584] = 25'b10111001_11011110_10010111_1;
      patterns[47585] = 25'b10111001_11011111_10011000_1;
      patterns[47586] = 25'b10111001_11100000_10011001_1;
      patterns[47587] = 25'b10111001_11100001_10011010_1;
      patterns[47588] = 25'b10111001_11100010_10011011_1;
      patterns[47589] = 25'b10111001_11100011_10011100_1;
      patterns[47590] = 25'b10111001_11100100_10011101_1;
      patterns[47591] = 25'b10111001_11100101_10011110_1;
      patterns[47592] = 25'b10111001_11100110_10011111_1;
      patterns[47593] = 25'b10111001_11100111_10100000_1;
      patterns[47594] = 25'b10111001_11101000_10100001_1;
      patterns[47595] = 25'b10111001_11101001_10100010_1;
      patterns[47596] = 25'b10111001_11101010_10100011_1;
      patterns[47597] = 25'b10111001_11101011_10100100_1;
      patterns[47598] = 25'b10111001_11101100_10100101_1;
      patterns[47599] = 25'b10111001_11101101_10100110_1;
      patterns[47600] = 25'b10111001_11101110_10100111_1;
      patterns[47601] = 25'b10111001_11101111_10101000_1;
      patterns[47602] = 25'b10111001_11110000_10101001_1;
      patterns[47603] = 25'b10111001_11110001_10101010_1;
      patterns[47604] = 25'b10111001_11110010_10101011_1;
      patterns[47605] = 25'b10111001_11110011_10101100_1;
      patterns[47606] = 25'b10111001_11110100_10101101_1;
      patterns[47607] = 25'b10111001_11110101_10101110_1;
      patterns[47608] = 25'b10111001_11110110_10101111_1;
      patterns[47609] = 25'b10111001_11110111_10110000_1;
      patterns[47610] = 25'b10111001_11111000_10110001_1;
      patterns[47611] = 25'b10111001_11111001_10110010_1;
      patterns[47612] = 25'b10111001_11111010_10110011_1;
      patterns[47613] = 25'b10111001_11111011_10110100_1;
      patterns[47614] = 25'b10111001_11111100_10110101_1;
      patterns[47615] = 25'b10111001_11111101_10110110_1;
      patterns[47616] = 25'b10111001_11111110_10110111_1;
      patterns[47617] = 25'b10111001_11111111_10111000_1;
      patterns[47618] = 25'b10111010_00000000_10111010_0;
      patterns[47619] = 25'b10111010_00000001_10111011_0;
      patterns[47620] = 25'b10111010_00000010_10111100_0;
      patterns[47621] = 25'b10111010_00000011_10111101_0;
      patterns[47622] = 25'b10111010_00000100_10111110_0;
      patterns[47623] = 25'b10111010_00000101_10111111_0;
      patterns[47624] = 25'b10111010_00000110_11000000_0;
      patterns[47625] = 25'b10111010_00000111_11000001_0;
      patterns[47626] = 25'b10111010_00001000_11000010_0;
      patterns[47627] = 25'b10111010_00001001_11000011_0;
      patterns[47628] = 25'b10111010_00001010_11000100_0;
      patterns[47629] = 25'b10111010_00001011_11000101_0;
      patterns[47630] = 25'b10111010_00001100_11000110_0;
      patterns[47631] = 25'b10111010_00001101_11000111_0;
      patterns[47632] = 25'b10111010_00001110_11001000_0;
      patterns[47633] = 25'b10111010_00001111_11001001_0;
      patterns[47634] = 25'b10111010_00010000_11001010_0;
      patterns[47635] = 25'b10111010_00010001_11001011_0;
      patterns[47636] = 25'b10111010_00010010_11001100_0;
      patterns[47637] = 25'b10111010_00010011_11001101_0;
      patterns[47638] = 25'b10111010_00010100_11001110_0;
      patterns[47639] = 25'b10111010_00010101_11001111_0;
      patterns[47640] = 25'b10111010_00010110_11010000_0;
      patterns[47641] = 25'b10111010_00010111_11010001_0;
      patterns[47642] = 25'b10111010_00011000_11010010_0;
      patterns[47643] = 25'b10111010_00011001_11010011_0;
      patterns[47644] = 25'b10111010_00011010_11010100_0;
      patterns[47645] = 25'b10111010_00011011_11010101_0;
      patterns[47646] = 25'b10111010_00011100_11010110_0;
      patterns[47647] = 25'b10111010_00011101_11010111_0;
      patterns[47648] = 25'b10111010_00011110_11011000_0;
      patterns[47649] = 25'b10111010_00011111_11011001_0;
      patterns[47650] = 25'b10111010_00100000_11011010_0;
      patterns[47651] = 25'b10111010_00100001_11011011_0;
      patterns[47652] = 25'b10111010_00100010_11011100_0;
      patterns[47653] = 25'b10111010_00100011_11011101_0;
      patterns[47654] = 25'b10111010_00100100_11011110_0;
      patterns[47655] = 25'b10111010_00100101_11011111_0;
      patterns[47656] = 25'b10111010_00100110_11100000_0;
      patterns[47657] = 25'b10111010_00100111_11100001_0;
      patterns[47658] = 25'b10111010_00101000_11100010_0;
      patterns[47659] = 25'b10111010_00101001_11100011_0;
      patterns[47660] = 25'b10111010_00101010_11100100_0;
      patterns[47661] = 25'b10111010_00101011_11100101_0;
      patterns[47662] = 25'b10111010_00101100_11100110_0;
      patterns[47663] = 25'b10111010_00101101_11100111_0;
      patterns[47664] = 25'b10111010_00101110_11101000_0;
      patterns[47665] = 25'b10111010_00101111_11101001_0;
      patterns[47666] = 25'b10111010_00110000_11101010_0;
      patterns[47667] = 25'b10111010_00110001_11101011_0;
      patterns[47668] = 25'b10111010_00110010_11101100_0;
      patterns[47669] = 25'b10111010_00110011_11101101_0;
      patterns[47670] = 25'b10111010_00110100_11101110_0;
      patterns[47671] = 25'b10111010_00110101_11101111_0;
      patterns[47672] = 25'b10111010_00110110_11110000_0;
      patterns[47673] = 25'b10111010_00110111_11110001_0;
      patterns[47674] = 25'b10111010_00111000_11110010_0;
      patterns[47675] = 25'b10111010_00111001_11110011_0;
      patterns[47676] = 25'b10111010_00111010_11110100_0;
      patterns[47677] = 25'b10111010_00111011_11110101_0;
      patterns[47678] = 25'b10111010_00111100_11110110_0;
      patterns[47679] = 25'b10111010_00111101_11110111_0;
      patterns[47680] = 25'b10111010_00111110_11111000_0;
      patterns[47681] = 25'b10111010_00111111_11111001_0;
      patterns[47682] = 25'b10111010_01000000_11111010_0;
      patterns[47683] = 25'b10111010_01000001_11111011_0;
      patterns[47684] = 25'b10111010_01000010_11111100_0;
      patterns[47685] = 25'b10111010_01000011_11111101_0;
      patterns[47686] = 25'b10111010_01000100_11111110_0;
      patterns[47687] = 25'b10111010_01000101_11111111_0;
      patterns[47688] = 25'b10111010_01000110_00000000_1;
      patterns[47689] = 25'b10111010_01000111_00000001_1;
      patterns[47690] = 25'b10111010_01001000_00000010_1;
      patterns[47691] = 25'b10111010_01001001_00000011_1;
      patterns[47692] = 25'b10111010_01001010_00000100_1;
      patterns[47693] = 25'b10111010_01001011_00000101_1;
      patterns[47694] = 25'b10111010_01001100_00000110_1;
      patterns[47695] = 25'b10111010_01001101_00000111_1;
      patterns[47696] = 25'b10111010_01001110_00001000_1;
      patterns[47697] = 25'b10111010_01001111_00001001_1;
      patterns[47698] = 25'b10111010_01010000_00001010_1;
      patterns[47699] = 25'b10111010_01010001_00001011_1;
      patterns[47700] = 25'b10111010_01010010_00001100_1;
      patterns[47701] = 25'b10111010_01010011_00001101_1;
      patterns[47702] = 25'b10111010_01010100_00001110_1;
      patterns[47703] = 25'b10111010_01010101_00001111_1;
      patterns[47704] = 25'b10111010_01010110_00010000_1;
      patterns[47705] = 25'b10111010_01010111_00010001_1;
      patterns[47706] = 25'b10111010_01011000_00010010_1;
      patterns[47707] = 25'b10111010_01011001_00010011_1;
      patterns[47708] = 25'b10111010_01011010_00010100_1;
      patterns[47709] = 25'b10111010_01011011_00010101_1;
      patterns[47710] = 25'b10111010_01011100_00010110_1;
      patterns[47711] = 25'b10111010_01011101_00010111_1;
      patterns[47712] = 25'b10111010_01011110_00011000_1;
      patterns[47713] = 25'b10111010_01011111_00011001_1;
      patterns[47714] = 25'b10111010_01100000_00011010_1;
      patterns[47715] = 25'b10111010_01100001_00011011_1;
      patterns[47716] = 25'b10111010_01100010_00011100_1;
      patterns[47717] = 25'b10111010_01100011_00011101_1;
      patterns[47718] = 25'b10111010_01100100_00011110_1;
      patterns[47719] = 25'b10111010_01100101_00011111_1;
      patterns[47720] = 25'b10111010_01100110_00100000_1;
      patterns[47721] = 25'b10111010_01100111_00100001_1;
      patterns[47722] = 25'b10111010_01101000_00100010_1;
      patterns[47723] = 25'b10111010_01101001_00100011_1;
      patterns[47724] = 25'b10111010_01101010_00100100_1;
      patterns[47725] = 25'b10111010_01101011_00100101_1;
      patterns[47726] = 25'b10111010_01101100_00100110_1;
      patterns[47727] = 25'b10111010_01101101_00100111_1;
      patterns[47728] = 25'b10111010_01101110_00101000_1;
      patterns[47729] = 25'b10111010_01101111_00101001_1;
      patterns[47730] = 25'b10111010_01110000_00101010_1;
      patterns[47731] = 25'b10111010_01110001_00101011_1;
      patterns[47732] = 25'b10111010_01110010_00101100_1;
      patterns[47733] = 25'b10111010_01110011_00101101_1;
      patterns[47734] = 25'b10111010_01110100_00101110_1;
      patterns[47735] = 25'b10111010_01110101_00101111_1;
      patterns[47736] = 25'b10111010_01110110_00110000_1;
      patterns[47737] = 25'b10111010_01110111_00110001_1;
      patterns[47738] = 25'b10111010_01111000_00110010_1;
      patterns[47739] = 25'b10111010_01111001_00110011_1;
      patterns[47740] = 25'b10111010_01111010_00110100_1;
      patterns[47741] = 25'b10111010_01111011_00110101_1;
      patterns[47742] = 25'b10111010_01111100_00110110_1;
      patterns[47743] = 25'b10111010_01111101_00110111_1;
      patterns[47744] = 25'b10111010_01111110_00111000_1;
      patterns[47745] = 25'b10111010_01111111_00111001_1;
      patterns[47746] = 25'b10111010_10000000_00111010_1;
      patterns[47747] = 25'b10111010_10000001_00111011_1;
      patterns[47748] = 25'b10111010_10000010_00111100_1;
      patterns[47749] = 25'b10111010_10000011_00111101_1;
      patterns[47750] = 25'b10111010_10000100_00111110_1;
      patterns[47751] = 25'b10111010_10000101_00111111_1;
      patterns[47752] = 25'b10111010_10000110_01000000_1;
      patterns[47753] = 25'b10111010_10000111_01000001_1;
      patterns[47754] = 25'b10111010_10001000_01000010_1;
      patterns[47755] = 25'b10111010_10001001_01000011_1;
      patterns[47756] = 25'b10111010_10001010_01000100_1;
      patterns[47757] = 25'b10111010_10001011_01000101_1;
      patterns[47758] = 25'b10111010_10001100_01000110_1;
      patterns[47759] = 25'b10111010_10001101_01000111_1;
      patterns[47760] = 25'b10111010_10001110_01001000_1;
      patterns[47761] = 25'b10111010_10001111_01001001_1;
      patterns[47762] = 25'b10111010_10010000_01001010_1;
      patterns[47763] = 25'b10111010_10010001_01001011_1;
      patterns[47764] = 25'b10111010_10010010_01001100_1;
      patterns[47765] = 25'b10111010_10010011_01001101_1;
      patterns[47766] = 25'b10111010_10010100_01001110_1;
      patterns[47767] = 25'b10111010_10010101_01001111_1;
      patterns[47768] = 25'b10111010_10010110_01010000_1;
      patterns[47769] = 25'b10111010_10010111_01010001_1;
      patterns[47770] = 25'b10111010_10011000_01010010_1;
      patterns[47771] = 25'b10111010_10011001_01010011_1;
      patterns[47772] = 25'b10111010_10011010_01010100_1;
      patterns[47773] = 25'b10111010_10011011_01010101_1;
      patterns[47774] = 25'b10111010_10011100_01010110_1;
      patterns[47775] = 25'b10111010_10011101_01010111_1;
      patterns[47776] = 25'b10111010_10011110_01011000_1;
      patterns[47777] = 25'b10111010_10011111_01011001_1;
      patterns[47778] = 25'b10111010_10100000_01011010_1;
      patterns[47779] = 25'b10111010_10100001_01011011_1;
      patterns[47780] = 25'b10111010_10100010_01011100_1;
      patterns[47781] = 25'b10111010_10100011_01011101_1;
      patterns[47782] = 25'b10111010_10100100_01011110_1;
      patterns[47783] = 25'b10111010_10100101_01011111_1;
      patterns[47784] = 25'b10111010_10100110_01100000_1;
      patterns[47785] = 25'b10111010_10100111_01100001_1;
      patterns[47786] = 25'b10111010_10101000_01100010_1;
      patterns[47787] = 25'b10111010_10101001_01100011_1;
      patterns[47788] = 25'b10111010_10101010_01100100_1;
      patterns[47789] = 25'b10111010_10101011_01100101_1;
      patterns[47790] = 25'b10111010_10101100_01100110_1;
      patterns[47791] = 25'b10111010_10101101_01100111_1;
      patterns[47792] = 25'b10111010_10101110_01101000_1;
      patterns[47793] = 25'b10111010_10101111_01101001_1;
      patterns[47794] = 25'b10111010_10110000_01101010_1;
      patterns[47795] = 25'b10111010_10110001_01101011_1;
      patterns[47796] = 25'b10111010_10110010_01101100_1;
      patterns[47797] = 25'b10111010_10110011_01101101_1;
      patterns[47798] = 25'b10111010_10110100_01101110_1;
      patterns[47799] = 25'b10111010_10110101_01101111_1;
      patterns[47800] = 25'b10111010_10110110_01110000_1;
      patterns[47801] = 25'b10111010_10110111_01110001_1;
      patterns[47802] = 25'b10111010_10111000_01110010_1;
      patterns[47803] = 25'b10111010_10111001_01110011_1;
      patterns[47804] = 25'b10111010_10111010_01110100_1;
      patterns[47805] = 25'b10111010_10111011_01110101_1;
      patterns[47806] = 25'b10111010_10111100_01110110_1;
      patterns[47807] = 25'b10111010_10111101_01110111_1;
      patterns[47808] = 25'b10111010_10111110_01111000_1;
      patterns[47809] = 25'b10111010_10111111_01111001_1;
      patterns[47810] = 25'b10111010_11000000_01111010_1;
      patterns[47811] = 25'b10111010_11000001_01111011_1;
      patterns[47812] = 25'b10111010_11000010_01111100_1;
      patterns[47813] = 25'b10111010_11000011_01111101_1;
      patterns[47814] = 25'b10111010_11000100_01111110_1;
      patterns[47815] = 25'b10111010_11000101_01111111_1;
      patterns[47816] = 25'b10111010_11000110_10000000_1;
      patterns[47817] = 25'b10111010_11000111_10000001_1;
      patterns[47818] = 25'b10111010_11001000_10000010_1;
      patterns[47819] = 25'b10111010_11001001_10000011_1;
      patterns[47820] = 25'b10111010_11001010_10000100_1;
      patterns[47821] = 25'b10111010_11001011_10000101_1;
      patterns[47822] = 25'b10111010_11001100_10000110_1;
      patterns[47823] = 25'b10111010_11001101_10000111_1;
      patterns[47824] = 25'b10111010_11001110_10001000_1;
      patterns[47825] = 25'b10111010_11001111_10001001_1;
      patterns[47826] = 25'b10111010_11010000_10001010_1;
      patterns[47827] = 25'b10111010_11010001_10001011_1;
      patterns[47828] = 25'b10111010_11010010_10001100_1;
      patterns[47829] = 25'b10111010_11010011_10001101_1;
      patterns[47830] = 25'b10111010_11010100_10001110_1;
      patterns[47831] = 25'b10111010_11010101_10001111_1;
      patterns[47832] = 25'b10111010_11010110_10010000_1;
      patterns[47833] = 25'b10111010_11010111_10010001_1;
      patterns[47834] = 25'b10111010_11011000_10010010_1;
      patterns[47835] = 25'b10111010_11011001_10010011_1;
      patterns[47836] = 25'b10111010_11011010_10010100_1;
      patterns[47837] = 25'b10111010_11011011_10010101_1;
      patterns[47838] = 25'b10111010_11011100_10010110_1;
      patterns[47839] = 25'b10111010_11011101_10010111_1;
      patterns[47840] = 25'b10111010_11011110_10011000_1;
      patterns[47841] = 25'b10111010_11011111_10011001_1;
      patterns[47842] = 25'b10111010_11100000_10011010_1;
      patterns[47843] = 25'b10111010_11100001_10011011_1;
      patterns[47844] = 25'b10111010_11100010_10011100_1;
      patterns[47845] = 25'b10111010_11100011_10011101_1;
      patterns[47846] = 25'b10111010_11100100_10011110_1;
      patterns[47847] = 25'b10111010_11100101_10011111_1;
      patterns[47848] = 25'b10111010_11100110_10100000_1;
      patterns[47849] = 25'b10111010_11100111_10100001_1;
      patterns[47850] = 25'b10111010_11101000_10100010_1;
      patterns[47851] = 25'b10111010_11101001_10100011_1;
      patterns[47852] = 25'b10111010_11101010_10100100_1;
      patterns[47853] = 25'b10111010_11101011_10100101_1;
      patterns[47854] = 25'b10111010_11101100_10100110_1;
      patterns[47855] = 25'b10111010_11101101_10100111_1;
      patterns[47856] = 25'b10111010_11101110_10101000_1;
      patterns[47857] = 25'b10111010_11101111_10101001_1;
      patterns[47858] = 25'b10111010_11110000_10101010_1;
      patterns[47859] = 25'b10111010_11110001_10101011_1;
      patterns[47860] = 25'b10111010_11110010_10101100_1;
      patterns[47861] = 25'b10111010_11110011_10101101_1;
      patterns[47862] = 25'b10111010_11110100_10101110_1;
      patterns[47863] = 25'b10111010_11110101_10101111_1;
      patterns[47864] = 25'b10111010_11110110_10110000_1;
      patterns[47865] = 25'b10111010_11110111_10110001_1;
      patterns[47866] = 25'b10111010_11111000_10110010_1;
      patterns[47867] = 25'b10111010_11111001_10110011_1;
      patterns[47868] = 25'b10111010_11111010_10110100_1;
      patterns[47869] = 25'b10111010_11111011_10110101_1;
      patterns[47870] = 25'b10111010_11111100_10110110_1;
      patterns[47871] = 25'b10111010_11111101_10110111_1;
      patterns[47872] = 25'b10111010_11111110_10111000_1;
      patterns[47873] = 25'b10111010_11111111_10111001_1;
      patterns[47874] = 25'b10111011_00000000_10111011_0;
      patterns[47875] = 25'b10111011_00000001_10111100_0;
      patterns[47876] = 25'b10111011_00000010_10111101_0;
      patterns[47877] = 25'b10111011_00000011_10111110_0;
      patterns[47878] = 25'b10111011_00000100_10111111_0;
      patterns[47879] = 25'b10111011_00000101_11000000_0;
      patterns[47880] = 25'b10111011_00000110_11000001_0;
      patterns[47881] = 25'b10111011_00000111_11000010_0;
      patterns[47882] = 25'b10111011_00001000_11000011_0;
      patterns[47883] = 25'b10111011_00001001_11000100_0;
      patterns[47884] = 25'b10111011_00001010_11000101_0;
      patterns[47885] = 25'b10111011_00001011_11000110_0;
      patterns[47886] = 25'b10111011_00001100_11000111_0;
      patterns[47887] = 25'b10111011_00001101_11001000_0;
      patterns[47888] = 25'b10111011_00001110_11001001_0;
      patterns[47889] = 25'b10111011_00001111_11001010_0;
      patterns[47890] = 25'b10111011_00010000_11001011_0;
      patterns[47891] = 25'b10111011_00010001_11001100_0;
      patterns[47892] = 25'b10111011_00010010_11001101_0;
      patterns[47893] = 25'b10111011_00010011_11001110_0;
      patterns[47894] = 25'b10111011_00010100_11001111_0;
      patterns[47895] = 25'b10111011_00010101_11010000_0;
      patterns[47896] = 25'b10111011_00010110_11010001_0;
      patterns[47897] = 25'b10111011_00010111_11010010_0;
      patterns[47898] = 25'b10111011_00011000_11010011_0;
      patterns[47899] = 25'b10111011_00011001_11010100_0;
      patterns[47900] = 25'b10111011_00011010_11010101_0;
      patterns[47901] = 25'b10111011_00011011_11010110_0;
      patterns[47902] = 25'b10111011_00011100_11010111_0;
      patterns[47903] = 25'b10111011_00011101_11011000_0;
      patterns[47904] = 25'b10111011_00011110_11011001_0;
      patterns[47905] = 25'b10111011_00011111_11011010_0;
      patterns[47906] = 25'b10111011_00100000_11011011_0;
      patterns[47907] = 25'b10111011_00100001_11011100_0;
      patterns[47908] = 25'b10111011_00100010_11011101_0;
      patterns[47909] = 25'b10111011_00100011_11011110_0;
      patterns[47910] = 25'b10111011_00100100_11011111_0;
      patterns[47911] = 25'b10111011_00100101_11100000_0;
      patterns[47912] = 25'b10111011_00100110_11100001_0;
      patterns[47913] = 25'b10111011_00100111_11100010_0;
      patterns[47914] = 25'b10111011_00101000_11100011_0;
      patterns[47915] = 25'b10111011_00101001_11100100_0;
      patterns[47916] = 25'b10111011_00101010_11100101_0;
      patterns[47917] = 25'b10111011_00101011_11100110_0;
      patterns[47918] = 25'b10111011_00101100_11100111_0;
      patterns[47919] = 25'b10111011_00101101_11101000_0;
      patterns[47920] = 25'b10111011_00101110_11101001_0;
      patterns[47921] = 25'b10111011_00101111_11101010_0;
      patterns[47922] = 25'b10111011_00110000_11101011_0;
      patterns[47923] = 25'b10111011_00110001_11101100_0;
      patterns[47924] = 25'b10111011_00110010_11101101_0;
      patterns[47925] = 25'b10111011_00110011_11101110_0;
      patterns[47926] = 25'b10111011_00110100_11101111_0;
      patterns[47927] = 25'b10111011_00110101_11110000_0;
      patterns[47928] = 25'b10111011_00110110_11110001_0;
      patterns[47929] = 25'b10111011_00110111_11110010_0;
      patterns[47930] = 25'b10111011_00111000_11110011_0;
      patterns[47931] = 25'b10111011_00111001_11110100_0;
      patterns[47932] = 25'b10111011_00111010_11110101_0;
      patterns[47933] = 25'b10111011_00111011_11110110_0;
      patterns[47934] = 25'b10111011_00111100_11110111_0;
      patterns[47935] = 25'b10111011_00111101_11111000_0;
      patterns[47936] = 25'b10111011_00111110_11111001_0;
      patterns[47937] = 25'b10111011_00111111_11111010_0;
      patterns[47938] = 25'b10111011_01000000_11111011_0;
      patterns[47939] = 25'b10111011_01000001_11111100_0;
      patterns[47940] = 25'b10111011_01000010_11111101_0;
      patterns[47941] = 25'b10111011_01000011_11111110_0;
      patterns[47942] = 25'b10111011_01000100_11111111_0;
      patterns[47943] = 25'b10111011_01000101_00000000_1;
      patterns[47944] = 25'b10111011_01000110_00000001_1;
      patterns[47945] = 25'b10111011_01000111_00000010_1;
      patterns[47946] = 25'b10111011_01001000_00000011_1;
      patterns[47947] = 25'b10111011_01001001_00000100_1;
      patterns[47948] = 25'b10111011_01001010_00000101_1;
      patterns[47949] = 25'b10111011_01001011_00000110_1;
      patterns[47950] = 25'b10111011_01001100_00000111_1;
      patterns[47951] = 25'b10111011_01001101_00001000_1;
      patterns[47952] = 25'b10111011_01001110_00001001_1;
      patterns[47953] = 25'b10111011_01001111_00001010_1;
      patterns[47954] = 25'b10111011_01010000_00001011_1;
      patterns[47955] = 25'b10111011_01010001_00001100_1;
      patterns[47956] = 25'b10111011_01010010_00001101_1;
      patterns[47957] = 25'b10111011_01010011_00001110_1;
      patterns[47958] = 25'b10111011_01010100_00001111_1;
      patterns[47959] = 25'b10111011_01010101_00010000_1;
      patterns[47960] = 25'b10111011_01010110_00010001_1;
      patterns[47961] = 25'b10111011_01010111_00010010_1;
      patterns[47962] = 25'b10111011_01011000_00010011_1;
      patterns[47963] = 25'b10111011_01011001_00010100_1;
      patterns[47964] = 25'b10111011_01011010_00010101_1;
      patterns[47965] = 25'b10111011_01011011_00010110_1;
      patterns[47966] = 25'b10111011_01011100_00010111_1;
      patterns[47967] = 25'b10111011_01011101_00011000_1;
      patterns[47968] = 25'b10111011_01011110_00011001_1;
      patterns[47969] = 25'b10111011_01011111_00011010_1;
      patterns[47970] = 25'b10111011_01100000_00011011_1;
      patterns[47971] = 25'b10111011_01100001_00011100_1;
      patterns[47972] = 25'b10111011_01100010_00011101_1;
      patterns[47973] = 25'b10111011_01100011_00011110_1;
      patterns[47974] = 25'b10111011_01100100_00011111_1;
      patterns[47975] = 25'b10111011_01100101_00100000_1;
      patterns[47976] = 25'b10111011_01100110_00100001_1;
      patterns[47977] = 25'b10111011_01100111_00100010_1;
      patterns[47978] = 25'b10111011_01101000_00100011_1;
      patterns[47979] = 25'b10111011_01101001_00100100_1;
      patterns[47980] = 25'b10111011_01101010_00100101_1;
      patterns[47981] = 25'b10111011_01101011_00100110_1;
      patterns[47982] = 25'b10111011_01101100_00100111_1;
      patterns[47983] = 25'b10111011_01101101_00101000_1;
      patterns[47984] = 25'b10111011_01101110_00101001_1;
      patterns[47985] = 25'b10111011_01101111_00101010_1;
      patterns[47986] = 25'b10111011_01110000_00101011_1;
      patterns[47987] = 25'b10111011_01110001_00101100_1;
      patterns[47988] = 25'b10111011_01110010_00101101_1;
      patterns[47989] = 25'b10111011_01110011_00101110_1;
      patterns[47990] = 25'b10111011_01110100_00101111_1;
      patterns[47991] = 25'b10111011_01110101_00110000_1;
      patterns[47992] = 25'b10111011_01110110_00110001_1;
      patterns[47993] = 25'b10111011_01110111_00110010_1;
      patterns[47994] = 25'b10111011_01111000_00110011_1;
      patterns[47995] = 25'b10111011_01111001_00110100_1;
      patterns[47996] = 25'b10111011_01111010_00110101_1;
      patterns[47997] = 25'b10111011_01111011_00110110_1;
      patterns[47998] = 25'b10111011_01111100_00110111_1;
      patterns[47999] = 25'b10111011_01111101_00111000_1;
      patterns[48000] = 25'b10111011_01111110_00111001_1;
      patterns[48001] = 25'b10111011_01111111_00111010_1;
      patterns[48002] = 25'b10111011_10000000_00111011_1;
      patterns[48003] = 25'b10111011_10000001_00111100_1;
      patterns[48004] = 25'b10111011_10000010_00111101_1;
      patterns[48005] = 25'b10111011_10000011_00111110_1;
      patterns[48006] = 25'b10111011_10000100_00111111_1;
      patterns[48007] = 25'b10111011_10000101_01000000_1;
      patterns[48008] = 25'b10111011_10000110_01000001_1;
      patterns[48009] = 25'b10111011_10000111_01000010_1;
      patterns[48010] = 25'b10111011_10001000_01000011_1;
      patterns[48011] = 25'b10111011_10001001_01000100_1;
      patterns[48012] = 25'b10111011_10001010_01000101_1;
      patterns[48013] = 25'b10111011_10001011_01000110_1;
      patterns[48014] = 25'b10111011_10001100_01000111_1;
      patterns[48015] = 25'b10111011_10001101_01001000_1;
      patterns[48016] = 25'b10111011_10001110_01001001_1;
      patterns[48017] = 25'b10111011_10001111_01001010_1;
      patterns[48018] = 25'b10111011_10010000_01001011_1;
      patterns[48019] = 25'b10111011_10010001_01001100_1;
      patterns[48020] = 25'b10111011_10010010_01001101_1;
      patterns[48021] = 25'b10111011_10010011_01001110_1;
      patterns[48022] = 25'b10111011_10010100_01001111_1;
      patterns[48023] = 25'b10111011_10010101_01010000_1;
      patterns[48024] = 25'b10111011_10010110_01010001_1;
      patterns[48025] = 25'b10111011_10010111_01010010_1;
      patterns[48026] = 25'b10111011_10011000_01010011_1;
      patterns[48027] = 25'b10111011_10011001_01010100_1;
      patterns[48028] = 25'b10111011_10011010_01010101_1;
      patterns[48029] = 25'b10111011_10011011_01010110_1;
      patterns[48030] = 25'b10111011_10011100_01010111_1;
      patterns[48031] = 25'b10111011_10011101_01011000_1;
      patterns[48032] = 25'b10111011_10011110_01011001_1;
      patterns[48033] = 25'b10111011_10011111_01011010_1;
      patterns[48034] = 25'b10111011_10100000_01011011_1;
      patterns[48035] = 25'b10111011_10100001_01011100_1;
      patterns[48036] = 25'b10111011_10100010_01011101_1;
      patterns[48037] = 25'b10111011_10100011_01011110_1;
      patterns[48038] = 25'b10111011_10100100_01011111_1;
      patterns[48039] = 25'b10111011_10100101_01100000_1;
      patterns[48040] = 25'b10111011_10100110_01100001_1;
      patterns[48041] = 25'b10111011_10100111_01100010_1;
      patterns[48042] = 25'b10111011_10101000_01100011_1;
      patterns[48043] = 25'b10111011_10101001_01100100_1;
      patterns[48044] = 25'b10111011_10101010_01100101_1;
      patterns[48045] = 25'b10111011_10101011_01100110_1;
      patterns[48046] = 25'b10111011_10101100_01100111_1;
      patterns[48047] = 25'b10111011_10101101_01101000_1;
      patterns[48048] = 25'b10111011_10101110_01101001_1;
      patterns[48049] = 25'b10111011_10101111_01101010_1;
      patterns[48050] = 25'b10111011_10110000_01101011_1;
      patterns[48051] = 25'b10111011_10110001_01101100_1;
      patterns[48052] = 25'b10111011_10110010_01101101_1;
      patterns[48053] = 25'b10111011_10110011_01101110_1;
      patterns[48054] = 25'b10111011_10110100_01101111_1;
      patterns[48055] = 25'b10111011_10110101_01110000_1;
      patterns[48056] = 25'b10111011_10110110_01110001_1;
      patterns[48057] = 25'b10111011_10110111_01110010_1;
      patterns[48058] = 25'b10111011_10111000_01110011_1;
      patterns[48059] = 25'b10111011_10111001_01110100_1;
      patterns[48060] = 25'b10111011_10111010_01110101_1;
      patterns[48061] = 25'b10111011_10111011_01110110_1;
      patterns[48062] = 25'b10111011_10111100_01110111_1;
      patterns[48063] = 25'b10111011_10111101_01111000_1;
      patterns[48064] = 25'b10111011_10111110_01111001_1;
      patterns[48065] = 25'b10111011_10111111_01111010_1;
      patterns[48066] = 25'b10111011_11000000_01111011_1;
      patterns[48067] = 25'b10111011_11000001_01111100_1;
      patterns[48068] = 25'b10111011_11000010_01111101_1;
      patterns[48069] = 25'b10111011_11000011_01111110_1;
      patterns[48070] = 25'b10111011_11000100_01111111_1;
      patterns[48071] = 25'b10111011_11000101_10000000_1;
      patterns[48072] = 25'b10111011_11000110_10000001_1;
      patterns[48073] = 25'b10111011_11000111_10000010_1;
      patterns[48074] = 25'b10111011_11001000_10000011_1;
      patterns[48075] = 25'b10111011_11001001_10000100_1;
      patterns[48076] = 25'b10111011_11001010_10000101_1;
      patterns[48077] = 25'b10111011_11001011_10000110_1;
      patterns[48078] = 25'b10111011_11001100_10000111_1;
      patterns[48079] = 25'b10111011_11001101_10001000_1;
      patterns[48080] = 25'b10111011_11001110_10001001_1;
      patterns[48081] = 25'b10111011_11001111_10001010_1;
      patterns[48082] = 25'b10111011_11010000_10001011_1;
      patterns[48083] = 25'b10111011_11010001_10001100_1;
      patterns[48084] = 25'b10111011_11010010_10001101_1;
      patterns[48085] = 25'b10111011_11010011_10001110_1;
      patterns[48086] = 25'b10111011_11010100_10001111_1;
      patterns[48087] = 25'b10111011_11010101_10010000_1;
      patterns[48088] = 25'b10111011_11010110_10010001_1;
      patterns[48089] = 25'b10111011_11010111_10010010_1;
      patterns[48090] = 25'b10111011_11011000_10010011_1;
      patterns[48091] = 25'b10111011_11011001_10010100_1;
      patterns[48092] = 25'b10111011_11011010_10010101_1;
      patterns[48093] = 25'b10111011_11011011_10010110_1;
      patterns[48094] = 25'b10111011_11011100_10010111_1;
      patterns[48095] = 25'b10111011_11011101_10011000_1;
      patterns[48096] = 25'b10111011_11011110_10011001_1;
      patterns[48097] = 25'b10111011_11011111_10011010_1;
      patterns[48098] = 25'b10111011_11100000_10011011_1;
      patterns[48099] = 25'b10111011_11100001_10011100_1;
      patterns[48100] = 25'b10111011_11100010_10011101_1;
      patterns[48101] = 25'b10111011_11100011_10011110_1;
      patterns[48102] = 25'b10111011_11100100_10011111_1;
      patterns[48103] = 25'b10111011_11100101_10100000_1;
      patterns[48104] = 25'b10111011_11100110_10100001_1;
      patterns[48105] = 25'b10111011_11100111_10100010_1;
      patterns[48106] = 25'b10111011_11101000_10100011_1;
      patterns[48107] = 25'b10111011_11101001_10100100_1;
      patterns[48108] = 25'b10111011_11101010_10100101_1;
      patterns[48109] = 25'b10111011_11101011_10100110_1;
      patterns[48110] = 25'b10111011_11101100_10100111_1;
      patterns[48111] = 25'b10111011_11101101_10101000_1;
      patterns[48112] = 25'b10111011_11101110_10101001_1;
      patterns[48113] = 25'b10111011_11101111_10101010_1;
      patterns[48114] = 25'b10111011_11110000_10101011_1;
      patterns[48115] = 25'b10111011_11110001_10101100_1;
      patterns[48116] = 25'b10111011_11110010_10101101_1;
      patterns[48117] = 25'b10111011_11110011_10101110_1;
      patterns[48118] = 25'b10111011_11110100_10101111_1;
      patterns[48119] = 25'b10111011_11110101_10110000_1;
      patterns[48120] = 25'b10111011_11110110_10110001_1;
      patterns[48121] = 25'b10111011_11110111_10110010_1;
      patterns[48122] = 25'b10111011_11111000_10110011_1;
      patterns[48123] = 25'b10111011_11111001_10110100_1;
      patterns[48124] = 25'b10111011_11111010_10110101_1;
      patterns[48125] = 25'b10111011_11111011_10110110_1;
      patterns[48126] = 25'b10111011_11111100_10110111_1;
      patterns[48127] = 25'b10111011_11111101_10111000_1;
      patterns[48128] = 25'b10111011_11111110_10111001_1;
      patterns[48129] = 25'b10111011_11111111_10111010_1;
      patterns[48130] = 25'b10111100_00000000_10111100_0;
      patterns[48131] = 25'b10111100_00000001_10111101_0;
      patterns[48132] = 25'b10111100_00000010_10111110_0;
      patterns[48133] = 25'b10111100_00000011_10111111_0;
      patterns[48134] = 25'b10111100_00000100_11000000_0;
      patterns[48135] = 25'b10111100_00000101_11000001_0;
      patterns[48136] = 25'b10111100_00000110_11000010_0;
      patterns[48137] = 25'b10111100_00000111_11000011_0;
      patterns[48138] = 25'b10111100_00001000_11000100_0;
      patterns[48139] = 25'b10111100_00001001_11000101_0;
      patterns[48140] = 25'b10111100_00001010_11000110_0;
      patterns[48141] = 25'b10111100_00001011_11000111_0;
      patterns[48142] = 25'b10111100_00001100_11001000_0;
      patterns[48143] = 25'b10111100_00001101_11001001_0;
      patterns[48144] = 25'b10111100_00001110_11001010_0;
      patterns[48145] = 25'b10111100_00001111_11001011_0;
      patterns[48146] = 25'b10111100_00010000_11001100_0;
      patterns[48147] = 25'b10111100_00010001_11001101_0;
      patterns[48148] = 25'b10111100_00010010_11001110_0;
      patterns[48149] = 25'b10111100_00010011_11001111_0;
      patterns[48150] = 25'b10111100_00010100_11010000_0;
      patterns[48151] = 25'b10111100_00010101_11010001_0;
      patterns[48152] = 25'b10111100_00010110_11010010_0;
      patterns[48153] = 25'b10111100_00010111_11010011_0;
      patterns[48154] = 25'b10111100_00011000_11010100_0;
      patterns[48155] = 25'b10111100_00011001_11010101_0;
      patterns[48156] = 25'b10111100_00011010_11010110_0;
      patterns[48157] = 25'b10111100_00011011_11010111_0;
      patterns[48158] = 25'b10111100_00011100_11011000_0;
      patterns[48159] = 25'b10111100_00011101_11011001_0;
      patterns[48160] = 25'b10111100_00011110_11011010_0;
      patterns[48161] = 25'b10111100_00011111_11011011_0;
      patterns[48162] = 25'b10111100_00100000_11011100_0;
      patterns[48163] = 25'b10111100_00100001_11011101_0;
      patterns[48164] = 25'b10111100_00100010_11011110_0;
      patterns[48165] = 25'b10111100_00100011_11011111_0;
      patterns[48166] = 25'b10111100_00100100_11100000_0;
      patterns[48167] = 25'b10111100_00100101_11100001_0;
      patterns[48168] = 25'b10111100_00100110_11100010_0;
      patterns[48169] = 25'b10111100_00100111_11100011_0;
      patterns[48170] = 25'b10111100_00101000_11100100_0;
      patterns[48171] = 25'b10111100_00101001_11100101_0;
      patterns[48172] = 25'b10111100_00101010_11100110_0;
      patterns[48173] = 25'b10111100_00101011_11100111_0;
      patterns[48174] = 25'b10111100_00101100_11101000_0;
      patterns[48175] = 25'b10111100_00101101_11101001_0;
      patterns[48176] = 25'b10111100_00101110_11101010_0;
      patterns[48177] = 25'b10111100_00101111_11101011_0;
      patterns[48178] = 25'b10111100_00110000_11101100_0;
      patterns[48179] = 25'b10111100_00110001_11101101_0;
      patterns[48180] = 25'b10111100_00110010_11101110_0;
      patterns[48181] = 25'b10111100_00110011_11101111_0;
      patterns[48182] = 25'b10111100_00110100_11110000_0;
      patterns[48183] = 25'b10111100_00110101_11110001_0;
      patterns[48184] = 25'b10111100_00110110_11110010_0;
      patterns[48185] = 25'b10111100_00110111_11110011_0;
      patterns[48186] = 25'b10111100_00111000_11110100_0;
      patterns[48187] = 25'b10111100_00111001_11110101_0;
      patterns[48188] = 25'b10111100_00111010_11110110_0;
      patterns[48189] = 25'b10111100_00111011_11110111_0;
      patterns[48190] = 25'b10111100_00111100_11111000_0;
      patterns[48191] = 25'b10111100_00111101_11111001_0;
      patterns[48192] = 25'b10111100_00111110_11111010_0;
      patterns[48193] = 25'b10111100_00111111_11111011_0;
      patterns[48194] = 25'b10111100_01000000_11111100_0;
      patterns[48195] = 25'b10111100_01000001_11111101_0;
      patterns[48196] = 25'b10111100_01000010_11111110_0;
      patterns[48197] = 25'b10111100_01000011_11111111_0;
      patterns[48198] = 25'b10111100_01000100_00000000_1;
      patterns[48199] = 25'b10111100_01000101_00000001_1;
      patterns[48200] = 25'b10111100_01000110_00000010_1;
      patterns[48201] = 25'b10111100_01000111_00000011_1;
      patterns[48202] = 25'b10111100_01001000_00000100_1;
      patterns[48203] = 25'b10111100_01001001_00000101_1;
      patterns[48204] = 25'b10111100_01001010_00000110_1;
      patterns[48205] = 25'b10111100_01001011_00000111_1;
      patterns[48206] = 25'b10111100_01001100_00001000_1;
      patterns[48207] = 25'b10111100_01001101_00001001_1;
      patterns[48208] = 25'b10111100_01001110_00001010_1;
      patterns[48209] = 25'b10111100_01001111_00001011_1;
      patterns[48210] = 25'b10111100_01010000_00001100_1;
      patterns[48211] = 25'b10111100_01010001_00001101_1;
      patterns[48212] = 25'b10111100_01010010_00001110_1;
      patterns[48213] = 25'b10111100_01010011_00001111_1;
      patterns[48214] = 25'b10111100_01010100_00010000_1;
      patterns[48215] = 25'b10111100_01010101_00010001_1;
      patterns[48216] = 25'b10111100_01010110_00010010_1;
      patterns[48217] = 25'b10111100_01010111_00010011_1;
      patterns[48218] = 25'b10111100_01011000_00010100_1;
      patterns[48219] = 25'b10111100_01011001_00010101_1;
      patterns[48220] = 25'b10111100_01011010_00010110_1;
      patterns[48221] = 25'b10111100_01011011_00010111_1;
      patterns[48222] = 25'b10111100_01011100_00011000_1;
      patterns[48223] = 25'b10111100_01011101_00011001_1;
      patterns[48224] = 25'b10111100_01011110_00011010_1;
      patterns[48225] = 25'b10111100_01011111_00011011_1;
      patterns[48226] = 25'b10111100_01100000_00011100_1;
      patterns[48227] = 25'b10111100_01100001_00011101_1;
      patterns[48228] = 25'b10111100_01100010_00011110_1;
      patterns[48229] = 25'b10111100_01100011_00011111_1;
      patterns[48230] = 25'b10111100_01100100_00100000_1;
      patterns[48231] = 25'b10111100_01100101_00100001_1;
      patterns[48232] = 25'b10111100_01100110_00100010_1;
      patterns[48233] = 25'b10111100_01100111_00100011_1;
      patterns[48234] = 25'b10111100_01101000_00100100_1;
      patterns[48235] = 25'b10111100_01101001_00100101_1;
      patterns[48236] = 25'b10111100_01101010_00100110_1;
      patterns[48237] = 25'b10111100_01101011_00100111_1;
      patterns[48238] = 25'b10111100_01101100_00101000_1;
      patterns[48239] = 25'b10111100_01101101_00101001_1;
      patterns[48240] = 25'b10111100_01101110_00101010_1;
      patterns[48241] = 25'b10111100_01101111_00101011_1;
      patterns[48242] = 25'b10111100_01110000_00101100_1;
      patterns[48243] = 25'b10111100_01110001_00101101_1;
      patterns[48244] = 25'b10111100_01110010_00101110_1;
      patterns[48245] = 25'b10111100_01110011_00101111_1;
      patterns[48246] = 25'b10111100_01110100_00110000_1;
      patterns[48247] = 25'b10111100_01110101_00110001_1;
      patterns[48248] = 25'b10111100_01110110_00110010_1;
      patterns[48249] = 25'b10111100_01110111_00110011_1;
      patterns[48250] = 25'b10111100_01111000_00110100_1;
      patterns[48251] = 25'b10111100_01111001_00110101_1;
      patterns[48252] = 25'b10111100_01111010_00110110_1;
      patterns[48253] = 25'b10111100_01111011_00110111_1;
      patterns[48254] = 25'b10111100_01111100_00111000_1;
      patterns[48255] = 25'b10111100_01111101_00111001_1;
      patterns[48256] = 25'b10111100_01111110_00111010_1;
      patterns[48257] = 25'b10111100_01111111_00111011_1;
      patterns[48258] = 25'b10111100_10000000_00111100_1;
      patterns[48259] = 25'b10111100_10000001_00111101_1;
      patterns[48260] = 25'b10111100_10000010_00111110_1;
      patterns[48261] = 25'b10111100_10000011_00111111_1;
      patterns[48262] = 25'b10111100_10000100_01000000_1;
      patterns[48263] = 25'b10111100_10000101_01000001_1;
      patterns[48264] = 25'b10111100_10000110_01000010_1;
      patterns[48265] = 25'b10111100_10000111_01000011_1;
      patterns[48266] = 25'b10111100_10001000_01000100_1;
      patterns[48267] = 25'b10111100_10001001_01000101_1;
      patterns[48268] = 25'b10111100_10001010_01000110_1;
      patterns[48269] = 25'b10111100_10001011_01000111_1;
      patterns[48270] = 25'b10111100_10001100_01001000_1;
      patterns[48271] = 25'b10111100_10001101_01001001_1;
      patterns[48272] = 25'b10111100_10001110_01001010_1;
      patterns[48273] = 25'b10111100_10001111_01001011_1;
      patterns[48274] = 25'b10111100_10010000_01001100_1;
      patterns[48275] = 25'b10111100_10010001_01001101_1;
      patterns[48276] = 25'b10111100_10010010_01001110_1;
      patterns[48277] = 25'b10111100_10010011_01001111_1;
      patterns[48278] = 25'b10111100_10010100_01010000_1;
      patterns[48279] = 25'b10111100_10010101_01010001_1;
      patterns[48280] = 25'b10111100_10010110_01010010_1;
      patterns[48281] = 25'b10111100_10010111_01010011_1;
      patterns[48282] = 25'b10111100_10011000_01010100_1;
      patterns[48283] = 25'b10111100_10011001_01010101_1;
      patterns[48284] = 25'b10111100_10011010_01010110_1;
      patterns[48285] = 25'b10111100_10011011_01010111_1;
      patterns[48286] = 25'b10111100_10011100_01011000_1;
      patterns[48287] = 25'b10111100_10011101_01011001_1;
      patterns[48288] = 25'b10111100_10011110_01011010_1;
      patterns[48289] = 25'b10111100_10011111_01011011_1;
      patterns[48290] = 25'b10111100_10100000_01011100_1;
      patterns[48291] = 25'b10111100_10100001_01011101_1;
      patterns[48292] = 25'b10111100_10100010_01011110_1;
      patterns[48293] = 25'b10111100_10100011_01011111_1;
      patterns[48294] = 25'b10111100_10100100_01100000_1;
      patterns[48295] = 25'b10111100_10100101_01100001_1;
      patterns[48296] = 25'b10111100_10100110_01100010_1;
      patterns[48297] = 25'b10111100_10100111_01100011_1;
      patterns[48298] = 25'b10111100_10101000_01100100_1;
      patterns[48299] = 25'b10111100_10101001_01100101_1;
      patterns[48300] = 25'b10111100_10101010_01100110_1;
      patterns[48301] = 25'b10111100_10101011_01100111_1;
      patterns[48302] = 25'b10111100_10101100_01101000_1;
      patterns[48303] = 25'b10111100_10101101_01101001_1;
      patterns[48304] = 25'b10111100_10101110_01101010_1;
      patterns[48305] = 25'b10111100_10101111_01101011_1;
      patterns[48306] = 25'b10111100_10110000_01101100_1;
      patterns[48307] = 25'b10111100_10110001_01101101_1;
      patterns[48308] = 25'b10111100_10110010_01101110_1;
      patterns[48309] = 25'b10111100_10110011_01101111_1;
      patterns[48310] = 25'b10111100_10110100_01110000_1;
      patterns[48311] = 25'b10111100_10110101_01110001_1;
      patterns[48312] = 25'b10111100_10110110_01110010_1;
      patterns[48313] = 25'b10111100_10110111_01110011_1;
      patterns[48314] = 25'b10111100_10111000_01110100_1;
      patterns[48315] = 25'b10111100_10111001_01110101_1;
      patterns[48316] = 25'b10111100_10111010_01110110_1;
      patterns[48317] = 25'b10111100_10111011_01110111_1;
      patterns[48318] = 25'b10111100_10111100_01111000_1;
      patterns[48319] = 25'b10111100_10111101_01111001_1;
      patterns[48320] = 25'b10111100_10111110_01111010_1;
      patterns[48321] = 25'b10111100_10111111_01111011_1;
      patterns[48322] = 25'b10111100_11000000_01111100_1;
      patterns[48323] = 25'b10111100_11000001_01111101_1;
      patterns[48324] = 25'b10111100_11000010_01111110_1;
      patterns[48325] = 25'b10111100_11000011_01111111_1;
      patterns[48326] = 25'b10111100_11000100_10000000_1;
      patterns[48327] = 25'b10111100_11000101_10000001_1;
      patterns[48328] = 25'b10111100_11000110_10000010_1;
      patterns[48329] = 25'b10111100_11000111_10000011_1;
      patterns[48330] = 25'b10111100_11001000_10000100_1;
      patterns[48331] = 25'b10111100_11001001_10000101_1;
      patterns[48332] = 25'b10111100_11001010_10000110_1;
      patterns[48333] = 25'b10111100_11001011_10000111_1;
      patterns[48334] = 25'b10111100_11001100_10001000_1;
      patterns[48335] = 25'b10111100_11001101_10001001_1;
      patterns[48336] = 25'b10111100_11001110_10001010_1;
      patterns[48337] = 25'b10111100_11001111_10001011_1;
      patterns[48338] = 25'b10111100_11010000_10001100_1;
      patterns[48339] = 25'b10111100_11010001_10001101_1;
      patterns[48340] = 25'b10111100_11010010_10001110_1;
      patterns[48341] = 25'b10111100_11010011_10001111_1;
      patterns[48342] = 25'b10111100_11010100_10010000_1;
      patterns[48343] = 25'b10111100_11010101_10010001_1;
      patterns[48344] = 25'b10111100_11010110_10010010_1;
      patterns[48345] = 25'b10111100_11010111_10010011_1;
      patterns[48346] = 25'b10111100_11011000_10010100_1;
      patterns[48347] = 25'b10111100_11011001_10010101_1;
      patterns[48348] = 25'b10111100_11011010_10010110_1;
      patterns[48349] = 25'b10111100_11011011_10010111_1;
      patterns[48350] = 25'b10111100_11011100_10011000_1;
      patterns[48351] = 25'b10111100_11011101_10011001_1;
      patterns[48352] = 25'b10111100_11011110_10011010_1;
      patterns[48353] = 25'b10111100_11011111_10011011_1;
      patterns[48354] = 25'b10111100_11100000_10011100_1;
      patterns[48355] = 25'b10111100_11100001_10011101_1;
      patterns[48356] = 25'b10111100_11100010_10011110_1;
      patterns[48357] = 25'b10111100_11100011_10011111_1;
      patterns[48358] = 25'b10111100_11100100_10100000_1;
      patterns[48359] = 25'b10111100_11100101_10100001_1;
      patterns[48360] = 25'b10111100_11100110_10100010_1;
      patterns[48361] = 25'b10111100_11100111_10100011_1;
      patterns[48362] = 25'b10111100_11101000_10100100_1;
      patterns[48363] = 25'b10111100_11101001_10100101_1;
      patterns[48364] = 25'b10111100_11101010_10100110_1;
      patterns[48365] = 25'b10111100_11101011_10100111_1;
      patterns[48366] = 25'b10111100_11101100_10101000_1;
      patterns[48367] = 25'b10111100_11101101_10101001_1;
      patterns[48368] = 25'b10111100_11101110_10101010_1;
      patterns[48369] = 25'b10111100_11101111_10101011_1;
      patterns[48370] = 25'b10111100_11110000_10101100_1;
      patterns[48371] = 25'b10111100_11110001_10101101_1;
      patterns[48372] = 25'b10111100_11110010_10101110_1;
      patterns[48373] = 25'b10111100_11110011_10101111_1;
      patterns[48374] = 25'b10111100_11110100_10110000_1;
      patterns[48375] = 25'b10111100_11110101_10110001_1;
      patterns[48376] = 25'b10111100_11110110_10110010_1;
      patterns[48377] = 25'b10111100_11110111_10110011_1;
      patterns[48378] = 25'b10111100_11111000_10110100_1;
      patterns[48379] = 25'b10111100_11111001_10110101_1;
      patterns[48380] = 25'b10111100_11111010_10110110_1;
      patterns[48381] = 25'b10111100_11111011_10110111_1;
      patterns[48382] = 25'b10111100_11111100_10111000_1;
      patterns[48383] = 25'b10111100_11111101_10111001_1;
      patterns[48384] = 25'b10111100_11111110_10111010_1;
      patterns[48385] = 25'b10111100_11111111_10111011_1;
      patterns[48386] = 25'b10111101_00000000_10111101_0;
      patterns[48387] = 25'b10111101_00000001_10111110_0;
      patterns[48388] = 25'b10111101_00000010_10111111_0;
      patterns[48389] = 25'b10111101_00000011_11000000_0;
      patterns[48390] = 25'b10111101_00000100_11000001_0;
      patterns[48391] = 25'b10111101_00000101_11000010_0;
      patterns[48392] = 25'b10111101_00000110_11000011_0;
      patterns[48393] = 25'b10111101_00000111_11000100_0;
      patterns[48394] = 25'b10111101_00001000_11000101_0;
      patterns[48395] = 25'b10111101_00001001_11000110_0;
      patterns[48396] = 25'b10111101_00001010_11000111_0;
      patterns[48397] = 25'b10111101_00001011_11001000_0;
      patterns[48398] = 25'b10111101_00001100_11001001_0;
      patterns[48399] = 25'b10111101_00001101_11001010_0;
      patterns[48400] = 25'b10111101_00001110_11001011_0;
      patterns[48401] = 25'b10111101_00001111_11001100_0;
      patterns[48402] = 25'b10111101_00010000_11001101_0;
      patterns[48403] = 25'b10111101_00010001_11001110_0;
      patterns[48404] = 25'b10111101_00010010_11001111_0;
      patterns[48405] = 25'b10111101_00010011_11010000_0;
      patterns[48406] = 25'b10111101_00010100_11010001_0;
      patterns[48407] = 25'b10111101_00010101_11010010_0;
      patterns[48408] = 25'b10111101_00010110_11010011_0;
      patterns[48409] = 25'b10111101_00010111_11010100_0;
      patterns[48410] = 25'b10111101_00011000_11010101_0;
      patterns[48411] = 25'b10111101_00011001_11010110_0;
      patterns[48412] = 25'b10111101_00011010_11010111_0;
      patterns[48413] = 25'b10111101_00011011_11011000_0;
      patterns[48414] = 25'b10111101_00011100_11011001_0;
      patterns[48415] = 25'b10111101_00011101_11011010_0;
      patterns[48416] = 25'b10111101_00011110_11011011_0;
      patterns[48417] = 25'b10111101_00011111_11011100_0;
      patterns[48418] = 25'b10111101_00100000_11011101_0;
      patterns[48419] = 25'b10111101_00100001_11011110_0;
      patterns[48420] = 25'b10111101_00100010_11011111_0;
      patterns[48421] = 25'b10111101_00100011_11100000_0;
      patterns[48422] = 25'b10111101_00100100_11100001_0;
      patterns[48423] = 25'b10111101_00100101_11100010_0;
      patterns[48424] = 25'b10111101_00100110_11100011_0;
      patterns[48425] = 25'b10111101_00100111_11100100_0;
      patterns[48426] = 25'b10111101_00101000_11100101_0;
      patterns[48427] = 25'b10111101_00101001_11100110_0;
      patterns[48428] = 25'b10111101_00101010_11100111_0;
      patterns[48429] = 25'b10111101_00101011_11101000_0;
      patterns[48430] = 25'b10111101_00101100_11101001_0;
      patterns[48431] = 25'b10111101_00101101_11101010_0;
      patterns[48432] = 25'b10111101_00101110_11101011_0;
      patterns[48433] = 25'b10111101_00101111_11101100_0;
      patterns[48434] = 25'b10111101_00110000_11101101_0;
      patterns[48435] = 25'b10111101_00110001_11101110_0;
      patterns[48436] = 25'b10111101_00110010_11101111_0;
      patterns[48437] = 25'b10111101_00110011_11110000_0;
      patterns[48438] = 25'b10111101_00110100_11110001_0;
      patterns[48439] = 25'b10111101_00110101_11110010_0;
      patterns[48440] = 25'b10111101_00110110_11110011_0;
      patterns[48441] = 25'b10111101_00110111_11110100_0;
      patterns[48442] = 25'b10111101_00111000_11110101_0;
      patterns[48443] = 25'b10111101_00111001_11110110_0;
      patterns[48444] = 25'b10111101_00111010_11110111_0;
      patterns[48445] = 25'b10111101_00111011_11111000_0;
      patterns[48446] = 25'b10111101_00111100_11111001_0;
      patterns[48447] = 25'b10111101_00111101_11111010_0;
      patterns[48448] = 25'b10111101_00111110_11111011_0;
      patterns[48449] = 25'b10111101_00111111_11111100_0;
      patterns[48450] = 25'b10111101_01000000_11111101_0;
      patterns[48451] = 25'b10111101_01000001_11111110_0;
      patterns[48452] = 25'b10111101_01000010_11111111_0;
      patterns[48453] = 25'b10111101_01000011_00000000_1;
      patterns[48454] = 25'b10111101_01000100_00000001_1;
      patterns[48455] = 25'b10111101_01000101_00000010_1;
      patterns[48456] = 25'b10111101_01000110_00000011_1;
      patterns[48457] = 25'b10111101_01000111_00000100_1;
      patterns[48458] = 25'b10111101_01001000_00000101_1;
      patterns[48459] = 25'b10111101_01001001_00000110_1;
      patterns[48460] = 25'b10111101_01001010_00000111_1;
      patterns[48461] = 25'b10111101_01001011_00001000_1;
      patterns[48462] = 25'b10111101_01001100_00001001_1;
      patterns[48463] = 25'b10111101_01001101_00001010_1;
      patterns[48464] = 25'b10111101_01001110_00001011_1;
      patterns[48465] = 25'b10111101_01001111_00001100_1;
      patterns[48466] = 25'b10111101_01010000_00001101_1;
      patterns[48467] = 25'b10111101_01010001_00001110_1;
      patterns[48468] = 25'b10111101_01010010_00001111_1;
      patterns[48469] = 25'b10111101_01010011_00010000_1;
      patterns[48470] = 25'b10111101_01010100_00010001_1;
      patterns[48471] = 25'b10111101_01010101_00010010_1;
      patterns[48472] = 25'b10111101_01010110_00010011_1;
      patterns[48473] = 25'b10111101_01010111_00010100_1;
      patterns[48474] = 25'b10111101_01011000_00010101_1;
      patterns[48475] = 25'b10111101_01011001_00010110_1;
      patterns[48476] = 25'b10111101_01011010_00010111_1;
      patterns[48477] = 25'b10111101_01011011_00011000_1;
      patterns[48478] = 25'b10111101_01011100_00011001_1;
      patterns[48479] = 25'b10111101_01011101_00011010_1;
      patterns[48480] = 25'b10111101_01011110_00011011_1;
      patterns[48481] = 25'b10111101_01011111_00011100_1;
      patterns[48482] = 25'b10111101_01100000_00011101_1;
      patterns[48483] = 25'b10111101_01100001_00011110_1;
      patterns[48484] = 25'b10111101_01100010_00011111_1;
      patterns[48485] = 25'b10111101_01100011_00100000_1;
      patterns[48486] = 25'b10111101_01100100_00100001_1;
      patterns[48487] = 25'b10111101_01100101_00100010_1;
      patterns[48488] = 25'b10111101_01100110_00100011_1;
      patterns[48489] = 25'b10111101_01100111_00100100_1;
      patterns[48490] = 25'b10111101_01101000_00100101_1;
      patterns[48491] = 25'b10111101_01101001_00100110_1;
      patterns[48492] = 25'b10111101_01101010_00100111_1;
      patterns[48493] = 25'b10111101_01101011_00101000_1;
      patterns[48494] = 25'b10111101_01101100_00101001_1;
      patterns[48495] = 25'b10111101_01101101_00101010_1;
      patterns[48496] = 25'b10111101_01101110_00101011_1;
      patterns[48497] = 25'b10111101_01101111_00101100_1;
      patterns[48498] = 25'b10111101_01110000_00101101_1;
      patterns[48499] = 25'b10111101_01110001_00101110_1;
      patterns[48500] = 25'b10111101_01110010_00101111_1;
      patterns[48501] = 25'b10111101_01110011_00110000_1;
      patterns[48502] = 25'b10111101_01110100_00110001_1;
      patterns[48503] = 25'b10111101_01110101_00110010_1;
      patterns[48504] = 25'b10111101_01110110_00110011_1;
      patterns[48505] = 25'b10111101_01110111_00110100_1;
      patterns[48506] = 25'b10111101_01111000_00110101_1;
      patterns[48507] = 25'b10111101_01111001_00110110_1;
      patterns[48508] = 25'b10111101_01111010_00110111_1;
      patterns[48509] = 25'b10111101_01111011_00111000_1;
      patterns[48510] = 25'b10111101_01111100_00111001_1;
      patterns[48511] = 25'b10111101_01111101_00111010_1;
      patterns[48512] = 25'b10111101_01111110_00111011_1;
      patterns[48513] = 25'b10111101_01111111_00111100_1;
      patterns[48514] = 25'b10111101_10000000_00111101_1;
      patterns[48515] = 25'b10111101_10000001_00111110_1;
      patterns[48516] = 25'b10111101_10000010_00111111_1;
      patterns[48517] = 25'b10111101_10000011_01000000_1;
      patterns[48518] = 25'b10111101_10000100_01000001_1;
      patterns[48519] = 25'b10111101_10000101_01000010_1;
      patterns[48520] = 25'b10111101_10000110_01000011_1;
      patterns[48521] = 25'b10111101_10000111_01000100_1;
      patterns[48522] = 25'b10111101_10001000_01000101_1;
      patterns[48523] = 25'b10111101_10001001_01000110_1;
      patterns[48524] = 25'b10111101_10001010_01000111_1;
      patterns[48525] = 25'b10111101_10001011_01001000_1;
      patterns[48526] = 25'b10111101_10001100_01001001_1;
      patterns[48527] = 25'b10111101_10001101_01001010_1;
      patterns[48528] = 25'b10111101_10001110_01001011_1;
      patterns[48529] = 25'b10111101_10001111_01001100_1;
      patterns[48530] = 25'b10111101_10010000_01001101_1;
      patterns[48531] = 25'b10111101_10010001_01001110_1;
      patterns[48532] = 25'b10111101_10010010_01001111_1;
      patterns[48533] = 25'b10111101_10010011_01010000_1;
      patterns[48534] = 25'b10111101_10010100_01010001_1;
      patterns[48535] = 25'b10111101_10010101_01010010_1;
      patterns[48536] = 25'b10111101_10010110_01010011_1;
      patterns[48537] = 25'b10111101_10010111_01010100_1;
      patterns[48538] = 25'b10111101_10011000_01010101_1;
      patterns[48539] = 25'b10111101_10011001_01010110_1;
      patterns[48540] = 25'b10111101_10011010_01010111_1;
      patterns[48541] = 25'b10111101_10011011_01011000_1;
      patterns[48542] = 25'b10111101_10011100_01011001_1;
      patterns[48543] = 25'b10111101_10011101_01011010_1;
      patterns[48544] = 25'b10111101_10011110_01011011_1;
      patterns[48545] = 25'b10111101_10011111_01011100_1;
      patterns[48546] = 25'b10111101_10100000_01011101_1;
      patterns[48547] = 25'b10111101_10100001_01011110_1;
      patterns[48548] = 25'b10111101_10100010_01011111_1;
      patterns[48549] = 25'b10111101_10100011_01100000_1;
      patterns[48550] = 25'b10111101_10100100_01100001_1;
      patterns[48551] = 25'b10111101_10100101_01100010_1;
      patterns[48552] = 25'b10111101_10100110_01100011_1;
      patterns[48553] = 25'b10111101_10100111_01100100_1;
      patterns[48554] = 25'b10111101_10101000_01100101_1;
      patterns[48555] = 25'b10111101_10101001_01100110_1;
      patterns[48556] = 25'b10111101_10101010_01100111_1;
      patterns[48557] = 25'b10111101_10101011_01101000_1;
      patterns[48558] = 25'b10111101_10101100_01101001_1;
      patterns[48559] = 25'b10111101_10101101_01101010_1;
      patterns[48560] = 25'b10111101_10101110_01101011_1;
      patterns[48561] = 25'b10111101_10101111_01101100_1;
      patterns[48562] = 25'b10111101_10110000_01101101_1;
      patterns[48563] = 25'b10111101_10110001_01101110_1;
      patterns[48564] = 25'b10111101_10110010_01101111_1;
      patterns[48565] = 25'b10111101_10110011_01110000_1;
      patterns[48566] = 25'b10111101_10110100_01110001_1;
      patterns[48567] = 25'b10111101_10110101_01110010_1;
      patterns[48568] = 25'b10111101_10110110_01110011_1;
      patterns[48569] = 25'b10111101_10110111_01110100_1;
      patterns[48570] = 25'b10111101_10111000_01110101_1;
      patterns[48571] = 25'b10111101_10111001_01110110_1;
      patterns[48572] = 25'b10111101_10111010_01110111_1;
      patterns[48573] = 25'b10111101_10111011_01111000_1;
      patterns[48574] = 25'b10111101_10111100_01111001_1;
      patterns[48575] = 25'b10111101_10111101_01111010_1;
      patterns[48576] = 25'b10111101_10111110_01111011_1;
      patterns[48577] = 25'b10111101_10111111_01111100_1;
      patterns[48578] = 25'b10111101_11000000_01111101_1;
      patterns[48579] = 25'b10111101_11000001_01111110_1;
      patterns[48580] = 25'b10111101_11000010_01111111_1;
      patterns[48581] = 25'b10111101_11000011_10000000_1;
      patterns[48582] = 25'b10111101_11000100_10000001_1;
      patterns[48583] = 25'b10111101_11000101_10000010_1;
      patterns[48584] = 25'b10111101_11000110_10000011_1;
      patterns[48585] = 25'b10111101_11000111_10000100_1;
      patterns[48586] = 25'b10111101_11001000_10000101_1;
      patterns[48587] = 25'b10111101_11001001_10000110_1;
      patterns[48588] = 25'b10111101_11001010_10000111_1;
      patterns[48589] = 25'b10111101_11001011_10001000_1;
      patterns[48590] = 25'b10111101_11001100_10001001_1;
      patterns[48591] = 25'b10111101_11001101_10001010_1;
      patterns[48592] = 25'b10111101_11001110_10001011_1;
      patterns[48593] = 25'b10111101_11001111_10001100_1;
      patterns[48594] = 25'b10111101_11010000_10001101_1;
      patterns[48595] = 25'b10111101_11010001_10001110_1;
      patterns[48596] = 25'b10111101_11010010_10001111_1;
      patterns[48597] = 25'b10111101_11010011_10010000_1;
      patterns[48598] = 25'b10111101_11010100_10010001_1;
      patterns[48599] = 25'b10111101_11010101_10010010_1;
      patterns[48600] = 25'b10111101_11010110_10010011_1;
      patterns[48601] = 25'b10111101_11010111_10010100_1;
      patterns[48602] = 25'b10111101_11011000_10010101_1;
      patterns[48603] = 25'b10111101_11011001_10010110_1;
      patterns[48604] = 25'b10111101_11011010_10010111_1;
      patterns[48605] = 25'b10111101_11011011_10011000_1;
      patterns[48606] = 25'b10111101_11011100_10011001_1;
      patterns[48607] = 25'b10111101_11011101_10011010_1;
      patterns[48608] = 25'b10111101_11011110_10011011_1;
      patterns[48609] = 25'b10111101_11011111_10011100_1;
      patterns[48610] = 25'b10111101_11100000_10011101_1;
      patterns[48611] = 25'b10111101_11100001_10011110_1;
      patterns[48612] = 25'b10111101_11100010_10011111_1;
      patterns[48613] = 25'b10111101_11100011_10100000_1;
      patterns[48614] = 25'b10111101_11100100_10100001_1;
      patterns[48615] = 25'b10111101_11100101_10100010_1;
      patterns[48616] = 25'b10111101_11100110_10100011_1;
      patterns[48617] = 25'b10111101_11100111_10100100_1;
      patterns[48618] = 25'b10111101_11101000_10100101_1;
      patterns[48619] = 25'b10111101_11101001_10100110_1;
      patterns[48620] = 25'b10111101_11101010_10100111_1;
      patterns[48621] = 25'b10111101_11101011_10101000_1;
      patterns[48622] = 25'b10111101_11101100_10101001_1;
      patterns[48623] = 25'b10111101_11101101_10101010_1;
      patterns[48624] = 25'b10111101_11101110_10101011_1;
      patterns[48625] = 25'b10111101_11101111_10101100_1;
      patterns[48626] = 25'b10111101_11110000_10101101_1;
      patterns[48627] = 25'b10111101_11110001_10101110_1;
      patterns[48628] = 25'b10111101_11110010_10101111_1;
      patterns[48629] = 25'b10111101_11110011_10110000_1;
      patterns[48630] = 25'b10111101_11110100_10110001_1;
      patterns[48631] = 25'b10111101_11110101_10110010_1;
      patterns[48632] = 25'b10111101_11110110_10110011_1;
      patterns[48633] = 25'b10111101_11110111_10110100_1;
      patterns[48634] = 25'b10111101_11111000_10110101_1;
      patterns[48635] = 25'b10111101_11111001_10110110_1;
      patterns[48636] = 25'b10111101_11111010_10110111_1;
      patterns[48637] = 25'b10111101_11111011_10111000_1;
      patterns[48638] = 25'b10111101_11111100_10111001_1;
      patterns[48639] = 25'b10111101_11111101_10111010_1;
      patterns[48640] = 25'b10111101_11111110_10111011_1;
      patterns[48641] = 25'b10111101_11111111_10111100_1;
      patterns[48642] = 25'b10111110_00000000_10111110_0;
      patterns[48643] = 25'b10111110_00000001_10111111_0;
      patterns[48644] = 25'b10111110_00000010_11000000_0;
      patterns[48645] = 25'b10111110_00000011_11000001_0;
      patterns[48646] = 25'b10111110_00000100_11000010_0;
      patterns[48647] = 25'b10111110_00000101_11000011_0;
      patterns[48648] = 25'b10111110_00000110_11000100_0;
      patterns[48649] = 25'b10111110_00000111_11000101_0;
      patterns[48650] = 25'b10111110_00001000_11000110_0;
      patterns[48651] = 25'b10111110_00001001_11000111_0;
      patterns[48652] = 25'b10111110_00001010_11001000_0;
      patterns[48653] = 25'b10111110_00001011_11001001_0;
      patterns[48654] = 25'b10111110_00001100_11001010_0;
      patterns[48655] = 25'b10111110_00001101_11001011_0;
      patterns[48656] = 25'b10111110_00001110_11001100_0;
      patterns[48657] = 25'b10111110_00001111_11001101_0;
      patterns[48658] = 25'b10111110_00010000_11001110_0;
      patterns[48659] = 25'b10111110_00010001_11001111_0;
      patterns[48660] = 25'b10111110_00010010_11010000_0;
      patterns[48661] = 25'b10111110_00010011_11010001_0;
      patterns[48662] = 25'b10111110_00010100_11010010_0;
      patterns[48663] = 25'b10111110_00010101_11010011_0;
      patterns[48664] = 25'b10111110_00010110_11010100_0;
      patterns[48665] = 25'b10111110_00010111_11010101_0;
      patterns[48666] = 25'b10111110_00011000_11010110_0;
      patterns[48667] = 25'b10111110_00011001_11010111_0;
      patterns[48668] = 25'b10111110_00011010_11011000_0;
      patterns[48669] = 25'b10111110_00011011_11011001_0;
      patterns[48670] = 25'b10111110_00011100_11011010_0;
      patterns[48671] = 25'b10111110_00011101_11011011_0;
      patterns[48672] = 25'b10111110_00011110_11011100_0;
      patterns[48673] = 25'b10111110_00011111_11011101_0;
      patterns[48674] = 25'b10111110_00100000_11011110_0;
      patterns[48675] = 25'b10111110_00100001_11011111_0;
      patterns[48676] = 25'b10111110_00100010_11100000_0;
      patterns[48677] = 25'b10111110_00100011_11100001_0;
      patterns[48678] = 25'b10111110_00100100_11100010_0;
      patterns[48679] = 25'b10111110_00100101_11100011_0;
      patterns[48680] = 25'b10111110_00100110_11100100_0;
      patterns[48681] = 25'b10111110_00100111_11100101_0;
      patterns[48682] = 25'b10111110_00101000_11100110_0;
      patterns[48683] = 25'b10111110_00101001_11100111_0;
      patterns[48684] = 25'b10111110_00101010_11101000_0;
      patterns[48685] = 25'b10111110_00101011_11101001_0;
      patterns[48686] = 25'b10111110_00101100_11101010_0;
      patterns[48687] = 25'b10111110_00101101_11101011_0;
      patterns[48688] = 25'b10111110_00101110_11101100_0;
      patterns[48689] = 25'b10111110_00101111_11101101_0;
      patterns[48690] = 25'b10111110_00110000_11101110_0;
      patterns[48691] = 25'b10111110_00110001_11101111_0;
      patterns[48692] = 25'b10111110_00110010_11110000_0;
      patterns[48693] = 25'b10111110_00110011_11110001_0;
      patterns[48694] = 25'b10111110_00110100_11110010_0;
      patterns[48695] = 25'b10111110_00110101_11110011_0;
      patterns[48696] = 25'b10111110_00110110_11110100_0;
      patterns[48697] = 25'b10111110_00110111_11110101_0;
      patterns[48698] = 25'b10111110_00111000_11110110_0;
      patterns[48699] = 25'b10111110_00111001_11110111_0;
      patterns[48700] = 25'b10111110_00111010_11111000_0;
      patterns[48701] = 25'b10111110_00111011_11111001_0;
      patterns[48702] = 25'b10111110_00111100_11111010_0;
      patterns[48703] = 25'b10111110_00111101_11111011_0;
      patterns[48704] = 25'b10111110_00111110_11111100_0;
      patterns[48705] = 25'b10111110_00111111_11111101_0;
      patterns[48706] = 25'b10111110_01000000_11111110_0;
      patterns[48707] = 25'b10111110_01000001_11111111_0;
      patterns[48708] = 25'b10111110_01000010_00000000_1;
      patterns[48709] = 25'b10111110_01000011_00000001_1;
      patterns[48710] = 25'b10111110_01000100_00000010_1;
      patterns[48711] = 25'b10111110_01000101_00000011_1;
      patterns[48712] = 25'b10111110_01000110_00000100_1;
      patterns[48713] = 25'b10111110_01000111_00000101_1;
      patterns[48714] = 25'b10111110_01001000_00000110_1;
      patterns[48715] = 25'b10111110_01001001_00000111_1;
      patterns[48716] = 25'b10111110_01001010_00001000_1;
      patterns[48717] = 25'b10111110_01001011_00001001_1;
      patterns[48718] = 25'b10111110_01001100_00001010_1;
      patterns[48719] = 25'b10111110_01001101_00001011_1;
      patterns[48720] = 25'b10111110_01001110_00001100_1;
      patterns[48721] = 25'b10111110_01001111_00001101_1;
      patterns[48722] = 25'b10111110_01010000_00001110_1;
      patterns[48723] = 25'b10111110_01010001_00001111_1;
      patterns[48724] = 25'b10111110_01010010_00010000_1;
      patterns[48725] = 25'b10111110_01010011_00010001_1;
      patterns[48726] = 25'b10111110_01010100_00010010_1;
      patterns[48727] = 25'b10111110_01010101_00010011_1;
      patterns[48728] = 25'b10111110_01010110_00010100_1;
      patterns[48729] = 25'b10111110_01010111_00010101_1;
      patterns[48730] = 25'b10111110_01011000_00010110_1;
      patterns[48731] = 25'b10111110_01011001_00010111_1;
      patterns[48732] = 25'b10111110_01011010_00011000_1;
      patterns[48733] = 25'b10111110_01011011_00011001_1;
      patterns[48734] = 25'b10111110_01011100_00011010_1;
      patterns[48735] = 25'b10111110_01011101_00011011_1;
      patterns[48736] = 25'b10111110_01011110_00011100_1;
      patterns[48737] = 25'b10111110_01011111_00011101_1;
      patterns[48738] = 25'b10111110_01100000_00011110_1;
      patterns[48739] = 25'b10111110_01100001_00011111_1;
      patterns[48740] = 25'b10111110_01100010_00100000_1;
      patterns[48741] = 25'b10111110_01100011_00100001_1;
      patterns[48742] = 25'b10111110_01100100_00100010_1;
      patterns[48743] = 25'b10111110_01100101_00100011_1;
      patterns[48744] = 25'b10111110_01100110_00100100_1;
      patterns[48745] = 25'b10111110_01100111_00100101_1;
      patterns[48746] = 25'b10111110_01101000_00100110_1;
      patterns[48747] = 25'b10111110_01101001_00100111_1;
      patterns[48748] = 25'b10111110_01101010_00101000_1;
      patterns[48749] = 25'b10111110_01101011_00101001_1;
      patterns[48750] = 25'b10111110_01101100_00101010_1;
      patterns[48751] = 25'b10111110_01101101_00101011_1;
      patterns[48752] = 25'b10111110_01101110_00101100_1;
      patterns[48753] = 25'b10111110_01101111_00101101_1;
      patterns[48754] = 25'b10111110_01110000_00101110_1;
      patterns[48755] = 25'b10111110_01110001_00101111_1;
      patterns[48756] = 25'b10111110_01110010_00110000_1;
      patterns[48757] = 25'b10111110_01110011_00110001_1;
      patterns[48758] = 25'b10111110_01110100_00110010_1;
      patterns[48759] = 25'b10111110_01110101_00110011_1;
      patterns[48760] = 25'b10111110_01110110_00110100_1;
      patterns[48761] = 25'b10111110_01110111_00110101_1;
      patterns[48762] = 25'b10111110_01111000_00110110_1;
      patterns[48763] = 25'b10111110_01111001_00110111_1;
      patterns[48764] = 25'b10111110_01111010_00111000_1;
      patterns[48765] = 25'b10111110_01111011_00111001_1;
      patterns[48766] = 25'b10111110_01111100_00111010_1;
      patterns[48767] = 25'b10111110_01111101_00111011_1;
      patterns[48768] = 25'b10111110_01111110_00111100_1;
      patterns[48769] = 25'b10111110_01111111_00111101_1;
      patterns[48770] = 25'b10111110_10000000_00111110_1;
      patterns[48771] = 25'b10111110_10000001_00111111_1;
      patterns[48772] = 25'b10111110_10000010_01000000_1;
      patterns[48773] = 25'b10111110_10000011_01000001_1;
      patterns[48774] = 25'b10111110_10000100_01000010_1;
      patterns[48775] = 25'b10111110_10000101_01000011_1;
      patterns[48776] = 25'b10111110_10000110_01000100_1;
      patterns[48777] = 25'b10111110_10000111_01000101_1;
      patterns[48778] = 25'b10111110_10001000_01000110_1;
      patterns[48779] = 25'b10111110_10001001_01000111_1;
      patterns[48780] = 25'b10111110_10001010_01001000_1;
      patterns[48781] = 25'b10111110_10001011_01001001_1;
      patterns[48782] = 25'b10111110_10001100_01001010_1;
      patterns[48783] = 25'b10111110_10001101_01001011_1;
      patterns[48784] = 25'b10111110_10001110_01001100_1;
      patterns[48785] = 25'b10111110_10001111_01001101_1;
      patterns[48786] = 25'b10111110_10010000_01001110_1;
      patterns[48787] = 25'b10111110_10010001_01001111_1;
      patterns[48788] = 25'b10111110_10010010_01010000_1;
      patterns[48789] = 25'b10111110_10010011_01010001_1;
      patterns[48790] = 25'b10111110_10010100_01010010_1;
      patterns[48791] = 25'b10111110_10010101_01010011_1;
      patterns[48792] = 25'b10111110_10010110_01010100_1;
      patterns[48793] = 25'b10111110_10010111_01010101_1;
      patterns[48794] = 25'b10111110_10011000_01010110_1;
      patterns[48795] = 25'b10111110_10011001_01010111_1;
      patterns[48796] = 25'b10111110_10011010_01011000_1;
      patterns[48797] = 25'b10111110_10011011_01011001_1;
      patterns[48798] = 25'b10111110_10011100_01011010_1;
      patterns[48799] = 25'b10111110_10011101_01011011_1;
      patterns[48800] = 25'b10111110_10011110_01011100_1;
      patterns[48801] = 25'b10111110_10011111_01011101_1;
      patterns[48802] = 25'b10111110_10100000_01011110_1;
      patterns[48803] = 25'b10111110_10100001_01011111_1;
      patterns[48804] = 25'b10111110_10100010_01100000_1;
      patterns[48805] = 25'b10111110_10100011_01100001_1;
      patterns[48806] = 25'b10111110_10100100_01100010_1;
      patterns[48807] = 25'b10111110_10100101_01100011_1;
      patterns[48808] = 25'b10111110_10100110_01100100_1;
      patterns[48809] = 25'b10111110_10100111_01100101_1;
      patterns[48810] = 25'b10111110_10101000_01100110_1;
      patterns[48811] = 25'b10111110_10101001_01100111_1;
      patterns[48812] = 25'b10111110_10101010_01101000_1;
      patterns[48813] = 25'b10111110_10101011_01101001_1;
      patterns[48814] = 25'b10111110_10101100_01101010_1;
      patterns[48815] = 25'b10111110_10101101_01101011_1;
      patterns[48816] = 25'b10111110_10101110_01101100_1;
      patterns[48817] = 25'b10111110_10101111_01101101_1;
      patterns[48818] = 25'b10111110_10110000_01101110_1;
      patterns[48819] = 25'b10111110_10110001_01101111_1;
      patterns[48820] = 25'b10111110_10110010_01110000_1;
      patterns[48821] = 25'b10111110_10110011_01110001_1;
      patterns[48822] = 25'b10111110_10110100_01110010_1;
      patterns[48823] = 25'b10111110_10110101_01110011_1;
      patterns[48824] = 25'b10111110_10110110_01110100_1;
      patterns[48825] = 25'b10111110_10110111_01110101_1;
      patterns[48826] = 25'b10111110_10111000_01110110_1;
      patterns[48827] = 25'b10111110_10111001_01110111_1;
      patterns[48828] = 25'b10111110_10111010_01111000_1;
      patterns[48829] = 25'b10111110_10111011_01111001_1;
      patterns[48830] = 25'b10111110_10111100_01111010_1;
      patterns[48831] = 25'b10111110_10111101_01111011_1;
      patterns[48832] = 25'b10111110_10111110_01111100_1;
      patterns[48833] = 25'b10111110_10111111_01111101_1;
      patterns[48834] = 25'b10111110_11000000_01111110_1;
      patterns[48835] = 25'b10111110_11000001_01111111_1;
      patterns[48836] = 25'b10111110_11000010_10000000_1;
      patterns[48837] = 25'b10111110_11000011_10000001_1;
      patterns[48838] = 25'b10111110_11000100_10000010_1;
      patterns[48839] = 25'b10111110_11000101_10000011_1;
      patterns[48840] = 25'b10111110_11000110_10000100_1;
      patterns[48841] = 25'b10111110_11000111_10000101_1;
      patterns[48842] = 25'b10111110_11001000_10000110_1;
      patterns[48843] = 25'b10111110_11001001_10000111_1;
      patterns[48844] = 25'b10111110_11001010_10001000_1;
      patterns[48845] = 25'b10111110_11001011_10001001_1;
      patterns[48846] = 25'b10111110_11001100_10001010_1;
      patterns[48847] = 25'b10111110_11001101_10001011_1;
      patterns[48848] = 25'b10111110_11001110_10001100_1;
      patterns[48849] = 25'b10111110_11001111_10001101_1;
      patterns[48850] = 25'b10111110_11010000_10001110_1;
      patterns[48851] = 25'b10111110_11010001_10001111_1;
      patterns[48852] = 25'b10111110_11010010_10010000_1;
      patterns[48853] = 25'b10111110_11010011_10010001_1;
      patterns[48854] = 25'b10111110_11010100_10010010_1;
      patterns[48855] = 25'b10111110_11010101_10010011_1;
      patterns[48856] = 25'b10111110_11010110_10010100_1;
      patterns[48857] = 25'b10111110_11010111_10010101_1;
      patterns[48858] = 25'b10111110_11011000_10010110_1;
      patterns[48859] = 25'b10111110_11011001_10010111_1;
      patterns[48860] = 25'b10111110_11011010_10011000_1;
      patterns[48861] = 25'b10111110_11011011_10011001_1;
      patterns[48862] = 25'b10111110_11011100_10011010_1;
      patterns[48863] = 25'b10111110_11011101_10011011_1;
      patterns[48864] = 25'b10111110_11011110_10011100_1;
      patterns[48865] = 25'b10111110_11011111_10011101_1;
      patterns[48866] = 25'b10111110_11100000_10011110_1;
      patterns[48867] = 25'b10111110_11100001_10011111_1;
      patterns[48868] = 25'b10111110_11100010_10100000_1;
      patterns[48869] = 25'b10111110_11100011_10100001_1;
      patterns[48870] = 25'b10111110_11100100_10100010_1;
      patterns[48871] = 25'b10111110_11100101_10100011_1;
      patterns[48872] = 25'b10111110_11100110_10100100_1;
      patterns[48873] = 25'b10111110_11100111_10100101_1;
      patterns[48874] = 25'b10111110_11101000_10100110_1;
      patterns[48875] = 25'b10111110_11101001_10100111_1;
      patterns[48876] = 25'b10111110_11101010_10101000_1;
      patterns[48877] = 25'b10111110_11101011_10101001_1;
      patterns[48878] = 25'b10111110_11101100_10101010_1;
      patterns[48879] = 25'b10111110_11101101_10101011_1;
      patterns[48880] = 25'b10111110_11101110_10101100_1;
      patterns[48881] = 25'b10111110_11101111_10101101_1;
      patterns[48882] = 25'b10111110_11110000_10101110_1;
      patterns[48883] = 25'b10111110_11110001_10101111_1;
      patterns[48884] = 25'b10111110_11110010_10110000_1;
      patterns[48885] = 25'b10111110_11110011_10110001_1;
      patterns[48886] = 25'b10111110_11110100_10110010_1;
      patterns[48887] = 25'b10111110_11110101_10110011_1;
      patterns[48888] = 25'b10111110_11110110_10110100_1;
      patterns[48889] = 25'b10111110_11110111_10110101_1;
      patterns[48890] = 25'b10111110_11111000_10110110_1;
      patterns[48891] = 25'b10111110_11111001_10110111_1;
      patterns[48892] = 25'b10111110_11111010_10111000_1;
      patterns[48893] = 25'b10111110_11111011_10111001_1;
      patterns[48894] = 25'b10111110_11111100_10111010_1;
      patterns[48895] = 25'b10111110_11111101_10111011_1;
      patterns[48896] = 25'b10111110_11111110_10111100_1;
      patterns[48897] = 25'b10111110_11111111_10111101_1;
      patterns[48898] = 25'b10111111_00000000_10111111_0;
      patterns[48899] = 25'b10111111_00000001_11000000_0;
      patterns[48900] = 25'b10111111_00000010_11000001_0;
      patterns[48901] = 25'b10111111_00000011_11000010_0;
      patterns[48902] = 25'b10111111_00000100_11000011_0;
      patterns[48903] = 25'b10111111_00000101_11000100_0;
      patterns[48904] = 25'b10111111_00000110_11000101_0;
      patterns[48905] = 25'b10111111_00000111_11000110_0;
      patterns[48906] = 25'b10111111_00001000_11000111_0;
      patterns[48907] = 25'b10111111_00001001_11001000_0;
      patterns[48908] = 25'b10111111_00001010_11001001_0;
      patterns[48909] = 25'b10111111_00001011_11001010_0;
      patterns[48910] = 25'b10111111_00001100_11001011_0;
      patterns[48911] = 25'b10111111_00001101_11001100_0;
      patterns[48912] = 25'b10111111_00001110_11001101_0;
      patterns[48913] = 25'b10111111_00001111_11001110_0;
      patterns[48914] = 25'b10111111_00010000_11001111_0;
      patterns[48915] = 25'b10111111_00010001_11010000_0;
      patterns[48916] = 25'b10111111_00010010_11010001_0;
      patterns[48917] = 25'b10111111_00010011_11010010_0;
      patterns[48918] = 25'b10111111_00010100_11010011_0;
      patterns[48919] = 25'b10111111_00010101_11010100_0;
      patterns[48920] = 25'b10111111_00010110_11010101_0;
      patterns[48921] = 25'b10111111_00010111_11010110_0;
      patterns[48922] = 25'b10111111_00011000_11010111_0;
      patterns[48923] = 25'b10111111_00011001_11011000_0;
      patterns[48924] = 25'b10111111_00011010_11011001_0;
      patterns[48925] = 25'b10111111_00011011_11011010_0;
      patterns[48926] = 25'b10111111_00011100_11011011_0;
      patterns[48927] = 25'b10111111_00011101_11011100_0;
      patterns[48928] = 25'b10111111_00011110_11011101_0;
      patterns[48929] = 25'b10111111_00011111_11011110_0;
      patterns[48930] = 25'b10111111_00100000_11011111_0;
      patterns[48931] = 25'b10111111_00100001_11100000_0;
      patterns[48932] = 25'b10111111_00100010_11100001_0;
      patterns[48933] = 25'b10111111_00100011_11100010_0;
      patterns[48934] = 25'b10111111_00100100_11100011_0;
      patterns[48935] = 25'b10111111_00100101_11100100_0;
      patterns[48936] = 25'b10111111_00100110_11100101_0;
      patterns[48937] = 25'b10111111_00100111_11100110_0;
      patterns[48938] = 25'b10111111_00101000_11100111_0;
      patterns[48939] = 25'b10111111_00101001_11101000_0;
      patterns[48940] = 25'b10111111_00101010_11101001_0;
      patterns[48941] = 25'b10111111_00101011_11101010_0;
      patterns[48942] = 25'b10111111_00101100_11101011_0;
      patterns[48943] = 25'b10111111_00101101_11101100_0;
      patterns[48944] = 25'b10111111_00101110_11101101_0;
      patterns[48945] = 25'b10111111_00101111_11101110_0;
      patterns[48946] = 25'b10111111_00110000_11101111_0;
      patterns[48947] = 25'b10111111_00110001_11110000_0;
      patterns[48948] = 25'b10111111_00110010_11110001_0;
      patterns[48949] = 25'b10111111_00110011_11110010_0;
      patterns[48950] = 25'b10111111_00110100_11110011_0;
      patterns[48951] = 25'b10111111_00110101_11110100_0;
      patterns[48952] = 25'b10111111_00110110_11110101_0;
      patterns[48953] = 25'b10111111_00110111_11110110_0;
      patterns[48954] = 25'b10111111_00111000_11110111_0;
      patterns[48955] = 25'b10111111_00111001_11111000_0;
      patterns[48956] = 25'b10111111_00111010_11111001_0;
      patterns[48957] = 25'b10111111_00111011_11111010_0;
      patterns[48958] = 25'b10111111_00111100_11111011_0;
      patterns[48959] = 25'b10111111_00111101_11111100_0;
      patterns[48960] = 25'b10111111_00111110_11111101_0;
      patterns[48961] = 25'b10111111_00111111_11111110_0;
      patterns[48962] = 25'b10111111_01000000_11111111_0;
      patterns[48963] = 25'b10111111_01000001_00000000_1;
      patterns[48964] = 25'b10111111_01000010_00000001_1;
      patterns[48965] = 25'b10111111_01000011_00000010_1;
      patterns[48966] = 25'b10111111_01000100_00000011_1;
      patterns[48967] = 25'b10111111_01000101_00000100_1;
      patterns[48968] = 25'b10111111_01000110_00000101_1;
      patterns[48969] = 25'b10111111_01000111_00000110_1;
      patterns[48970] = 25'b10111111_01001000_00000111_1;
      patterns[48971] = 25'b10111111_01001001_00001000_1;
      patterns[48972] = 25'b10111111_01001010_00001001_1;
      patterns[48973] = 25'b10111111_01001011_00001010_1;
      patterns[48974] = 25'b10111111_01001100_00001011_1;
      patterns[48975] = 25'b10111111_01001101_00001100_1;
      patterns[48976] = 25'b10111111_01001110_00001101_1;
      patterns[48977] = 25'b10111111_01001111_00001110_1;
      patterns[48978] = 25'b10111111_01010000_00001111_1;
      patterns[48979] = 25'b10111111_01010001_00010000_1;
      patterns[48980] = 25'b10111111_01010010_00010001_1;
      patterns[48981] = 25'b10111111_01010011_00010010_1;
      patterns[48982] = 25'b10111111_01010100_00010011_1;
      patterns[48983] = 25'b10111111_01010101_00010100_1;
      patterns[48984] = 25'b10111111_01010110_00010101_1;
      patterns[48985] = 25'b10111111_01010111_00010110_1;
      patterns[48986] = 25'b10111111_01011000_00010111_1;
      patterns[48987] = 25'b10111111_01011001_00011000_1;
      patterns[48988] = 25'b10111111_01011010_00011001_1;
      patterns[48989] = 25'b10111111_01011011_00011010_1;
      patterns[48990] = 25'b10111111_01011100_00011011_1;
      patterns[48991] = 25'b10111111_01011101_00011100_1;
      patterns[48992] = 25'b10111111_01011110_00011101_1;
      patterns[48993] = 25'b10111111_01011111_00011110_1;
      patterns[48994] = 25'b10111111_01100000_00011111_1;
      patterns[48995] = 25'b10111111_01100001_00100000_1;
      patterns[48996] = 25'b10111111_01100010_00100001_1;
      patterns[48997] = 25'b10111111_01100011_00100010_1;
      patterns[48998] = 25'b10111111_01100100_00100011_1;
      patterns[48999] = 25'b10111111_01100101_00100100_1;
      patterns[49000] = 25'b10111111_01100110_00100101_1;
      patterns[49001] = 25'b10111111_01100111_00100110_1;
      patterns[49002] = 25'b10111111_01101000_00100111_1;
      patterns[49003] = 25'b10111111_01101001_00101000_1;
      patterns[49004] = 25'b10111111_01101010_00101001_1;
      patterns[49005] = 25'b10111111_01101011_00101010_1;
      patterns[49006] = 25'b10111111_01101100_00101011_1;
      patterns[49007] = 25'b10111111_01101101_00101100_1;
      patterns[49008] = 25'b10111111_01101110_00101101_1;
      patterns[49009] = 25'b10111111_01101111_00101110_1;
      patterns[49010] = 25'b10111111_01110000_00101111_1;
      patterns[49011] = 25'b10111111_01110001_00110000_1;
      patterns[49012] = 25'b10111111_01110010_00110001_1;
      patterns[49013] = 25'b10111111_01110011_00110010_1;
      patterns[49014] = 25'b10111111_01110100_00110011_1;
      patterns[49015] = 25'b10111111_01110101_00110100_1;
      patterns[49016] = 25'b10111111_01110110_00110101_1;
      patterns[49017] = 25'b10111111_01110111_00110110_1;
      patterns[49018] = 25'b10111111_01111000_00110111_1;
      patterns[49019] = 25'b10111111_01111001_00111000_1;
      patterns[49020] = 25'b10111111_01111010_00111001_1;
      patterns[49021] = 25'b10111111_01111011_00111010_1;
      patterns[49022] = 25'b10111111_01111100_00111011_1;
      patterns[49023] = 25'b10111111_01111101_00111100_1;
      patterns[49024] = 25'b10111111_01111110_00111101_1;
      patterns[49025] = 25'b10111111_01111111_00111110_1;
      patterns[49026] = 25'b10111111_10000000_00111111_1;
      patterns[49027] = 25'b10111111_10000001_01000000_1;
      patterns[49028] = 25'b10111111_10000010_01000001_1;
      patterns[49029] = 25'b10111111_10000011_01000010_1;
      patterns[49030] = 25'b10111111_10000100_01000011_1;
      patterns[49031] = 25'b10111111_10000101_01000100_1;
      patterns[49032] = 25'b10111111_10000110_01000101_1;
      patterns[49033] = 25'b10111111_10000111_01000110_1;
      patterns[49034] = 25'b10111111_10001000_01000111_1;
      patterns[49035] = 25'b10111111_10001001_01001000_1;
      patterns[49036] = 25'b10111111_10001010_01001001_1;
      patterns[49037] = 25'b10111111_10001011_01001010_1;
      patterns[49038] = 25'b10111111_10001100_01001011_1;
      patterns[49039] = 25'b10111111_10001101_01001100_1;
      patterns[49040] = 25'b10111111_10001110_01001101_1;
      patterns[49041] = 25'b10111111_10001111_01001110_1;
      patterns[49042] = 25'b10111111_10010000_01001111_1;
      patterns[49043] = 25'b10111111_10010001_01010000_1;
      patterns[49044] = 25'b10111111_10010010_01010001_1;
      patterns[49045] = 25'b10111111_10010011_01010010_1;
      patterns[49046] = 25'b10111111_10010100_01010011_1;
      patterns[49047] = 25'b10111111_10010101_01010100_1;
      patterns[49048] = 25'b10111111_10010110_01010101_1;
      patterns[49049] = 25'b10111111_10010111_01010110_1;
      patterns[49050] = 25'b10111111_10011000_01010111_1;
      patterns[49051] = 25'b10111111_10011001_01011000_1;
      patterns[49052] = 25'b10111111_10011010_01011001_1;
      patterns[49053] = 25'b10111111_10011011_01011010_1;
      patterns[49054] = 25'b10111111_10011100_01011011_1;
      patterns[49055] = 25'b10111111_10011101_01011100_1;
      patterns[49056] = 25'b10111111_10011110_01011101_1;
      patterns[49057] = 25'b10111111_10011111_01011110_1;
      patterns[49058] = 25'b10111111_10100000_01011111_1;
      patterns[49059] = 25'b10111111_10100001_01100000_1;
      patterns[49060] = 25'b10111111_10100010_01100001_1;
      patterns[49061] = 25'b10111111_10100011_01100010_1;
      patterns[49062] = 25'b10111111_10100100_01100011_1;
      patterns[49063] = 25'b10111111_10100101_01100100_1;
      patterns[49064] = 25'b10111111_10100110_01100101_1;
      patterns[49065] = 25'b10111111_10100111_01100110_1;
      patterns[49066] = 25'b10111111_10101000_01100111_1;
      patterns[49067] = 25'b10111111_10101001_01101000_1;
      patterns[49068] = 25'b10111111_10101010_01101001_1;
      patterns[49069] = 25'b10111111_10101011_01101010_1;
      patterns[49070] = 25'b10111111_10101100_01101011_1;
      patterns[49071] = 25'b10111111_10101101_01101100_1;
      patterns[49072] = 25'b10111111_10101110_01101101_1;
      patterns[49073] = 25'b10111111_10101111_01101110_1;
      patterns[49074] = 25'b10111111_10110000_01101111_1;
      patterns[49075] = 25'b10111111_10110001_01110000_1;
      patterns[49076] = 25'b10111111_10110010_01110001_1;
      patterns[49077] = 25'b10111111_10110011_01110010_1;
      patterns[49078] = 25'b10111111_10110100_01110011_1;
      patterns[49079] = 25'b10111111_10110101_01110100_1;
      patterns[49080] = 25'b10111111_10110110_01110101_1;
      patterns[49081] = 25'b10111111_10110111_01110110_1;
      patterns[49082] = 25'b10111111_10111000_01110111_1;
      patterns[49083] = 25'b10111111_10111001_01111000_1;
      patterns[49084] = 25'b10111111_10111010_01111001_1;
      patterns[49085] = 25'b10111111_10111011_01111010_1;
      patterns[49086] = 25'b10111111_10111100_01111011_1;
      patterns[49087] = 25'b10111111_10111101_01111100_1;
      patterns[49088] = 25'b10111111_10111110_01111101_1;
      patterns[49089] = 25'b10111111_10111111_01111110_1;
      patterns[49090] = 25'b10111111_11000000_01111111_1;
      patterns[49091] = 25'b10111111_11000001_10000000_1;
      patterns[49092] = 25'b10111111_11000010_10000001_1;
      patterns[49093] = 25'b10111111_11000011_10000010_1;
      patterns[49094] = 25'b10111111_11000100_10000011_1;
      patterns[49095] = 25'b10111111_11000101_10000100_1;
      patterns[49096] = 25'b10111111_11000110_10000101_1;
      patterns[49097] = 25'b10111111_11000111_10000110_1;
      patterns[49098] = 25'b10111111_11001000_10000111_1;
      patterns[49099] = 25'b10111111_11001001_10001000_1;
      patterns[49100] = 25'b10111111_11001010_10001001_1;
      patterns[49101] = 25'b10111111_11001011_10001010_1;
      patterns[49102] = 25'b10111111_11001100_10001011_1;
      patterns[49103] = 25'b10111111_11001101_10001100_1;
      patterns[49104] = 25'b10111111_11001110_10001101_1;
      patterns[49105] = 25'b10111111_11001111_10001110_1;
      patterns[49106] = 25'b10111111_11010000_10001111_1;
      patterns[49107] = 25'b10111111_11010001_10010000_1;
      patterns[49108] = 25'b10111111_11010010_10010001_1;
      patterns[49109] = 25'b10111111_11010011_10010010_1;
      patterns[49110] = 25'b10111111_11010100_10010011_1;
      patterns[49111] = 25'b10111111_11010101_10010100_1;
      patterns[49112] = 25'b10111111_11010110_10010101_1;
      patterns[49113] = 25'b10111111_11010111_10010110_1;
      patterns[49114] = 25'b10111111_11011000_10010111_1;
      patterns[49115] = 25'b10111111_11011001_10011000_1;
      patterns[49116] = 25'b10111111_11011010_10011001_1;
      patterns[49117] = 25'b10111111_11011011_10011010_1;
      patterns[49118] = 25'b10111111_11011100_10011011_1;
      patterns[49119] = 25'b10111111_11011101_10011100_1;
      patterns[49120] = 25'b10111111_11011110_10011101_1;
      patterns[49121] = 25'b10111111_11011111_10011110_1;
      patterns[49122] = 25'b10111111_11100000_10011111_1;
      patterns[49123] = 25'b10111111_11100001_10100000_1;
      patterns[49124] = 25'b10111111_11100010_10100001_1;
      patterns[49125] = 25'b10111111_11100011_10100010_1;
      patterns[49126] = 25'b10111111_11100100_10100011_1;
      patterns[49127] = 25'b10111111_11100101_10100100_1;
      patterns[49128] = 25'b10111111_11100110_10100101_1;
      patterns[49129] = 25'b10111111_11100111_10100110_1;
      patterns[49130] = 25'b10111111_11101000_10100111_1;
      patterns[49131] = 25'b10111111_11101001_10101000_1;
      patterns[49132] = 25'b10111111_11101010_10101001_1;
      patterns[49133] = 25'b10111111_11101011_10101010_1;
      patterns[49134] = 25'b10111111_11101100_10101011_1;
      patterns[49135] = 25'b10111111_11101101_10101100_1;
      patterns[49136] = 25'b10111111_11101110_10101101_1;
      patterns[49137] = 25'b10111111_11101111_10101110_1;
      patterns[49138] = 25'b10111111_11110000_10101111_1;
      patterns[49139] = 25'b10111111_11110001_10110000_1;
      patterns[49140] = 25'b10111111_11110010_10110001_1;
      patterns[49141] = 25'b10111111_11110011_10110010_1;
      patterns[49142] = 25'b10111111_11110100_10110011_1;
      patterns[49143] = 25'b10111111_11110101_10110100_1;
      patterns[49144] = 25'b10111111_11110110_10110101_1;
      patterns[49145] = 25'b10111111_11110111_10110110_1;
      patterns[49146] = 25'b10111111_11111000_10110111_1;
      patterns[49147] = 25'b10111111_11111001_10111000_1;
      patterns[49148] = 25'b10111111_11111010_10111001_1;
      patterns[49149] = 25'b10111111_11111011_10111010_1;
      patterns[49150] = 25'b10111111_11111100_10111011_1;
      patterns[49151] = 25'b10111111_11111101_10111100_1;
      patterns[49152] = 25'b10111111_11111110_10111101_1;
      patterns[49153] = 25'b10111111_11111111_10111110_1;
      patterns[49154] = 25'b11000000_00000000_11000000_0;
      patterns[49155] = 25'b11000000_00000001_11000001_0;
      patterns[49156] = 25'b11000000_00000010_11000010_0;
      patterns[49157] = 25'b11000000_00000011_11000011_0;
      patterns[49158] = 25'b11000000_00000100_11000100_0;
      patterns[49159] = 25'b11000000_00000101_11000101_0;
      patterns[49160] = 25'b11000000_00000110_11000110_0;
      patterns[49161] = 25'b11000000_00000111_11000111_0;
      patterns[49162] = 25'b11000000_00001000_11001000_0;
      patterns[49163] = 25'b11000000_00001001_11001001_0;
      patterns[49164] = 25'b11000000_00001010_11001010_0;
      patterns[49165] = 25'b11000000_00001011_11001011_0;
      patterns[49166] = 25'b11000000_00001100_11001100_0;
      patterns[49167] = 25'b11000000_00001101_11001101_0;
      patterns[49168] = 25'b11000000_00001110_11001110_0;
      patterns[49169] = 25'b11000000_00001111_11001111_0;
      patterns[49170] = 25'b11000000_00010000_11010000_0;
      patterns[49171] = 25'b11000000_00010001_11010001_0;
      patterns[49172] = 25'b11000000_00010010_11010010_0;
      patterns[49173] = 25'b11000000_00010011_11010011_0;
      patterns[49174] = 25'b11000000_00010100_11010100_0;
      patterns[49175] = 25'b11000000_00010101_11010101_0;
      patterns[49176] = 25'b11000000_00010110_11010110_0;
      patterns[49177] = 25'b11000000_00010111_11010111_0;
      patterns[49178] = 25'b11000000_00011000_11011000_0;
      patterns[49179] = 25'b11000000_00011001_11011001_0;
      patterns[49180] = 25'b11000000_00011010_11011010_0;
      patterns[49181] = 25'b11000000_00011011_11011011_0;
      patterns[49182] = 25'b11000000_00011100_11011100_0;
      patterns[49183] = 25'b11000000_00011101_11011101_0;
      patterns[49184] = 25'b11000000_00011110_11011110_0;
      patterns[49185] = 25'b11000000_00011111_11011111_0;
      patterns[49186] = 25'b11000000_00100000_11100000_0;
      patterns[49187] = 25'b11000000_00100001_11100001_0;
      patterns[49188] = 25'b11000000_00100010_11100010_0;
      patterns[49189] = 25'b11000000_00100011_11100011_0;
      patterns[49190] = 25'b11000000_00100100_11100100_0;
      patterns[49191] = 25'b11000000_00100101_11100101_0;
      patterns[49192] = 25'b11000000_00100110_11100110_0;
      patterns[49193] = 25'b11000000_00100111_11100111_0;
      patterns[49194] = 25'b11000000_00101000_11101000_0;
      patterns[49195] = 25'b11000000_00101001_11101001_0;
      patterns[49196] = 25'b11000000_00101010_11101010_0;
      patterns[49197] = 25'b11000000_00101011_11101011_0;
      patterns[49198] = 25'b11000000_00101100_11101100_0;
      patterns[49199] = 25'b11000000_00101101_11101101_0;
      patterns[49200] = 25'b11000000_00101110_11101110_0;
      patterns[49201] = 25'b11000000_00101111_11101111_0;
      patterns[49202] = 25'b11000000_00110000_11110000_0;
      patterns[49203] = 25'b11000000_00110001_11110001_0;
      patterns[49204] = 25'b11000000_00110010_11110010_0;
      patterns[49205] = 25'b11000000_00110011_11110011_0;
      patterns[49206] = 25'b11000000_00110100_11110100_0;
      patterns[49207] = 25'b11000000_00110101_11110101_0;
      patterns[49208] = 25'b11000000_00110110_11110110_0;
      patterns[49209] = 25'b11000000_00110111_11110111_0;
      patterns[49210] = 25'b11000000_00111000_11111000_0;
      patterns[49211] = 25'b11000000_00111001_11111001_0;
      patterns[49212] = 25'b11000000_00111010_11111010_0;
      patterns[49213] = 25'b11000000_00111011_11111011_0;
      patterns[49214] = 25'b11000000_00111100_11111100_0;
      patterns[49215] = 25'b11000000_00111101_11111101_0;
      patterns[49216] = 25'b11000000_00111110_11111110_0;
      patterns[49217] = 25'b11000000_00111111_11111111_0;
      patterns[49218] = 25'b11000000_01000000_00000000_1;
      patterns[49219] = 25'b11000000_01000001_00000001_1;
      patterns[49220] = 25'b11000000_01000010_00000010_1;
      patterns[49221] = 25'b11000000_01000011_00000011_1;
      patterns[49222] = 25'b11000000_01000100_00000100_1;
      patterns[49223] = 25'b11000000_01000101_00000101_1;
      patterns[49224] = 25'b11000000_01000110_00000110_1;
      patterns[49225] = 25'b11000000_01000111_00000111_1;
      patterns[49226] = 25'b11000000_01001000_00001000_1;
      patterns[49227] = 25'b11000000_01001001_00001001_1;
      patterns[49228] = 25'b11000000_01001010_00001010_1;
      patterns[49229] = 25'b11000000_01001011_00001011_1;
      patterns[49230] = 25'b11000000_01001100_00001100_1;
      patterns[49231] = 25'b11000000_01001101_00001101_1;
      patterns[49232] = 25'b11000000_01001110_00001110_1;
      patterns[49233] = 25'b11000000_01001111_00001111_1;
      patterns[49234] = 25'b11000000_01010000_00010000_1;
      patterns[49235] = 25'b11000000_01010001_00010001_1;
      patterns[49236] = 25'b11000000_01010010_00010010_1;
      patterns[49237] = 25'b11000000_01010011_00010011_1;
      patterns[49238] = 25'b11000000_01010100_00010100_1;
      patterns[49239] = 25'b11000000_01010101_00010101_1;
      patterns[49240] = 25'b11000000_01010110_00010110_1;
      patterns[49241] = 25'b11000000_01010111_00010111_1;
      patterns[49242] = 25'b11000000_01011000_00011000_1;
      patterns[49243] = 25'b11000000_01011001_00011001_1;
      patterns[49244] = 25'b11000000_01011010_00011010_1;
      patterns[49245] = 25'b11000000_01011011_00011011_1;
      patterns[49246] = 25'b11000000_01011100_00011100_1;
      patterns[49247] = 25'b11000000_01011101_00011101_1;
      patterns[49248] = 25'b11000000_01011110_00011110_1;
      patterns[49249] = 25'b11000000_01011111_00011111_1;
      patterns[49250] = 25'b11000000_01100000_00100000_1;
      patterns[49251] = 25'b11000000_01100001_00100001_1;
      patterns[49252] = 25'b11000000_01100010_00100010_1;
      patterns[49253] = 25'b11000000_01100011_00100011_1;
      patterns[49254] = 25'b11000000_01100100_00100100_1;
      patterns[49255] = 25'b11000000_01100101_00100101_1;
      patterns[49256] = 25'b11000000_01100110_00100110_1;
      patterns[49257] = 25'b11000000_01100111_00100111_1;
      patterns[49258] = 25'b11000000_01101000_00101000_1;
      patterns[49259] = 25'b11000000_01101001_00101001_1;
      patterns[49260] = 25'b11000000_01101010_00101010_1;
      patterns[49261] = 25'b11000000_01101011_00101011_1;
      patterns[49262] = 25'b11000000_01101100_00101100_1;
      patterns[49263] = 25'b11000000_01101101_00101101_1;
      patterns[49264] = 25'b11000000_01101110_00101110_1;
      patterns[49265] = 25'b11000000_01101111_00101111_1;
      patterns[49266] = 25'b11000000_01110000_00110000_1;
      patterns[49267] = 25'b11000000_01110001_00110001_1;
      patterns[49268] = 25'b11000000_01110010_00110010_1;
      patterns[49269] = 25'b11000000_01110011_00110011_1;
      patterns[49270] = 25'b11000000_01110100_00110100_1;
      patterns[49271] = 25'b11000000_01110101_00110101_1;
      patterns[49272] = 25'b11000000_01110110_00110110_1;
      patterns[49273] = 25'b11000000_01110111_00110111_1;
      patterns[49274] = 25'b11000000_01111000_00111000_1;
      patterns[49275] = 25'b11000000_01111001_00111001_1;
      patterns[49276] = 25'b11000000_01111010_00111010_1;
      patterns[49277] = 25'b11000000_01111011_00111011_1;
      patterns[49278] = 25'b11000000_01111100_00111100_1;
      patterns[49279] = 25'b11000000_01111101_00111101_1;
      patterns[49280] = 25'b11000000_01111110_00111110_1;
      patterns[49281] = 25'b11000000_01111111_00111111_1;
      patterns[49282] = 25'b11000000_10000000_01000000_1;
      patterns[49283] = 25'b11000000_10000001_01000001_1;
      patterns[49284] = 25'b11000000_10000010_01000010_1;
      patterns[49285] = 25'b11000000_10000011_01000011_1;
      patterns[49286] = 25'b11000000_10000100_01000100_1;
      patterns[49287] = 25'b11000000_10000101_01000101_1;
      patterns[49288] = 25'b11000000_10000110_01000110_1;
      patterns[49289] = 25'b11000000_10000111_01000111_1;
      patterns[49290] = 25'b11000000_10001000_01001000_1;
      patterns[49291] = 25'b11000000_10001001_01001001_1;
      patterns[49292] = 25'b11000000_10001010_01001010_1;
      patterns[49293] = 25'b11000000_10001011_01001011_1;
      patterns[49294] = 25'b11000000_10001100_01001100_1;
      patterns[49295] = 25'b11000000_10001101_01001101_1;
      patterns[49296] = 25'b11000000_10001110_01001110_1;
      patterns[49297] = 25'b11000000_10001111_01001111_1;
      patterns[49298] = 25'b11000000_10010000_01010000_1;
      patterns[49299] = 25'b11000000_10010001_01010001_1;
      patterns[49300] = 25'b11000000_10010010_01010010_1;
      patterns[49301] = 25'b11000000_10010011_01010011_1;
      patterns[49302] = 25'b11000000_10010100_01010100_1;
      patterns[49303] = 25'b11000000_10010101_01010101_1;
      patterns[49304] = 25'b11000000_10010110_01010110_1;
      patterns[49305] = 25'b11000000_10010111_01010111_1;
      patterns[49306] = 25'b11000000_10011000_01011000_1;
      patterns[49307] = 25'b11000000_10011001_01011001_1;
      patterns[49308] = 25'b11000000_10011010_01011010_1;
      patterns[49309] = 25'b11000000_10011011_01011011_1;
      patterns[49310] = 25'b11000000_10011100_01011100_1;
      patterns[49311] = 25'b11000000_10011101_01011101_1;
      patterns[49312] = 25'b11000000_10011110_01011110_1;
      patterns[49313] = 25'b11000000_10011111_01011111_1;
      patterns[49314] = 25'b11000000_10100000_01100000_1;
      patterns[49315] = 25'b11000000_10100001_01100001_1;
      patterns[49316] = 25'b11000000_10100010_01100010_1;
      patterns[49317] = 25'b11000000_10100011_01100011_1;
      patterns[49318] = 25'b11000000_10100100_01100100_1;
      patterns[49319] = 25'b11000000_10100101_01100101_1;
      patterns[49320] = 25'b11000000_10100110_01100110_1;
      patterns[49321] = 25'b11000000_10100111_01100111_1;
      patterns[49322] = 25'b11000000_10101000_01101000_1;
      patterns[49323] = 25'b11000000_10101001_01101001_1;
      patterns[49324] = 25'b11000000_10101010_01101010_1;
      patterns[49325] = 25'b11000000_10101011_01101011_1;
      patterns[49326] = 25'b11000000_10101100_01101100_1;
      patterns[49327] = 25'b11000000_10101101_01101101_1;
      patterns[49328] = 25'b11000000_10101110_01101110_1;
      patterns[49329] = 25'b11000000_10101111_01101111_1;
      patterns[49330] = 25'b11000000_10110000_01110000_1;
      patterns[49331] = 25'b11000000_10110001_01110001_1;
      patterns[49332] = 25'b11000000_10110010_01110010_1;
      patterns[49333] = 25'b11000000_10110011_01110011_1;
      patterns[49334] = 25'b11000000_10110100_01110100_1;
      patterns[49335] = 25'b11000000_10110101_01110101_1;
      patterns[49336] = 25'b11000000_10110110_01110110_1;
      patterns[49337] = 25'b11000000_10110111_01110111_1;
      patterns[49338] = 25'b11000000_10111000_01111000_1;
      patterns[49339] = 25'b11000000_10111001_01111001_1;
      patterns[49340] = 25'b11000000_10111010_01111010_1;
      patterns[49341] = 25'b11000000_10111011_01111011_1;
      patterns[49342] = 25'b11000000_10111100_01111100_1;
      patterns[49343] = 25'b11000000_10111101_01111101_1;
      patterns[49344] = 25'b11000000_10111110_01111110_1;
      patterns[49345] = 25'b11000000_10111111_01111111_1;
      patterns[49346] = 25'b11000000_11000000_10000000_1;
      patterns[49347] = 25'b11000000_11000001_10000001_1;
      patterns[49348] = 25'b11000000_11000010_10000010_1;
      patterns[49349] = 25'b11000000_11000011_10000011_1;
      patterns[49350] = 25'b11000000_11000100_10000100_1;
      patterns[49351] = 25'b11000000_11000101_10000101_1;
      patterns[49352] = 25'b11000000_11000110_10000110_1;
      patterns[49353] = 25'b11000000_11000111_10000111_1;
      patterns[49354] = 25'b11000000_11001000_10001000_1;
      patterns[49355] = 25'b11000000_11001001_10001001_1;
      patterns[49356] = 25'b11000000_11001010_10001010_1;
      patterns[49357] = 25'b11000000_11001011_10001011_1;
      patterns[49358] = 25'b11000000_11001100_10001100_1;
      patterns[49359] = 25'b11000000_11001101_10001101_1;
      patterns[49360] = 25'b11000000_11001110_10001110_1;
      patterns[49361] = 25'b11000000_11001111_10001111_1;
      patterns[49362] = 25'b11000000_11010000_10010000_1;
      patterns[49363] = 25'b11000000_11010001_10010001_1;
      patterns[49364] = 25'b11000000_11010010_10010010_1;
      patterns[49365] = 25'b11000000_11010011_10010011_1;
      patterns[49366] = 25'b11000000_11010100_10010100_1;
      patterns[49367] = 25'b11000000_11010101_10010101_1;
      patterns[49368] = 25'b11000000_11010110_10010110_1;
      patterns[49369] = 25'b11000000_11010111_10010111_1;
      patterns[49370] = 25'b11000000_11011000_10011000_1;
      patterns[49371] = 25'b11000000_11011001_10011001_1;
      patterns[49372] = 25'b11000000_11011010_10011010_1;
      patterns[49373] = 25'b11000000_11011011_10011011_1;
      patterns[49374] = 25'b11000000_11011100_10011100_1;
      patterns[49375] = 25'b11000000_11011101_10011101_1;
      patterns[49376] = 25'b11000000_11011110_10011110_1;
      patterns[49377] = 25'b11000000_11011111_10011111_1;
      patterns[49378] = 25'b11000000_11100000_10100000_1;
      patterns[49379] = 25'b11000000_11100001_10100001_1;
      patterns[49380] = 25'b11000000_11100010_10100010_1;
      patterns[49381] = 25'b11000000_11100011_10100011_1;
      patterns[49382] = 25'b11000000_11100100_10100100_1;
      patterns[49383] = 25'b11000000_11100101_10100101_1;
      patterns[49384] = 25'b11000000_11100110_10100110_1;
      patterns[49385] = 25'b11000000_11100111_10100111_1;
      patterns[49386] = 25'b11000000_11101000_10101000_1;
      patterns[49387] = 25'b11000000_11101001_10101001_1;
      patterns[49388] = 25'b11000000_11101010_10101010_1;
      patterns[49389] = 25'b11000000_11101011_10101011_1;
      patterns[49390] = 25'b11000000_11101100_10101100_1;
      patterns[49391] = 25'b11000000_11101101_10101101_1;
      patterns[49392] = 25'b11000000_11101110_10101110_1;
      patterns[49393] = 25'b11000000_11101111_10101111_1;
      patterns[49394] = 25'b11000000_11110000_10110000_1;
      patterns[49395] = 25'b11000000_11110001_10110001_1;
      patterns[49396] = 25'b11000000_11110010_10110010_1;
      patterns[49397] = 25'b11000000_11110011_10110011_1;
      patterns[49398] = 25'b11000000_11110100_10110100_1;
      patterns[49399] = 25'b11000000_11110101_10110101_1;
      patterns[49400] = 25'b11000000_11110110_10110110_1;
      patterns[49401] = 25'b11000000_11110111_10110111_1;
      patterns[49402] = 25'b11000000_11111000_10111000_1;
      patterns[49403] = 25'b11000000_11111001_10111001_1;
      patterns[49404] = 25'b11000000_11111010_10111010_1;
      patterns[49405] = 25'b11000000_11111011_10111011_1;
      patterns[49406] = 25'b11000000_11111100_10111100_1;
      patterns[49407] = 25'b11000000_11111101_10111101_1;
      patterns[49408] = 25'b11000000_11111110_10111110_1;
      patterns[49409] = 25'b11000000_11111111_10111111_1;
      patterns[49410] = 25'b11000001_00000000_11000001_0;
      patterns[49411] = 25'b11000001_00000001_11000010_0;
      patterns[49412] = 25'b11000001_00000010_11000011_0;
      patterns[49413] = 25'b11000001_00000011_11000100_0;
      patterns[49414] = 25'b11000001_00000100_11000101_0;
      patterns[49415] = 25'b11000001_00000101_11000110_0;
      patterns[49416] = 25'b11000001_00000110_11000111_0;
      patterns[49417] = 25'b11000001_00000111_11001000_0;
      patterns[49418] = 25'b11000001_00001000_11001001_0;
      patterns[49419] = 25'b11000001_00001001_11001010_0;
      patterns[49420] = 25'b11000001_00001010_11001011_0;
      patterns[49421] = 25'b11000001_00001011_11001100_0;
      patterns[49422] = 25'b11000001_00001100_11001101_0;
      patterns[49423] = 25'b11000001_00001101_11001110_0;
      patterns[49424] = 25'b11000001_00001110_11001111_0;
      patterns[49425] = 25'b11000001_00001111_11010000_0;
      patterns[49426] = 25'b11000001_00010000_11010001_0;
      patterns[49427] = 25'b11000001_00010001_11010010_0;
      patterns[49428] = 25'b11000001_00010010_11010011_0;
      patterns[49429] = 25'b11000001_00010011_11010100_0;
      patterns[49430] = 25'b11000001_00010100_11010101_0;
      patterns[49431] = 25'b11000001_00010101_11010110_0;
      patterns[49432] = 25'b11000001_00010110_11010111_0;
      patterns[49433] = 25'b11000001_00010111_11011000_0;
      patterns[49434] = 25'b11000001_00011000_11011001_0;
      patterns[49435] = 25'b11000001_00011001_11011010_0;
      patterns[49436] = 25'b11000001_00011010_11011011_0;
      patterns[49437] = 25'b11000001_00011011_11011100_0;
      patterns[49438] = 25'b11000001_00011100_11011101_0;
      patterns[49439] = 25'b11000001_00011101_11011110_0;
      patterns[49440] = 25'b11000001_00011110_11011111_0;
      patterns[49441] = 25'b11000001_00011111_11100000_0;
      patterns[49442] = 25'b11000001_00100000_11100001_0;
      patterns[49443] = 25'b11000001_00100001_11100010_0;
      patterns[49444] = 25'b11000001_00100010_11100011_0;
      patterns[49445] = 25'b11000001_00100011_11100100_0;
      patterns[49446] = 25'b11000001_00100100_11100101_0;
      patterns[49447] = 25'b11000001_00100101_11100110_0;
      patterns[49448] = 25'b11000001_00100110_11100111_0;
      patterns[49449] = 25'b11000001_00100111_11101000_0;
      patterns[49450] = 25'b11000001_00101000_11101001_0;
      patterns[49451] = 25'b11000001_00101001_11101010_0;
      patterns[49452] = 25'b11000001_00101010_11101011_0;
      patterns[49453] = 25'b11000001_00101011_11101100_0;
      patterns[49454] = 25'b11000001_00101100_11101101_0;
      patterns[49455] = 25'b11000001_00101101_11101110_0;
      patterns[49456] = 25'b11000001_00101110_11101111_0;
      patterns[49457] = 25'b11000001_00101111_11110000_0;
      patterns[49458] = 25'b11000001_00110000_11110001_0;
      patterns[49459] = 25'b11000001_00110001_11110010_0;
      patterns[49460] = 25'b11000001_00110010_11110011_0;
      patterns[49461] = 25'b11000001_00110011_11110100_0;
      patterns[49462] = 25'b11000001_00110100_11110101_0;
      patterns[49463] = 25'b11000001_00110101_11110110_0;
      patterns[49464] = 25'b11000001_00110110_11110111_0;
      patterns[49465] = 25'b11000001_00110111_11111000_0;
      patterns[49466] = 25'b11000001_00111000_11111001_0;
      patterns[49467] = 25'b11000001_00111001_11111010_0;
      patterns[49468] = 25'b11000001_00111010_11111011_0;
      patterns[49469] = 25'b11000001_00111011_11111100_0;
      patterns[49470] = 25'b11000001_00111100_11111101_0;
      patterns[49471] = 25'b11000001_00111101_11111110_0;
      patterns[49472] = 25'b11000001_00111110_11111111_0;
      patterns[49473] = 25'b11000001_00111111_00000000_1;
      patterns[49474] = 25'b11000001_01000000_00000001_1;
      patterns[49475] = 25'b11000001_01000001_00000010_1;
      patterns[49476] = 25'b11000001_01000010_00000011_1;
      patterns[49477] = 25'b11000001_01000011_00000100_1;
      patterns[49478] = 25'b11000001_01000100_00000101_1;
      patterns[49479] = 25'b11000001_01000101_00000110_1;
      patterns[49480] = 25'b11000001_01000110_00000111_1;
      patterns[49481] = 25'b11000001_01000111_00001000_1;
      patterns[49482] = 25'b11000001_01001000_00001001_1;
      patterns[49483] = 25'b11000001_01001001_00001010_1;
      patterns[49484] = 25'b11000001_01001010_00001011_1;
      patterns[49485] = 25'b11000001_01001011_00001100_1;
      patterns[49486] = 25'b11000001_01001100_00001101_1;
      patterns[49487] = 25'b11000001_01001101_00001110_1;
      patterns[49488] = 25'b11000001_01001110_00001111_1;
      patterns[49489] = 25'b11000001_01001111_00010000_1;
      patterns[49490] = 25'b11000001_01010000_00010001_1;
      patterns[49491] = 25'b11000001_01010001_00010010_1;
      patterns[49492] = 25'b11000001_01010010_00010011_1;
      patterns[49493] = 25'b11000001_01010011_00010100_1;
      patterns[49494] = 25'b11000001_01010100_00010101_1;
      patterns[49495] = 25'b11000001_01010101_00010110_1;
      patterns[49496] = 25'b11000001_01010110_00010111_1;
      patterns[49497] = 25'b11000001_01010111_00011000_1;
      patterns[49498] = 25'b11000001_01011000_00011001_1;
      patterns[49499] = 25'b11000001_01011001_00011010_1;
      patterns[49500] = 25'b11000001_01011010_00011011_1;
      patterns[49501] = 25'b11000001_01011011_00011100_1;
      patterns[49502] = 25'b11000001_01011100_00011101_1;
      patterns[49503] = 25'b11000001_01011101_00011110_1;
      patterns[49504] = 25'b11000001_01011110_00011111_1;
      patterns[49505] = 25'b11000001_01011111_00100000_1;
      patterns[49506] = 25'b11000001_01100000_00100001_1;
      patterns[49507] = 25'b11000001_01100001_00100010_1;
      patterns[49508] = 25'b11000001_01100010_00100011_1;
      patterns[49509] = 25'b11000001_01100011_00100100_1;
      patterns[49510] = 25'b11000001_01100100_00100101_1;
      patterns[49511] = 25'b11000001_01100101_00100110_1;
      patterns[49512] = 25'b11000001_01100110_00100111_1;
      patterns[49513] = 25'b11000001_01100111_00101000_1;
      patterns[49514] = 25'b11000001_01101000_00101001_1;
      patterns[49515] = 25'b11000001_01101001_00101010_1;
      patterns[49516] = 25'b11000001_01101010_00101011_1;
      patterns[49517] = 25'b11000001_01101011_00101100_1;
      patterns[49518] = 25'b11000001_01101100_00101101_1;
      patterns[49519] = 25'b11000001_01101101_00101110_1;
      patterns[49520] = 25'b11000001_01101110_00101111_1;
      patterns[49521] = 25'b11000001_01101111_00110000_1;
      patterns[49522] = 25'b11000001_01110000_00110001_1;
      patterns[49523] = 25'b11000001_01110001_00110010_1;
      patterns[49524] = 25'b11000001_01110010_00110011_1;
      patterns[49525] = 25'b11000001_01110011_00110100_1;
      patterns[49526] = 25'b11000001_01110100_00110101_1;
      patterns[49527] = 25'b11000001_01110101_00110110_1;
      patterns[49528] = 25'b11000001_01110110_00110111_1;
      patterns[49529] = 25'b11000001_01110111_00111000_1;
      patterns[49530] = 25'b11000001_01111000_00111001_1;
      patterns[49531] = 25'b11000001_01111001_00111010_1;
      patterns[49532] = 25'b11000001_01111010_00111011_1;
      patterns[49533] = 25'b11000001_01111011_00111100_1;
      patterns[49534] = 25'b11000001_01111100_00111101_1;
      patterns[49535] = 25'b11000001_01111101_00111110_1;
      patterns[49536] = 25'b11000001_01111110_00111111_1;
      patterns[49537] = 25'b11000001_01111111_01000000_1;
      patterns[49538] = 25'b11000001_10000000_01000001_1;
      patterns[49539] = 25'b11000001_10000001_01000010_1;
      patterns[49540] = 25'b11000001_10000010_01000011_1;
      patterns[49541] = 25'b11000001_10000011_01000100_1;
      patterns[49542] = 25'b11000001_10000100_01000101_1;
      patterns[49543] = 25'b11000001_10000101_01000110_1;
      patterns[49544] = 25'b11000001_10000110_01000111_1;
      patterns[49545] = 25'b11000001_10000111_01001000_1;
      patterns[49546] = 25'b11000001_10001000_01001001_1;
      patterns[49547] = 25'b11000001_10001001_01001010_1;
      patterns[49548] = 25'b11000001_10001010_01001011_1;
      patterns[49549] = 25'b11000001_10001011_01001100_1;
      patterns[49550] = 25'b11000001_10001100_01001101_1;
      patterns[49551] = 25'b11000001_10001101_01001110_1;
      patterns[49552] = 25'b11000001_10001110_01001111_1;
      patterns[49553] = 25'b11000001_10001111_01010000_1;
      patterns[49554] = 25'b11000001_10010000_01010001_1;
      patterns[49555] = 25'b11000001_10010001_01010010_1;
      patterns[49556] = 25'b11000001_10010010_01010011_1;
      patterns[49557] = 25'b11000001_10010011_01010100_1;
      patterns[49558] = 25'b11000001_10010100_01010101_1;
      patterns[49559] = 25'b11000001_10010101_01010110_1;
      patterns[49560] = 25'b11000001_10010110_01010111_1;
      patterns[49561] = 25'b11000001_10010111_01011000_1;
      patterns[49562] = 25'b11000001_10011000_01011001_1;
      patterns[49563] = 25'b11000001_10011001_01011010_1;
      patterns[49564] = 25'b11000001_10011010_01011011_1;
      patterns[49565] = 25'b11000001_10011011_01011100_1;
      patterns[49566] = 25'b11000001_10011100_01011101_1;
      patterns[49567] = 25'b11000001_10011101_01011110_1;
      patterns[49568] = 25'b11000001_10011110_01011111_1;
      patterns[49569] = 25'b11000001_10011111_01100000_1;
      patterns[49570] = 25'b11000001_10100000_01100001_1;
      patterns[49571] = 25'b11000001_10100001_01100010_1;
      patterns[49572] = 25'b11000001_10100010_01100011_1;
      patterns[49573] = 25'b11000001_10100011_01100100_1;
      patterns[49574] = 25'b11000001_10100100_01100101_1;
      patterns[49575] = 25'b11000001_10100101_01100110_1;
      patterns[49576] = 25'b11000001_10100110_01100111_1;
      patterns[49577] = 25'b11000001_10100111_01101000_1;
      patterns[49578] = 25'b11000001_10101000_01101001_1;
      patterns[49579] = 25'b11000001_10101001_01101010_1;
      patterns[49580] = 25'b11000001_10101010_01101011_1;
      patterns[49581] = 25'b11000001_10101011_01101100_1;
      patterns[49582] = 25'b11000001_10101100_01101101_1;
      patterns[49583] = 25'b11000001_10101101_01101110_1;
      patterns[49584] = 25'b11000001_10101110_01101111_1;
      patterns[49585] = 25'b11000001_10101111_01110000_1;
      patterns[49586] = 25'b11000001_10110000_01110001_1;
      patterns[49587] = 25'b11000001_10110001_01110010_1;
      patterns[49588] = 25'b11000001_10110010_01110011_1;
      patterns[49589] = 25'b11000001_10110011_01110100_1;
      patterns[49590] = 25'b11000001_10110100_01110101_1;
      patterns[49591] = 25'b11000001_10110101_01110110_1;
      patterns[49592] = 25'b11000001_10110110_01110111_1;
      patterns[49593] = 25'b11000001_10110111_01111000_1;
      patterns[49594] = 25'b11000001_10111000_01111001_1;
      patterns[49595] = 25'b11000001_10111001_01111010_1;
      patterns[49596] = 25'b11000001_10111010_01111011_1;
      patterns[49597] = 25'b11000001_10111011_01111100_1;
      patterns[49598] = 25'b11000001_10111100_01111101_1;
      patterns[49599] = 25'b11000001_10111101_01111110_1;
      patterns[49600] = 25'b11000001_10111110_01111111_1;
      patterns[49601] = 25'b11000001_10111111_10000000_1;
      patterns[49602] = 25'b11000001_11000000_10000001_1;
      patterns[49603] = 25'b11000001_11000001_10000010_1;
      patterns[49604] = 25'b11000001_11000010_10000011_1;
      patterns[49605] = 25'b11000001_11000011_10000100_1;
      patterns[49606] = 25'b11000001_11000100_10000101_1;
      patterns[49607] = 25'b11000001_11000101_10000110_1;
      patterns[49608] = 25'b11000001_11000110_10000111_1;
      patterns[49609] = 25'b11000001_11000111_10001000_1;
      patterns[49610] = 25'b11000001_11001000_10001001_1;
      patterns[49611] = 25'b11000001_11001001_10001010_1;
      patterns[49612] = 25'b11000001_11001010_10001011_1;
      patterns[49613] = 25'b11000001_11001011_10001100_1;
      patterns[49614] = 25'b11000001_11001100_10001101_1;
      patterns[49615] = 25'b11000001_11001101_10001110_1;
      patterns[49616] = 25'b11000001_11001110_10001111_1;
      patterns[49617] = 25'b11000001_11001111_10010000_1;
      patterns[49618] = 25'b11000001_11010000_10010001_1;
      patterns[49619] = 25'b11000001_11010001_10010010_1;
      patterns[49620] = 25'b11000001_11010010_10010011_1;
      patterns[49621] = 25'b11000001_11010011_10010100_1;
      patterns[49622] = 25'b11000001_11010100_10010101_1;
      patterns[49623] = 25'b11000001_11010101_10010110_1;
      patterns[49624] = 25'b11000001_11010110_10010111_1;
      patterns[49625] = 25'b11000001_11010111_10011000_1;
      patterns[49626] = 25'b11000001_11011000_10011001_1;
      patterns[49627] = 25'b11000001_11011001_10011010_1;
      patterns[49628] = 25'b11000001_11011010_10011011_1;
      patterns[49629] = 25'b11000001_11011011_10011100_1;
      patterns[49630] = 25'b11000001_11011100_10011101_1;
      patterns[49631] = 25'b11000001_11011101_10011110_1;
      patterns[49632] = 25'b11000001_11011110_10011111_1;
      patterns[49633] = 25'b11000001_11011111_10100000_1;
      patterns[49634] = 25'b11000001_11100000_10100001_1;
      patterns[49635] = 25'b11000001_11100001_10100010_1;
      patterns[49636] = 25'b11000001_11100010_10100011_1;
      patterns[49637] = 25'b11000001_11100011_10100100_1;
      patterns[49638] = 25'b11000001_11100100_10100101_1;
      patterns[49639] = 25'b11000001_11100101_10100110_1;
      patterns[49640] = 25'b11000001_11100110_10100111_1;
      patterns[49641] = 25'b11000001_11100111_10101000_1;
      patterns[49642] = 25'b11000001_11101000_10101001_1;
      patterns[49643] = 25'b11000001_11101001_10101010_1;
      patterns[49644] = 25'b11000001_11101010_10101011_1;
      patterns[49645] = 25'b11000001_11101011_10101100_1;
      patterns[49646] = 25'b11000001_11101100_10101101_1;
      patterns[49647] = 25'b11000001_11101101_10101110_1;
      patterns[49648] = 25'b11000001_11101110_10101111_1;
      patterns[49649] = 25'b11000001_11101111_10110000_1;
      patterns[49650] = 25'b11000001_11110000_10110001_1;
      patterns[49651] = 25'b11000001_11110001_10110010_1;
      patterns[49652] = 25'b11000001_11110010_10110011_1;
      patterns[49653] = 25'b11000001_11110011_10110100_1;
      patterns[49654] = 25'b11000001_11110100_10110101_1;
      patterns[49655] = 25'b11000001_11110101_10110110_1;
      patterns[49656] = 25'b11000001_11110110_10110111_1;
      patterns[49657] = 25'b11000001_11110111_10111000_1;
      patterns[49658] = 25'b11000001_11111000_10111001_1;
      patterns[49659] = 25'b11000001_11111001_10111010_1;
      patterns[49660] = 25'b11000001_11111010_10111011_1;
      patterns[49661] = 25'b11000001_11111011_10111100_1;
      patterns[49662] = 25'b11000001_11111100_10111101_1;
      patterns[49663] = 25'b11000001_11111101_10111110_1;
      patterns[49664] = 25'b11000001_11111110_10111111_1;
      patterns[49665] = 25'b11000001_11111111_11000000_1;
      patterns[49666] = 25'b11000010_00000000_11000010_0;
      patterns[49667] = 25'b11000010_00000001_11000011_0;
      patterns[49668] = 25'b11000010_00000010_11000100_0;
      patterns[49669] = 25'b11000010_00000011_11000101_0;
      patterns[49670] = 25'b11000010_00000100_11000110_0;
      patterns[49671] = 25'b11000010_00000101_11000111_0;
      patterns[49672] = 25'b11000010_00000110_11001000_0;
      patterns[49673] = 25'b11000010_00000111_11001001_0;
      patterns[49674] = 25'b11000010_00001000_11001010_0;
      patterns[49675] = 25'b11000010_00001001_11001011_0;
      patterns[49676] = 25'b11000010_00001010_11001100_0;
      patterns[49677] = 25'b11000010_00001011_11001101_0;
      patterns[49678] = 25'b11000010_00001100_11001110_0;
      patterns[49679] = 25'b11000010_00001101_11001111_0;
      patterns[49680] = 25'b11000010_00001110_11010000_0;
      patterns[49681] = 25'b11000010_00001111_11010001_0;
      patterns[49682] = 25'b11000010_00010000_11010010_0;
      patterns[49683] = 25'b11000010_00010001_11010011_0;
      patterns[49684] = 25'b11000010_00010010_11010100_0;
      patterns[49685] = 25'b11000010_00010011_11010101_0;
      patterns[49686] = 25'b11000010_00010100_11010110_0;
      patterns[49687] = 25'b11000010_00010101_11010111_0;
      patterns[49688] = 25'b11000010_00010110_11011000_0;
      patterns[49689] = 25'b11000010_00010111_11011001_0;
      patterns[49690] = 25'b11000010_00011000_11011010_0;
      patterns[49691] = 25'b11000010_00011001_11011011_0;
      patterns[49692] = 25'b11000010_00011010_11011100_0;
      patterns[49693] = 25'b11000010_00011011_11011101_0;
      patterns[49694] = 25'b11000010_00011100_11011110_0;
      patterns[49695] = 25'b11000010_00011101_11011111_0;
      patterns[49696] = 25'b11000010_00011110_11100000_0;
      patterns[49697] = 25'b11000010_00011111_11100001_0;
      patterns[49698] = 25'b11000010_00100000_11100010_0;
      patterns[49699] = 25'b11000010_00100001_11100011_0;
      patterns[49700] = 25'b11000010_00100010_11100100_0;
      patterns[49701] = 25'b11000010_00100011_11100101_0;
      patterns[49702] = 25'b11000010_00100100_11100110_0;
      patterns[49703] = 25'b11000010_00100101_11100111_0;
      patterns[49704] = 25'b11000010_00100110_11101000_0;
      patterns[49705] = 25'b11000010_00100111_11101001_0;
      patterns[49706] = 25'b11000010_00101000_11101010_0;
      patterns[49707] = 25'b11000010_00101001_11101011_0;
      patterns[49708] = 25'b11000010_00101010_11101100_0;
      patterns[49709] = 25'b11000010_00101011_11101101_0;
      patterns[49710] = 25'b11000010_00101100_11101110_0;
      patterns[49711] = 25'b11000010_00101101_11101111_0;
      patterns[49712] = 25'b11000010_00101110_11110000_0;
      patterns[49713] = 25'b11000010_00101111_11110001_0;
      patterns[49714] = 25'b11000010_00110000_11110010_0;
      patterns[49715] = 25'b11000010_00110001_11110011_0;
      patterns[49716] = 25'b11000010_00110010_11110100_0;
      patterns[49717] = 25'b11000010_00110011_11110101_0;
      patterns[49718] = 25'b11000010_00110100_11110110_0;
      patterns[49719] = 25'b11000010_00110101_11110111_0;
      patterns[49720] = 25'b11000010_00110110_11111000_0;
      patterns[49721] = 25'b11000010_00110111_11111001_0;
      patterns[49722] = 25'b11000010_00111000_11111010_0;
      patterns[49723] = 25'b11000010_00111001_11111011_0;
      patterns[49724] = 25'b11000010_00111010_11111100_0;
      patterns[49725] = 25'b11000010_00111011_11111101_0;
      patterns[49726] = 25'b11000010_00111100_11111110_0;
      patterns[49727] = 25'b11000010_00111101_11111111_0;
      patterns[49728] = 25'b11000010_00111110_00000000_1;
      patterns[49729] = 25'b11000010_00111111_00000001_1;
      patterns[49730] = 25'b11000010_01000000_00000010_1;
      patterns[49731] = 25'b11000010_01000001_00000011_1;
      patterns[49732] = 25'b11000010_01000010_00000100_1;
      patterns[49733] = 25'b11000010_01000011_00000101_1;
      patterns[49734] = 25'b11000010_01000100_00000110_1;
      patterns[49735] = 25'b11000010_01000101_00000111_1;
      patterns[49736] = 25'b11000010_01000110_00001000_1;
      patterns[49737] = 25'b11000010_01000111_00001001_1;
      patterns[49738] = 25'b11000010_01001000_00001010_1;
      patterns[49739] = 25'b11000010_01001001_00001011_1;
      patterns[49740] = 25'b11000010_01001010_00001100_1;
      patterns[49741] = 25'b11000010_01001011_00001101_1;
      patterns[49742] = 25'b11000010_01001100_00001110_1;
      patterns[49743] = 25'b11000010_01001101_00001111_1;
      patterns[49744] = 25'b11000010_01001110_00010000_1;
      patterns[49745] = 25'b11000010_01001111_00010001_1;
      patterns[49746] = 25'b11000010_01010000_00010010_1;
      patterns[49747] = 25'b11000010_01010001_00010011_1;
      patterns[49748] = 25'b11000010_01010010_00010100_1;
      patterns[49749] = 25'b11000010_01010011_00010101_1;
      patterns[49750] = 25'b11000010_01010100_00010110_1;
      patterns[49751] = 25'b11000010_01010101_00010111_1;
      patterns[49752] = 25'b11000010_01010110_00011000_1;
      patterns[49753] = 25'b11000010_01010111_00011001_1;
      patterns[49754] = 25'b11000010_01011000_00011010_1;
      patterns[49755] = 25'b11000010_01011001_00011011_1;
      patterns[49756] = 25'b11000010_01011010_00011100_1;
      patterns[49757] = 25'b11000010_01011011_00011101_1;
      patterns[49758] = 25'b11000010_01011100_00011110_1;
      patterns[49759] = 25'b11000010_01011101_00011111_1;
      patterns[49760] = 25'b11000010_01011110_00100000_1;
      patterns[49761] = 25'b11000010_01011111_00100001_1;
      patterns[49762] = 25'b11000010_01100000_00100010_1;
      patterns[49763] = 25'b11000010_01100001_00100011_1;
      patterns[49764] = 25'b11000010_01100010_00100100_1;
      patterns[49765] = 25'b11000010_01100011_00100101_1;
      patterns[49766] = 25'b11000010_01100100_00100110_1;
      patterns[49767] = 25'b11000010_01100101_00100111_1;
      patterns[49768] = 25'b11000010_01100110_00101000_1;
      patterns[49769] = 25'b11000010_01100111_00101001_1;
      patterns[49770] = 25'b11000010_01101000_00101010_1;
      patterns[49771] = 25'b11000010_01101001_00101011_1;
      patterns[49772] = 25'b11000010_01101010_00101100_1;
      patterns[49773] = 25'b11000010_01101011_00101101_1;
      patterns[49774] = 25'b11000010_01101100_00101110_1;
      patterns[49775] = 25'b11000010_01101101_00101111_1;
      patterns[49776] = 25'b11000010_01101110_00110000_1;
      patterns[49777] = 25'b11000010_01101111_00110001_1;
      patterns[49778] = 25'b11000010_01110000_00110010_1;
      patterns[49779] = 25'b11000010_01110001_00110011_1;
      patterns[49780] = 25'b11000010_01110010_00110100_1;
      patterns[49781] = 25'b11000010_01110011_00110101_1;
      patterns[49782] = 25'b11000010_01110100_00110110_1;
      patterns[49783] = 25'b11000010_01110101_00110111_1;
      patterns[49784] = 25'b11000010_01110110_00111000_1;
      patterns[49785] = 25'b11000010_01110111_00111001_1;
      patterns[49786] = 25'b11000010_01111000_00111010_1;
      patterns[49787] = 25'b11000010_01111001_00111011_1;
      patterns[49788] = 25'b11000010_01111010_00111100_1;
      patterns[49789] = 25'b11000010_01111011_00111101_1;
      patterns[49790] = 25'b11000010_01111100_00111110_1;
      patterns[49791] = 25'b11000010_01111101_00111111_1;
      patterns[49792] = 25'b11000010_01111110_01000000_1;
      patterns[49793] = 25'b11000010_01111111_01000001_1;
      patterns[49794] = 25'b11000010_10000000_01000010_1;
      patterns[49795] = 25'b11000010_10000001_01000011_1;
      patterns[49796] = 25'b11000010_10000010_01000100_1;
      patterns[49797] = 25'b11000010_10000011_01000101_1;
      patterns[49798] = 25'b11000010_10000100_01000110_1;
      patterns[49799] = 25'b11000010_10000101_01000111_1;
      patterns[49800] = 25'b11000010_10000110_01001000_1;
      patterns[49801] = 25'b11000010_10000111_01001001_1;
      patterns[49802] = 25'b11000010_10001000_01001010_1;
      patterns[49803] = 25'b11000010_10001001_01001011_1;
      patterns[49804] = 25'b11000010_10001010_01001100_1;
      patterns[49805] = 25'b11000010_10001011_01001101_1;
      patterns[49806] = 25'b11000010_10001100_01001110_1;
      patterns[49807] = 25'b11000010_10001101_01001111_1;
      patterns[49808] = 25'b11000010_10001110_01010000_1;
      patterns[49809] = 25'b11000010_10001111_01010001_1;
      patterns[49810] = 25'b11000010_10010000_01010010_1;
      patterns[49811] = 25'b11000010_10010001_01010011_1;
      patterns[49812] = 25'b11000010_10010010_01010100_1;
      patterns[49813] = 25'b11000010_10010011_01010101_1;
      patterns[49814] = 25'b11000010_10010100_01010110_1;
      patterns[49815] = 25'b11000010_10010101_01010111_1;
      patterns[49816] = 25'b11000010_10010110_01011000_1;
      patterns[49817] = 25'b11000010_10010111_01011001_1;
      patterns[49818] = 25'b11000010_10011000_01011010_1;
      patterns[49819] = 25'b11000010_10011001_01011011_1;
      patterns[49820] = 25'b11000010_10011010_01011100_1;
      patterns[49821] = 25'b11000010_10011011_01011101_1;
      patterns[49822] = 25'b11000010_10011100_01011110_1;
      patterns[49823] = 25'b11000010_10011101_01011111_1;
      patterns[49824] = 25'b11000010_10011110_01100000_1;
      patterns[49825] = 25'b11000010_10011111_01100001_1;
      patterns[49826] = 25'b11000010_10100000_01100010_1;
      patterns[49827] = 25'b11000010_10100001_01100011_1;
      patterns[49828] = 25'b11000010_10100010_01100100_1;
      patterns[49829] = 25'b11000010_10100011_01100101_1;
      patterns[49830] = 25'b11000010_10100100_01100110_1;
      patterns[49831] = 25'b11000010_10100101_01100111_1;
      patterns[49832] = 25'b11000010_10100110_01101000_1;
      patterns[49833] = 25'b11000010_10100111_01101001_1;
      patterns[49834] = 25'b11000010_10101000_01101010_1;
      patterns[49835] = 25'b11000010_10101001_01101011_1;
      patterns[49836] = 25'b11000010_10101010_01101100_1;
      patterns[49837] = 25'b11000010_10101011_01101101_1;
      patterns[49838] = 25'b11000010_10101100_01101110_1;
      patterns[49839] = 25'b11000010_10101101_01101111_1;
      patterns[49840] = 25'b11000010_10101110_01110000_1;
      patterns[49841] = 25'b11000010_10101111_01110001_1;
      patterns[49842] = 25'b11000010_10110000_01110010_1;
      patterns[49843] = 25'b11000010_10110001_01110011_1;
      patterns[49844] = 25'b11000010_10110010_01110100_1;
      patterns[49845] = 25'b11000010_10110011_01110101_1;
      patterns[49846] = 25'b11000010_10110100_01110110_1;
      patterns[49847] = 25'b11000010_10110101_01110111_1;
      patterns[49848] = 25'b11000010_10110110_01111000_1;
      patterns[49849] = 25'b11000010_10110111_01111001_1;
      patterns[49850] = 25'b11000010_10111000_01111010_1;
      patterns[49851] = 25'b11000010_10111001_01111011_1;
      patterns[49852] = 25'b11000010_10111010_01111100_1;
      patterns[49853] = 25'b11000010_10111011_01111101_1;
      patterns[49854] = 25'b11000010_10111100_01111110_1;
      patterns[49855] = 25'b11000010_10111101_01111111_1;
      patterns[49856] = 25'b11000010_10111110_10000000_1;
      patterns[49857] = 25'b11000010_10111111_10000001_1;
      patterns[49858] = 25'b11000010_11000000_10000010_1;
      patterns[49859] = 25'b11000010_11000001_10000011_1;
      patterns[49860] = 25'b11000010_11000010_10000100_1;
      patterns[49861] = 25'b11000010_11000011_10000101_1;
      patterns[49862] = 25'b11000010_11000100_10000110_1;
      patterns[49863] = 25'b11000010_11000101_10000111_1;
      patterns[49864] = 25'b11000010_11000110_10001000_1;
      patterns[49865] = 25'b11000010_11000111_10001001_1;
      patterns[49866] = 25'b11000010_11001000_10001010_1;
      patterns[49867] = 25'b11000010_11001001_10001011_1;
      patterns[49868] = 25'b11000010_11001010_10001100_1;
      patterns[49869] = 25'b11000010_11001011_10001101_1;
      patterns[49870] = 25'b11000010_11001100_10001110_1;
      patterns[49871] = 25'b11000010_11001101_10001111_1;
      patterns[49872] = 25'b11000010_11001110_10010000_1;
      patterns[49873] = 25'b11000010_11001111_10010001_1;
      patterns[49874] = 25'b11000010_11010000_10010010_1;
      patterns[49875] = 25'b11000010_11010001_10010011_1;
      patterns[49876] = 25'b11000010_11010010_10010100_1;
      patterns[49877] = 25'b11000010_11010011_10010101_1;
      patterns[49878] = 25'b11000010_11010100_10010110_1;
      patterns[49879] = 25'b11000010_11010101_10010111_1;
      patterns[49880] = 25'b11000010_11010110_10011000_1;
      patterns[49881] = 25'b11000010_11010111_10011001_1;
      patterns[49882] = 25'b11000010_11011000_10011010_1;
      patterns[49883] = 25'b11000010_11011001_10011011_1;
      patterns[49884] = 25'b11000010_11011010_10011100_1;
      patterns[49885] = 25'b11000010_11011011_10011101_1;
      patterns[49886] = 25'b11000010_11011100_10011110_1;
      patterns[49887] = 25'b11000010_11011101_10011111_1;
      patterns[49888] = 25'b11000010_11011110_10100000_1;
      patterns[49889] = 25'b11000010_11011111_10100001_1;
      patterns[49890] = 25'b11000010_11100000_10100010_1;
      patterns[49891] = 25'b11000010_11100001_10100011_1;
      patterns[49892] = 25'b11000010_11100010_10100100_1;
      patterns[49893] = 25'b11000010_11100011_10100101_1;
      patterns[49894] = 25'b11000010_11100100_10100110_1;
      patterns[49895] = 25'b11000010_11100101_10100111_1;
      patterns[49896] = 25'b11000010_11100110_10101000_1;
      patterns[49897] = 25'b11000010_11100111_10101001_1;
      patterns[49898] = 25'b11000010_11101000_10101010_1;
      patterns[49899] = 25'b11000010_11101001_10101011_1;
      patterns[49900] = 25'b11000010_11101010_10101100_1;
      patterns[49901] = 25'b11000010_11101011_10101101_1;
      patterns[49902] = 25'b11000010_11101100_10101110_1;
      patterns[49903] = 25'b11000010_11101101_10101111_1;
      patterns[49904] = 25'b11000010_11101110_10110000_1;
      patterns[49905] = 25'b11000010_11101111_10110001_1;
      patterns[49906] = 25'b11000010_11110000_10110010_1;
      patterns[49907] = 25'b11000010_11110001_10110011_1;
      patterns[49908] = 25'b11000010_11110010_10110100_1;
      patterns[49909] = 25'b11000010_11110011_10110101_1;
      patterns[49910] = 25'b11000010_11110100_10110110_1;
      patterns[49911] = 25'b11000010_11110101_10110111_1;
      patterns[49912] = 25'b11000010_11110110_10111000_1;
      patterns[49913] = 25'b11000010_11110111_10111001_1;
      patterns[49914] = 25'b11000010_11111000_10111010_1;
      patterns[49915] = 25'b11000010_11111001_10111011_1;
      patterns[49916] = 25'b11000010_11111010_10111100_1;
      patterns[49917] = 25'b11000010_11111011_10111101_1;
      patterns[49918] = 25'b11000010_11111100_10111110_1;
      patterns[49919] = 25'b11000010_11111101_10111111_1;
      patterns[49920] = 25'b11000010_11111110_11000000_1;
      patterns[49921] = 25'b11000010_11111111_11000001_1;
      patterns[49922] = 25'b11000011_00000000_11000011_0;
      patterns[49923] = 25'b11000011_00000001_11000100_0;
      patterns[49924] = 25'b11000011_00000010_11000101_0;
      patterns[49925] = 25'b11000011_00000011_11000110_0;
      patterns[49926] = 25'b11000011_00000100_11000111_0;
      patterns[49927] = 25'b11000011_00000101_11001000_0;
      patterns[49928] = 25'b11000011_00000110_11001001_0;
      patterns[49929] = 25'b11000011_00000111_11001010_0;
      patterns[49930] = 25'b11000011_00001000_11001011_0;
      patterns[49931] = 25'b11000011_00001001_11001100_0;
      patterns[49932] = 25'b11000011_00001010_11001101_0;
      patterns[49933] = 25'b11000011_00001011_11001110_0;
      patterns[49934] = 25'b11000011_00001100_11001111_0;
      patterns[49935] = 25'b11000011_00001101_11010000_0;
      patterns[49936] = 25'b11000011_00001110_11010001_0;
      patterns[49937] = 25'b11000011_00001111_11010010_0;
      patterns[49938] = 25'b11000011_00010000_11010011_0;
      patterns[49939] = 25'b11000011_00010001_11010100_0;
      patterns[49940] = 25'b11000011_00010010_11010101_0;
      patterns[49941] = 25'b11000011_00010011_11010110_0;
      patterns[49942] = 25'b11000011_00010100_11010111_0;
      patterns[49943] = 25'b11000011_00010101_11011000_0;
      patterns[49944] = 25'b11000011_00010110_11011001_0;
      patterns[49945] = 25'b11000011_00010111_11011010_0;
      patterns[49946] = 25'b11000011_00011000_11011011_0;
      patterns[49947] = 25'b11000011_00011001_11011100_0;
      patterns[49948] = 25'b11000011_00011010_11011101_0;
      patterns[49949] = 25'b11000011_00011011_11011110_0;
      patterns[49950] = 25'b11000011_00011100_11011111_0;
      patterns[49951] = 25'b11000011_00011101_11100000_0;
      patterns[49952] = 25'b11000011_00011110_11100001_0;
      patterns[49953] = 25'b11000011_00011111_11100010_0;
      patterns[49954] = 25'b11000011_00100000_11100011_0;
      patterns[49955] = 25'b11000011_00100001_11100100_0;
      patterns[49956] = 25'b11000011_00100010_11100101_0;
      patterns[49957] = 25'b11000011_00100011_11100110_0;
      patterns[49958] = 25'b11000011_00100100_11100111_0;
      patterns[49959] = 25'b11000011_00100101_11101000_0;
      patterns[49960] = 25'b11000011_00100110_11101001_0;
      patterns[49961] = 25'b11000011_00100111_11101010_0;
      patterns[49962] = 25'b11000011_00101000_11101011_0;
      patterns[49963] = 25'b11000011_00101001_11101100_0;
      patterns[49964] = 25'b11000011_00101010_11101101_0;
      patterns[49965] = 25'b11000011_00101011_11101110_0;
      patterns[49966] = 25'b11000011_00101100_11101111_0;
      patterns[49967] = 25'b11000011_00101101_11110000_0;
      patterns[49968] = 25'b11000011_00101110_11110001_0;
      patterns[49969] = 25'b11000011_00101111_11110010_0;
      patterns[49970] = 25'b11000011_00110000_11110011_0;
      patterns[49971] = 25'b11000011_00110001_11110100_0;
      patterns[49972] = 25'b11000011_00110010_11110101_0;
      patterns[49973] = 25'b11000011_00110011_11110110_0;
      patterns[49974] = 25'b11000011_00110100_11110111_0;
      patterns[49975] = 25'b11000011_00110101_11111000_0;
      patterns[49976] = 25'b11000011_00110110_11111001_0;
      patterns[49977] = 25'b11000011_00110111_11111010_0;
      patterns[49978] = 25'b11000011_00111000_11111011_0;
      patterns[49979] = 25'b11000011_00111001_11111100_0;
      patterns[49980] = 25'b11000011_00111010_11111101_0;
      patterns[49981] = 25'b11000011_00111011_11111110_0;
      patterns[49982] = 25'b11000011_00111100_11111111_0;
      patterns[49983] = 25'b11000011_00111101_00000000_1;
      patterns[49984] = 25'b11000011_00111110_00000001_1;
      patterns[49985] = 25'b11000011_00111111_00000010_1;
      patterns[49986] = 25'b11000011_01000000_00000011_1;
      patterns[49987] = 25'b11000011_01000001_00000100_1;
      patterns[49988] = 25'b11000011_01000010_00000101_1;
      patterns[49989] = 25'b11000011_01000011_00000110_1;
      patterns[49990] = 25'b11000011_01000100_00000111_1;
      patterns[49991] = 25'b11000011_01000101_00001000_1;
      patterns[49992] = 25'b11000011_01000110_00001001_1;
      patterns[49993] = 25'b11000011_01000111_00001010_1;
      patterns[49994] = 25'b11000011_01001000_00001011_1;
      patterns[49995] = 25'b11000011_01001001_00001100_1;
      patterns[49996] = 25'b11000011_01001010_00001101_1;
      patterns[49997] = 25'b11000011_01001011_00001110_1;
      patterns[49998] = 25'b11000011_01001100_00001111_1;
      patterns[49999] = 25'b11000011_01001101_00010000_1;
      patterns[50000] = 25'b11000011_01001110_00010001_1;
      patterns[50001] = 25'b11000011_01001111_00010010_1;
      patterns[50002] = 25'b11000011_01010000_00010011_1;
      patterns[50003] = 25'b11000011_01010001_00010100_1;
      patterns[50004] = 25'b11000011_01010010_00010101_1;
      patterns[50005] = 25'b11000011_01010011_00010110_1;
      patterns[50006] = 25'b11000011_01010100_00010111_1;
      patterns[50007] = 25'b11000011_01010101_00011000_1;
      patterns[50008] = 25'b11000011_01010110_00011001_1;
      patterns[50009] = 25'b11000011_01010111_00011010_1;
      patterns[50010] = 25'b11000011_01011000_00011011_1;
      patterns[50011] = 25'b11000011_01011001_00011100_1;
      patterns[50012] = 25'b11000011_01011010_00011101_1;
      patterns[50013] = 25'b11000011_01011011_00011110_1;
      patterns[50014] = 25'b11000011_01011100_00011111_1;
      patterns[50015] = 25'b11000011_01011101_00100000_1;
      patterns[50016] = 25'b11000011_01011110_00100001_1;
      patterns[50017] = 25'b11000011_01011111_00100010_1;
      patterns[50018] = 25'b11000011_01100000_00100011_1;
      patterns[50019] = 25'b11000011_01100001_00100100_1;
      patterns[50020] = 25'b11000011_01100010_00100101_1;
      patterns[50021] = 25'b11000011_01100011_00100110_1;
      patterns[50022] = 25'b11000011_01100100_00100111_1;
      patterns[50023] = 25'b11000011_01100101_00101000_1;
      patterns[50024] = 25'b11000011_01100110_00101001_1;
      patterns[50025] = 25'b11000011_01100111_00101010_1;
      patterns[50026] = 25'b11000011_01101000_00101011_1;
      patterns[50027] = 25'b11000011_01101001_00101100_1;
      patterns[50028] = 25'b11000011_01101010_00101101_1;
      patterns[50029] = 25'b11000011_01101011_00101110_1;
      patterns[50030] = 25'b11000011_01101100_00101111_1;
      patterns[50031] = 25'b11000011_01101101_00110000_1;
      patterns[50032] = 25'b11000011_01101110_00110001_1;
      patterns[50033] = 25'b11000011_01101111_00110010_1;
      patterns[50034] = 25'b11000011_01110000_00110011_1;
      patterns[50035] = 25'b11000011_01110001_00110100_1;
      patterns[50036] = 25'b11000011_01110010_00110101_1;
      patterns[50037] = 25'b11000011_01110011_00110110_1;
      patterns[50038] = 25'b11000011_01110100_00110111_1;
      patterns[50039] = 25'b11000011_01110101_00111000_1;
      patterns[50040] = 25'b11000011_01110110_00111001_1;
      patterns[50041] = 25'b11000011_01110111_00111010_1;
      patterns[50042] = 25'b11000011_01111000_00111011_1;
      patterns[50043] = 25'b11000011_01111001_00111100_1;
      patterns[50044] = 25'b11000011_01111010_00111101_1;
      patterns[50045] = 25'b11000011_01111011_00111110_1;
      patterns[50046] = 25'b11000011_01111100_00111111_1;
      patterns[50047] = 25'b11000011_01111101_01000000_1;
      patterns[50048] = 25'b11000011_01111110_01000001_1;
      patterns[50049] = 25'b11000011_01111111_01000010_1;
      patterns[50050] = 25'b11000011_10000000_01000011_1;
      patterns[50051] = 25'b11000011_10000001_01000100_1;
      patterns[50052] = 25'b11000011_10000010_01000101_1;
      patterns[50053] = 25'b11000011_10000011_01000110_1;
      patterns[50054] = 25'b11000011_10000100_01000111_1;
      patterns[50055] = 25'b11000011_10000101_01001000_1;
      patterns[50056] = 25'b11000011_10000110_01001001_1;
      patterns[50057] = 25'b11000011_10000111_01001010_1;
      patterns[50058] = 25'b11000011_10001000_01001011_1;
      patterns[50059] = 25'b11000011_10001001_01001100_1;
      patterns[50060] = 25'b11000011_10001010_01001101_1;
      patterns[50061] = 25'b11000011_10001011_01001110_1;
      patterns[50062] = 25'b11000011_10001100_01001111_1;
      patterns[50063] = 25'b11000011_10001101_01010000_1;
      patterns[50064] = 25'b11000011_10001110_01010001_1;
      patterns[50065] = 25'b11000011_10001111_01010010_1;
      patterns[50066] = 25'b11000011_10010000_01010011_1;
      patterns[50067] = 25'b11000011_10010001_01010100_1;
      patterns[50068] = 25'b11000011_10010010_01010101_1;
      patterns[50069] = 25'b11000011_10010011_01010110_1;
      patterns[50070] = 25'b11000011_10010100_01010111_1;
      patterns[50071] = 25'b11000011_10010101_01011000_1;
      patterns[50072] = 25'b11000011_10010110_01011001_1;
      patterns[50073] = 25'b11000011_10010111_01011010_1;
      patterns[50074] = 25'b11000011_10011000_01011011_1;
      patterns[50075] = 25'b11000011_10011001_01011100_1;
      patterns[50076] = 25'b11000011_10011010_01011101_1;
      patterns[50077] = 25'b11000011_10011011_01011110_1;
      patterns[50078] = 25'b11000011_10011100_01011111_1;
      patterns[50079] = 25'b11000011_10011101_01100000_1;
      patterns[50080] = 25'b11000011_10011110_01100001_1;
      patterns[50081] = 25'b11000011_10011111_01100010_1;
      patterns[50082] = 25'b11000011_10100000_01100011_1;
      patterns[50083] = 25'b11000011_10100001_01100100_1;
      patterns[50084] = 25'b11000011_10100010_01100101_1;
      patterns[50085] = 25'b11000011_10100011_01100110_1;
      patterns[50086] = 25'b11000011_10100100_01100111_1;
      patterns[50087] = 25'b11000011_10100101_01101000_1;
      patterns[50088] = 25'b11000011_10100110_01101001_1;
      patterns[50089] = 25'b11000011_10100111_01101010_1;
      patterns[50090] = 25'b11000011_10101000_01101011_1;
      patterns[50091] = 25'b11000011_10101001_01101100_1;
      patterns[50092] = 25'b11000011_10101010_01101101_1;
      patterns[50093] = 25'b11000011_10101011_01101110_1;
      patterns[50094] = 25'b11000011_10101100_01101111_1;
      patterns[50095] = 25'b11000011_10101101_01110000_1;
      patterns[50096] = 25'b11000011_10101110_01110001_1;
      patterns[50097] = 25'b11000011_10101111_01110010_1;
      patterns[50098] = 25'b11000011_10110000_01110011_1;
      patterns[50099] = 25'b11000011_10110001_01110100_1;
      patterns[50100] = 25'b11000011_10110010_01110101_1;
      patterns[50101] = 25'b11000011_10110011_01110110_1;
      patterns[50102] = 25'b11000011_10110100_01110111_1;
      patterns[50103] = 25'b11000011_10110101_01111000_1;
      patterns[50104] = 25'b11000011_10110110_01111001_1;
      patterns[50105] = 25'b11000011_10110111_01111010_1;
      patterns[50106] = 25'b11000011_10111000_01111011_1;
      patterns[50107] = 25'b11000011_10111001_01111100_1;
      patterns[50108] = 25'b11000011_10111010_01111101_1;
      patterns[50109] = 25'b11000011_10111011_01111110_1;
      patterns[50110] = 25'b11000011_10111100_01111111_1;
      patterns[50111] = 25'b11000011_10111101_10000000_1;
      patterns[50112] = 25'b11000011_10111110_10000001_1;
      patterns[50113] = 25'b11000011_10111111_10000010_1;
      patterns[50114] = 25'b11000011_11000000_10000011_1;
      patterns[50115] = 25'b11000011_11000001_10000100_1;
      patterns[50116] = 25'b11000011_11000010_10000101_1;
      patterns[50117] = 25'b11000011_11000011_10000110_1;
      patterns[50118] = 25'b11000011_11000100_10000111_1;
      patterns[50119] = 25'b11000011_11000101_10001000_1;
      patterns[50120] = 25'b11000011_11000110_10001001_1;
      patterns[50121] = 25'b11000011_11000111_10001010_1;
      patterns[50122] = 25'b11000011_11001000_10001011_1;
      patterns[50123] = 25'b11000011_11001001_10001100_1;
      patterns[50124] = 25'b11000011_11001010_10001101_1;
      patterns[50125] = 25'b11000011_11001011_10001110_1;
      patterns[50126] = 25'b11000011_11001100_10001111_1;
      patterns[50127] = 25'b11000011_11001101_10010000_1;
      patterns[50128] = 25'b11000011_11001110_10010001_1;
      patterns[50129] = 25'b11000011_11001111_10010010_1;
      patterns[50130] = 25'b11000011_11010000_10010011_1;
      patterns[50131] = 25'b11000011_11010001_10010100_1;
      patterns[50132] = 25'b11000011_11010010_10010101_1;
      patterns[50133] = 25'b11000011_11010011_10010110_1;
      patterns[50134] = 25'b11000011_11010100_10010111_1;
      patterns[50135] = 25'b11000011_11010101_10011000_1;
      patterns[50136] = 25'b11000011_11010110_10011001_1;
      patterns[50137] = 25'b11000011_11010111_10011010_1;
      patterns[50138] = 25'b11000011_11011000_10011011_1;
      patterns[50139] = 25'b11000011_11011001_10011100_1;
      patterns[50140] = 25'b11000011_11011010_10011101_1;
      patterns[50141] = 25'b11000011_11011011_10011110_1;
      patterns[50142] = 25'b11000011_11011100_10011111_1;
      patterns[50143] = 25'b11000011_11011101_10100000_1;
      patterns[50144] = 25'b11000011_11011110_10100001_1;
      patterns[50145] = 25'b11000011_11011111_10100010_1;
      patterns[50146] = 25'b11000011_11100000_10100011_1;
      patterns[50147] = 25'b11000011_11100001_10100100_1;
      patterns[50148] = 25'b11000011_11100010_10100101_1;
      patterns[50149] = 25'b11000011_11100011_10100110_1;
      patterns[50150] = 25'b11000011_11100100_10100111_1;
      patterns[50151] = 25'b11000011_11100101_10101000_1;
      patterns[50152] = 25'b11000011_11100110_10101001_1;
      patterns[50153] = 25'b11000011_11100111_10101010_1;
      patterns[50154] = 25'b11000011_11101000_10101011_1;
      patterns[50155] = 25'b11000011_11101001_10101100_1;
      patterns[50156] = 25'b11000011_11101010_10101101_1;
      patterns[50157] = 25'b11000011_11101011_10101110_1;
      patterns[50158] = 25'b11000011_11101100_10101111_1;
      patterns[50159] = 25'b11000011_11101101_10110000_1;
      patterns[50160] = 25'b11000011_11101110_10110001_1;
      patterns[50161] = 25'b11000011_11101111_10110010_1;
      patterns[50162] = 25'b11000011_11110000_10110011_1;
      patterns[50163] = 25'b11000011_11110001_10110100_1;
      patterns[50164] = 25'b11000011_11110010_10110101_1;
      patterns[50165] = 25'b11000011_11110011_10110110_1;
      patterns[50166] = 25'b11000011_11110100_10110111_1;
      patterns[50167] = 25'b11000011_11110101_10111000_1;
      patterns[50168] = 25'b11000011_11110110_10111001_1;
      patterns[50169] = 25'b11000011_11110111_10111010_1;
      patterns[50170] = 25'b11000011_11111000_10111011_1;
      patterns[50171] = 25'b11000011_11111001_10111100_1;
      patterns[50172] = 25'b11000011_11111010_10111101_1;
      patterns[50173] = 25'b11000011_11111011_10111110_1;
      patterns[50174] = 25'b11000011_11111100_10111111_1;
      patterns[50175] = 25'b11000011_11111101_11000000_1;
      patterns[50176] = 25'b11000011_11111110_11000001_1;
      patterns[50177] = 25'b11000011_11111111_11000010_1;
      patterns[50178] = 25'b11000100_00000000_11000100_0;
      patterns[50179] = 25'b11000100_00000001_11000101_0;
      patterns[50180] = 25'b11000100_00000010_11000110_0;
      patterns[50181] = 25'b11000100_00000011_11000111_0;
      patterns[50182] = 25'b11000100_00000100_11001000_0;
      patterns[50183] = 25'b11000100_00000101_11001001_0;
      patterns[50184] = 25'b11000100_00000110_11001010_0;
      patterns[50185] = 25'b11000100_00000111_11001011_0;
      patterns[50186] = 25'b11000100_00001000_11001100_0;
      patterns[50187] = 25'b11000100_00001001_11001101_0;
      patterns[50188] = 25'b11000100_00001010_11001110_0;
      patterns[50189] = 25'b11000100_00001011_11001111_0;
      patterns[50190] = 25'b11000100_00001100_11010000_0;
      patterns[50191] = 25'b11000100_00001101_11010001_0;
      patterns[50192] = 25'b11000100_00001110_11010010_0;
      patterns[50193] = 25'b11000100_00001111_11010011_0;
      patterns[50194] = 25'b11000100_00010000_11010100_0;
      patterns[50195] = 25'b11000100_00010001_11010101_0;
      patterns[50196] = 25'b11000100_00010010_11010110_0;
      patterns[50197] = 25'b11000100_00010011_11010111_0;
      patterns[50198] = 25'b11000100_00010100_11011000_0;
      patterns[50199] = 25'b11000100_00010101_11011001_0;
      patterns[50200] = 25'b11000100_00010110_11011010_0;
      patterns[50201] = 25'b11000100_00010111_11011011_0;
      patterns[50202] = 25'b11000100_00011000_11011100_0;
      patterns[50203] = 25'b11000100_00011001_11011101_0;
      patterns[50204] = 25'b11000100_00011010_11011110_0;
      patterns[50205] = 25'b11000100_00011011_11011111_0;
      patterns[50206] = 25'b11000100_00011100_11100000_0;
      patterns[50207] = 25'b11000100_00011101_11100001_0;
      patterns[50208] = 25'b11000100_00011110_11100010_0;
      patterns[50209] = 25'b11000100_00011111_11100011_0;
      patterns[50210] = 25'b11000100_00100000_11100100_0;
      patterns[50211] = 25'b11000100_00100001_11100101_0;
      patterns[50212] = 25'b11000100_00100010_11100110_0;
      patterns[50213] = 25'b11000100_00100011_11100111_0;
      patterns[50214] = 25'b11000100_00100100_11101000_0;
      patterns[50215] = 25'b11000100_00100101_11101001_0;
      patterns[50216] = 25'b11000100_00100110_11101010_0;
      patterns[50217] = 25'b11000100_00100111_11101011_0;
      patterns[50218] = 25'b11000100_00101000_11101100_0;
      patterns[50219] = 25'b11000100_00101001_11101101_0;
      patterns[50220] = 25'b11000100_00101010_11101110_0;
      patterns[50221] = 25'b11000100_00101011_11101111_0;
      patterns[50222] = 25'b11000100_00101100_11110000_0;
      patterns[50223] = 25'b11000100_00101101_11110001_0;
      patterns[50224] = 25'b11000100_00101110_11110010_0;
      patterns[50225] = 25'b11000100_00101111_11110011_0;
      patterns[50226] = 25'b11000100_00110000_11110100_0;
      patterns[50227] = 25'b11000100_00110001_11110101_0;
      patterns[50228] = 25'b11000100_00110010_11110110_0;
      patterns[50229] = 25'b11000100_00110011_11110111_0;
      patterns[50230] = 25'b11000100_00110100_11111000_0;
      patterns[50231] = 25'b11000100_00110101_11111001_0;
      patterns[50232] = 25'b11000100_00110110_11111010_0;
      patterns[50233] = 25'b11000100_00110111_11111011_0;
      patterns[50234] = 25'b11000100_00111000_11111100_0;
      patterns[50235] = 25'b11000100_00111001_11111101_0;
      patterns[50236] = 25'b11000100_00111010_11111110_0;
      patterns[50237] = 25'b11000100_00111011_11111111_0;
      patterns[50238] = 25'b11000100_00111100_00000000_1;
      patterns[50239] = 25'b11000100_00111101_00000001_1;
      patterns[50240] = 25'b11000100_00111110_00000010_1;
      patterns[50241] = 25'b11000100_00111111_00000011_1;
      patterns[50242] = 25'b11000100_01000000_00000100_1;
      patterns[50243] = 25'b11000100_01000001_00000101_1;
      patterns[50244] = 25'b11000100_01000010_00000110_1;
      patterns[50245] = 25'b11000100_01000011_00000111_1;
      patterns[50246] = 25'b11000100_01000100_00001000_1;
      patterns[50247] = 25'b11000100_01000101_00001001_1;
      patterns[50248] = 25'b11000100_01000110_00001010_1;
      patterns[50249] = 25'b11000100_01000111_00001011_1;
      patterns[50250] = 25'b11000100_01001000_00001100_1;
      patterns[50251] = 25'b11000100_01001001_00001101_1;
      patterns[50252] = 25'b11000100_01001010_00001110_1;
      patterns[50253] = 25'b11000100_01001011_00001111_1;
      patterns[50254] = 25'b11000100_01001100_00010000_1;
      patterns[50255] = 25'b11000100_01001101_00010001_1;
      patterns[50256] = 25'b11000100_01001110_00010010_1;
      patterns[50257] = 25'b11000100_01001111_00010011_1;
      patterns[50258] = 25'b11000100_01010000_00010100_1;
      patterns[50259] = 25'b11000100_01010001_00010101_1;
      patterns[50260] = 25'b11000100_01010010_00010110_1;
      patterns[50261] = 25'b11000100_01010011_00010111_1;
      patterns[50262] = 25'b11000100_01010100_00011000_1;
      patterns[50263] = 25'b11000100_01010101_00011001_1;
      patterns[50264] = 25'b11000100_01010110_00011010_1;
      patterns[50265] = 25'b11000100_01010111_00011011_1;
      patterns[50266] = 25'b11000100_01011000_00011100_1;
      patterns[50267] = 25'b11000100_01011001_00011101_1;
      patterns[50268] = 25'b11000100_01011010_00011110_1;
      patterns[50269] = 25'b11000100_01011011_00011111_1;
      patterns[50270] = 25'b11000100_01011100_00100000_1;
      patterns[50271] = 25'b11000100_01011101_00100001_1;
      patterns[50272] = 25'b11000100_01011110_00100010_1;
      patterns[50273] = 25'b11000100_01011111_00100011_1;
      patterns[50274] = 25'b11000100_01100000_00100100_1;
      patterns[50275] = 25'b11000100_01100001_00100101_1;
      patterns[50276] = 25'b11000100_01100010_00100110_1;
      patterns[50277] = 25'b11000100_01100011_00100111_1;
      patterns[50278] = 25'b11000100_01100100_00101000_1;
      patterns[50279] = 25'b11000100_01100101_00101001_1;
      patterns[50280] = 25'b11000100_01100110_00101010_1;
      patterns[50281] = 25'b11000100_01100111_00101011_1;
      patterns[50282] = 25'b11000100_01101000_00101100_1;
      patterns[50283] = 25'b11000100_01101001_00101101_1;
      patterns[50284] = 25'b11000100_01101010_00101110_1;
      patterns[50285] = 25'b11000100_01101011_00101111_1;
      patterns[50286] = 25'b11000100_01101100_00110000_1;
      patterns[50287] = 25'b11000100_01101101_00110001_1;
      patterns[50288] = 25'b11000100_01101110_00110010_1;
      patterns[50289] = 25'b11000100_01101111_00110011_1;
      patterns[50290] = 25'b11000100_01110000_00110100_1;
      patterns[50291] = 25'b11000100_01110001_00110101_1;
      patterns[50292] = 25'b11000100_01110010_00110110_1;
      patterns[50293] = 25'b11000100_01110011_00110111_1;
      patterns[50294] = 25'b11000100_01110100_00111000_1;
      patterns[50295] = 25'b11000100_01110101_00111001_1;
      patterns[50296] = 25'b11000100_01110110_00111010_1;
      patterns[50297] = 25'b11000100_01110111_00111011_1;
      patterns[50298] = 25'b11000100_01111000_00111100_1;
      patterns[50299] = 25'b11000100_01111001_00111101_1;
      patterns[50300] = 25'b11000100_01111010_00111110_1;
      patterns[50301] = 25'b11000100_01111011_00111111_1;
      patterns[50302] = 25'b11000100_01111100_01000000_1;
      patterns[50303] = 25'b11000100_01111101_01000001_1;
      patterns[50304] = 25'b11000100_01111110_01000010_1;
      patterns[50305] = 25'b11000100_01111111_01000011_1;
      patterns[50306] = 25'b11000100_10000000_01000100_1;
      patterns[50307] = 25'b11000100_10000001_01000101_1;
      patterns[50308] = 25'b11000100_10000010_01000110_1;
      patterns[50309] = 25'b11000100_10000011_01000111_1;
      patterns[50310] = 25'b11000100_10000100_01001000_1;
      patterns[50311] = 25'b11000100_10000101_01001001_1;
      patterns[50312] = 25'b11000100_10000110_01001010_1;
      patterns[50313] = 25'b11000100_10000111_01001011_1;
      patterns[50314] = 25'b11000100_10001000_01001100_1;
      patterns[50315] = 25'b11000100_10001001_01001101_1;
      patterns[50316] = 25'b11000100_10001010_01001110_1;
      patterns[50317] = 25'b11000100_10001011_01001111_1;
      patterns[50318] = 25'b11000100_10001100_01010000_1;
      patterns[50319] = 25'b11000100_10001101_01010001_1;
      patterns[50320] = 25'b11000100_10001110_01010010_1;
      patterns[50321] = 25'b11000100_10001111_01010011_1;
      patterns[50322] = 25'b11000100_10010000_01010100_1;
      patterns[50323] = 25'b11000100_10010001_01010101_1;
      patterns[50324] = 25'b11000100_10010010_01010110_1;
      patterns[50325] = 25'b11000100_10010011_01010111_1;
      patterns[50326] = 25'b11000100_10010100_01011000_1;
      patterns[50327] = 25'b11000100_10010101_01011001_1;
      patterns[50328] = 25'b11000100_10010110_01011010_1;
      patterns[50329] = 25'b11000100_10010111_01011011_1;
      patterns[50330] = 25'b11000100_10011000_01011100_1;
      patterns[50331] = 25'b11000100_10011001_01011101_1;
      patterns[50332] = 25'b11000100_10011010_01011110_1;
      patterns[50333] = 25'b11000100_10011011_01011111_1;
      patterns[50334] = 25'b11000100_10011100_01100000_1;
      patterns[50335] = 25'b11000100_10011101_01100001_1;
      patterns[50336] = 25'b11000100_10011110_01100010_1;
      patterns[50337] = 25'b11000100_10011111_01100011_1;
      patterns[50338] = 25'b11000100_10100000_01100100_1;
      patterns[50339] = 25'b11000100_10100001_01100101_1;
      patterns[50340] = 25'b11000100_10100010_01100110_1;
      patterns[50341] = 25'b11000100_10100011_01100111_1;
      patterns[50342] = 25'b11000100_10100100_01101000_1;
      patterns[50343] = 25'b11000100_10100101_01101001_1;
      patterns[50344] = 25'b11000100_10100110_01101010_1;
      patterns[50345] = 25'b11000100_10100111_01101011_1;
      patterns[50346] = 25'b11000100_10101000_01101100_1;
      patterns[50347] = 25'b11000100_10101001_01101101_1;
      patterns[50348] = 25'b11000100_10101010_01101110_1;
      patterns[50349] = 25'b11000100_10101011_01101111_1;
      patterns[50350] = 25'b11000100_10101100_01110000_1;
      patterns[50351] = 25'b11000100_10101101_01110001_1;
      patterns[50352] = 25'b11000100_10101110_01110010_1;
      patterns[50353] = 25'b11000100_10101111_01110011_1;
      patterns[50354] = 25'b11000100_10110000_01110100_1;
      patterns[50355] = 25'b11000100_10110001_01110101_1;
      patterns[50356] = 25'b11000100_10110010_01110110_1;
      patterns[50357] = 25'b11000100_10110011_01110111_1;
      patterns[50358] = 25'b11000100_10110100_01111000_1;
      patterns[50359] = 25'b11000100_10110101_01111001_1;
      patterns[50360] = 25'b11000100_10110110_01111010_1;
      patterns[50361] = 25'b11000100_10110111_01111011_1;
      patterns[50362] = 25'b11000100_10111000_01111100_1;
      patterns[50363] = 25'b11000100_10111001_01111101_1;
      patterns[50364] = 25'b11000100_10111010_01111110_1;
      patterns[50365] = 25'b11000100_10111011_01111111_1;
      patterns[50366] = 25'b11000100_10111100_10000000_1;
      patterns[50367] = 25'b11000100_10111101_10000001_1;
      patterns[50368] = 25'b11000100_10111110_10000010_1;
      patterns[50369] = 25'b11000100_10111111_10000011_1;
      patterns[50370] = 25'b11000100_11000000_10000100_1;
      patterns[50371] = 25'b11000100_11000001_10000101_1;
      patterns[50372] = 25'b11000100_11000010_10000110_1;
      patterns[50373] = 25'b11000100_11000011_10000111_1;
      patterns[50374] = 25'b11000100_11000100_10001000_1;
      patterns[50375] = 25'b11000100_11000101_10001001_1;
      patterns[50376] = 25'b11000100_11000110_10001010_1;
      patterns[50377] = 25'b11000100_11000111_10001011_1;
      patterns[50378] = 25'b11000100_11001000_10001100_1;
      patterns[50379] = 25'b11000100_11001001_10001101_1;
      patterns[50380] = 25'b11000100_11001010_10001110_1;
      patterns[50381] = 25'b11000100_11001011_10001111_1;
      patterns[50382] = 25'b11000100_11001100_10010000_1;
      patterns[50383] = 25'b11000100_11001101_10010001_1;
      patterns[50384] = 25'b11000100_11001110_10010010_1;
      patterns[50385] = 25'b11000100_11001111_10010011_1;
      patterns[50386] = 25'b11000100_11010000_10010100_1;
      patterns[50387] = 25'b11000100_11010001_10010101_1;
      patterns[50388] = 25'b11000100_11010010_10010110_1;
      patterns[50389] = 25'b11000100_11010011_10010111_1;
      patterns[50390] = 25'b11000100_11010100_10011000_1;
      patterns[50391] = 25'b11000100_11010101_10011001_1;
      patterns[50392] = 25'b11000100_11010110_10011010_1;
      patterns[50393] = 25'b11000100_11010111_10011011_1;
      patterns[50394] = 25'b11000100_11011000_10011100_1;
      patterns[50395] = 25'b11000100_11011001_10011101_1;
      patterns[50396] = 25'b11000100_11011010_10011110_1;
      patterns[50397] = 25'b11000100_11011011_10011111_1;
      patterns[50398] = 25'b11000100_11011100_10100000_1;
      patterns[50399] = 25'b11000100_11011101_10100001_1;
      patterns[50400] = 25'b11000100_11011110_10100010_1;
      patterns[50401] = 25'b11000100_11011111_10100011_1;
      patterns[50402] = 25'b11000100_11100000_10100100_1;
      patterns[50403] = 25'b11000100_11100001_10100101_1;
      patterns[50404] = 25'b11000100_11100010_10100110_1;
      patterns[50405] = 25'b11000100_11100011_10100111_1;
      patterns[50406] = 25'b11000100_11100100_10101000_1;
      patterns[50407] = 25'b11000100_11100101_10101001_1;
      patterns[50408] = 25'b11000100_11100110_10101010_1;
      patterns[50409] = 25'b11000100_11100111_10101011_1;
      patterns[50410] = 25'b11000100_11101000_10101100_1;
      patterns[50411] = 25'b11000100_11101001_10101101_1;
      patterns[50412] = 25'b11000100_11101010_10101110_1;
      patterns[50413] = 25'b11000100_11101011_10101111_1;
      patterns[50414] = 25'b11000100_11101100_10110000_1;
      patterns[50415] = 25'b11000100_11101101_10110001_1;
      patterns[50416] = 25'b11000100_11101110_10110010_1;
      patterns[50417] = 25'b11000100_11101111_10110011_1;
      patterns[50418] = 25'b11000100_11110000_10110100_1;
      patterns[50419] = 25'b11000100_11110001_10110101_1;
      patterns[50420] = 25'b11000100_11110010_10110110_1;
      patterns[50421] = 25'b11000100_11110011_10110111_1;
      patterns[50422] = 25'b11000100_11110100_10111000_1;
      patterns[50423] = 25'b11000100_11110101_10111001_1;
      patterns[50424] = 25'b11000100_11110110_10111010_1;
      patterns[50425] = 25'b11000100_11110111_10111011_1;
      patterns[50426] = 25'b11000100_11111000_10111100_1;
      patterns[50427] = 25'b11000100_11111001_10111101_1;
      patterns[50428] = 25'b11000100_11111010_10111110_1;
      patterns[50429] = 25'b11000100_11111011_10111111_1;
      patterns[50430] = 25'b11000100_11111100_11000000_1;
      patterns[50431] = 25'b11000100_11111101_11000001_1;
      patterns[50432] = 25'b11000100_11111110_11000010_1;
      patterns[50433] = 25'b11000100_11111111_11000011_1;
      patterns[50434] = 25'b11000101_00000000_11000101_0;
      patterns[50435] = 25'b11000101_00000001_11000110_0;
      patterns[50436] = 25'b11000101_00000010_11000111_0;
      patterns[50437] = 25'b11000101_00000011_11001000_0;
      patterns[50438] = 25'b11000101_00000100_11001001_0;
      patterns[50439] = 25'b11000101_00000101_11001010_0;
      patterns[50440] = 25'b11000101_00000110_11001011_0;
      patterns[50441] = 25'b11000101_00000111_11001100_0;
      patterns[50442] = 25'b11000101_00001000_11001101_0;
      patterns[50443] = 25'b11000101_00001001_11001110_0;
      patterns[50444] = 25'b11000101_00001010_11001111_0;
      patterns[50445] = 25'b11000101_00001011_11010000_0;
      patterns[50446] = 25'b11000101_00001100_11010001_0;
      patterns[50447] = 25'b11000101_00001101_11010010_0;
      patterns[50448] = 25'b11000101_00001110_11010011_0;
      patterns[50449] = 25'b11000101_00001111_11010100_0;
      patterns[50450] = 25'b11000101_00010000_11010101_0;
      patterns[50451] = 25'b11000101_00010001_11010110_0;
      patterns[50452] = 25'b11000101_00010010_11010111_0;
      patterns[50453] = 25'b11000101_00010011_11011000_0;
      patterns[50454] = 25'b11000101_00010100_11011001_0;
      patterns[50455] = 25'b11000101_00010101_11011010_0;
      patterns[50456] = 25'b11000101_00010110_11011011_0;
      patterns[50457] = 25'b11000101_00010111_11011100_0;
      patterns[50458] = 25'b11000101_00011000_11011101_0;
      patterns[50459] = 25'b11000101_00011001_11011110_0;
      patterns[50460] = 25'b11000101_00011010_11011111_0;
      patterns[50461] = 25'b11000101_00011011_11100000_0;
      patterns[50462] = 25'b11000101_00011100_11100001_0;
      patterns[50463] = 25'b11000101_00011101_11100010_0;
      patterns[50464] = 25'b11000101_00011110_11100011_0;
      patterns[50465] = 25'b11000101_00011111_11100100_0;
      patterns[50466] = 25'b11000101_00100000_11100101_0;
      patterns[50467] = 25'b11000101_00100001_11100110_0;
      patterns[50468] = 25'b11000101_00100010_11100111_0;
      patterns[50469] = 25'b11000101_00100011_11101000_0;
      patterns[50470] = 25'b11000101_00100100_11101001_0;
      patterns[50471] = 25'b11000101_00100101_11101010_0;
      patterns[50472] = 25'b11000101_00100110_11101011_0;
      patterns[50473] = 25'b11000101_00100111_11101100_0;
      patterns[50474] = 25'b11000101_00101000_11101101_0;
      patterns[50475] = 25'b11000101_00101001_11101110_0;
      patterns[50476] = 25'b11000101_00101010_11101111_0;
      patterns[50477] = 25'b11000101_00101011_11110000_0;
      patterns[50478] = 25'b11000101_00101100_11110001_0;
      patterns[50479] = 25'b11000101_00101101_11110010_0;
      patterns[50480] = 25'b11000101_00101110_11110011_0;
      patterns[50481] = 25'b11000101_00101111_11110100_0;
      patterns[50482] = 25'b11000101_00110000_11110101_0;
      patterns[50483] = 25'b11000101_00110001_11110110_0;
      patterns[50484] = 25'b11000101_00110010_11110111_0;
      patterns[50485] = 25'b11000101_00110011_11111000_0;
      patterns[50486] = 25'b11000101_00110100_11111001_0;
      patterns[50487] = 25'b11000101_00110101_11111010_0;
      patterns[50488] = 25'b11000101_00110110_11111011_0;
      patterns[50489] = 25'b11000101_00110111_11111100_0;
      patterns[50490] = 25'b11000101_00111000_11111101_0;
      patterns[50491] = 25'b11000101_00111001_11111110_0;
      patterns[50492] = 25'b11000101_00111010_11111111_0;
      patterns[50493] = 25'b11000101_00111011_00000000_1;
      patterns[50494] = 25'b11000101_00111100_00000001_1;
      patterns[50495] = 25'b11000101_00111101_00000010_1;
      patterns[50496] = 25'b11000101_00111110_00000011_1;
      patterns[50497] = 25'b11000101_00111111_00000100_1;
      patterns[50498] = 25'b11000101_01000000_00000101_1;
      patterns[50499] = 25'b11000101_01000001_00000110_1;
      patterns[50500] = 25'b11000101_01000010_00000111_1;
      patterns[50501] = 25'b11000101_01000011_00001000_1;
      patterns[50502] = 25'b11000101_01000100_00001001_1;
      patterns[50503] = 25'b11000101_01000101_00001010_1;
      patterns[50504] = 25'b11000101_01000110_00001011_1;
      patterns[50505] = 25'b11000101_01000111_00001100_1;
      patterns[50506] = 25'b11000101_01001000_00001101_1;
      patterns[50507] = 25'b11000101_01001001_00001110_1;
      patterns[50508] = 25'b11000101_01001010_00001111_1;
      patterns[50509] = 25'b11000101_01001011_00010000_1;
      patterns[50510] = 25'b11000101_01001100_00010001_1;
      patterns[50511] = 25'b11000101_01001101_00010010_1;
      patterns[50512] = 25'b11000101_01001110_00010011_1;
      patterns[50513] = 25'b11000101_01001111_00010100_1;
      patterns[50514] = 25'b11000101_01010000_00010101_1;
      patterns[50515] = 25'b11000101_01010001_00010110_1;
      patterns[50516] = 25'b11000101_01010010_00010111_1;
      patterns[50517] = 25'b11000101_01010011_00011000_1;
      patterns[50518] = 25'b11000101_01010100_00011001_1;
      patterns[50519] = 25'b11000101_01010101_00011010_1;
      patterns[50520] = 25'b11000101_01010110_00011011_1;
      patterns[50521] = 25'b11000101_01010111_00011100_1;
      patterns[50522] = 25'b11000101_01011000_00011101_1;
      patterns[50523] = 25'b11000101_01011001_00011110_1;
      patterns[50524] = 25'b11000101_01011010_00011111_1;
      patterns[50525] = 25'b11000101_01011011_00100000_1;
      patterns[50526] = 25'b11000101_01011100_00100001_1;
      patterns[50527] = 25'b11000101_01011101_00100010_1;
      patterns[50528] = 25'b11000101_01011110_00100011_1;
      patterns[50529] = 25'b11000101_01011111_00100100_1;
      patterns[50530] = 25'b11000101_01100000_00100101_1;
      patterns[50531] = 25'b11000101_01100001_00100110_1;
      patterns[50532] = 25'b11000101_01100010_00100111_1;
      patterns[50533] = 25'b11000101_01100011_00101000_1;
      patterns[50534] = 25'b11000101_01100100_00101001_1;
      patterns[50535] = 25'b11000101_01100101_00101010_1;
      patterns[50536] = 25'b11000101_01100110_00101011_1;
      patterns[50537] = 25'b11000101_01100111_00101100_1;
      patterns[50538] = 25'b11000101_01101000_00101101_1;
      patterns[50539] = 25'b11000101_01101001_00101110_1;
      patterns[50540] = 25'b11000101_01101010_00101111_1;
      patterns[50541] = 25'b11000101_01101011_00110000_1;
      patterns[50542] = 25'b11000101_01101100_00110001_1;
      patterns[50543] = 25'b11000101_01101101_00110010_1;
      patterns[50544] = 25'b11000101_01101110_00110011_1;
      patterns[50545] = 25'b11000101_01101111_00110100_1;
      patterns[50546] = 25'b11000101_01110000_00110101_1;
      patterns[50547] = 25'b11000101_01110001_00110110_1;
      patterns[50548] = 25'b11000101_01110010_00110111_1;
      patterns[50549] = 25'b11000101_01110011_00111000_1;
      patterns[50550] = 25'b11000101_01110100_00111001_1;
      patterns[50551] = 25'b11000101_01110101_00111010_1;
      patterns[50552] = 25'b11000101_01110110_00111011_1;
      patterns[50553] = 25'b11000101_01110111_00111100_1;
      patterns[50554] = 25'b11000101_01111000_00111101_1;
      patterns[50555] = 25'b11000101_01111001_00111110_1;
      patterns[50556] = 25'b11000101_01111010_00111111_1;
      patterns[50557] = 25'b11000101_01111011_01000000_1;
      patterns[50558] = 25'b11000101_01111100_01000001_1;
      patterns[50559] = 25'b11000101_01111101_01000010_1;
      patterns[50560] = 25'b11000101_01111110_01000011_1;
      patterns[50561] = 25'b11000101_01111111_01000100_1;
      patterns[50562] = 25'b11000101_10000000_01000101_1;
      patterns[50563] = 25'b11000101_10000001_01000110_1;
      patterns[50564] = 25'b11000101_10000010_01000111_1;
      patterns[50565] = 25'b11000101_10000011_01001000_1;
      patterns[50566] = 25'b11000101_10000100_01001001_1;
      patterns[50567] = 25'b11000101_10000101_01001010_1;
      patterns[50568] = 25'b11000101_10000110_01001011_1;
      patterns[50569] = 25'b11000101_10000111_01001100_1;
      patterns[50570] = 25'b11000101_10001000_01001101_1;
      patterns[50571] = 25'b11000101_10001001_01001110_1;
      patterns[50572] = 25'b11000101_10001010_01001111_1;
      patterns[50573] = 25'b11000101_10001011_01010000_1;
      patterns[50574] = 25'b11000101_10001100_01010001_1;
      patterns[50575] = 25'b11000101_10001101_01010010_1;
      patterns[50576] = 25'b11000101_10001110_01010011_1;
      patterns[50577] = 25'b11000101_10001111_01010100_1;
      patterns[50578] = 25'b11000101_10010000_01010101_1;
      patterns[50579] = 25'b11000101_10010001_01010110_1;
      patterns[50580] = 25'b11000101_10010010_01010111_1;
      patterns[50581] = 25'b11000101_10010011_01011000_1;
      patterns[50582] = 25'b11000101_10010100_01011001_1;
      patterns[50583] = 25'b11000101_10010101_01011010_1;
      patterns[50584] = 25'b11000101_10010110_01011011_1;
      patterns[50585] = 25'b11000101_10010111_01011100_1;
      patterns[50586] = 25'b11000101_10011000_01011101_1;
      patterns[50587] = 25'b11000101_10011001_01011110_1;
      patterns[50588] = 25'b11000101_10011010_01011111_1;
      patterns[50589] = 25'b11000101_10011011_01100000_1;
      patterns[50590] = 25'b11000101_10011100_01100001_1;
      patterns[50591] = 25'b11000101_10011101_01100010_1;
      patterns[50592] = 25'b11000101_10011110_01100011_1;
      patterns[50593] = 25'b11000101_10011111_01100100_1;
      patterns[50594] = 25'b11000101_10100000_01100101_1;
      patterns[50595] = 25'b11000101_10100001_01100110_1;
      patterns[50596] = 25'b11000101_10100010_01100111_1;
      patterns[50597] = 25'b11000101_10100011_01101000_1;
      patterns[50598] = 25'b11000101_10100100_01101001_1;
      patterns[50599] = 25'b11000101_10100101_01101010_1;
      patterns[50600] = 25'b11000101_10100110_01101011_1;
      patterns[50601] = 25'b11000101_10100111_01101100_1;
      patterns[50602] = 25'b11000101_10101000_01101101_1;
      patterns[50603] = 25'b11000101_10101001_01101110_1;
      patterns[50604] = 25'b11000101_10101010_01101111_1;
      patterns[50605] = 25'b11000101_10101011_01110000_1;
      patterns[50606] = 25'b11000101_10101100_01110001_1;
      patterns[50607] = 25'b11000101_10101101_01110010_1;
      patterns[50608] = 25'b11000101_10101110_01110011_1;
      patterns[50609] = 25'b11000101_10101111_01110100_1;
      patterns[50610] = 25'b11000101_10110000_01110101_1;
      patterns[50611] = 25'b11000101_10110001_01110110_1;
      patterns[50612] = 25'b11000101_10110010_01110111_1;
      patterns[50613] = 25'b11000101_10110011_01111000_1;
      patterns[50614] = 25'b11000101_10110100_01111001_1;
      patterns[50615] = 25'b11000101_10110101_01111010_1;
      patterns[50616] = 25'b11000101_10110110_01111011_1;
      patterns[50617] = 25'b11000101_10110111_01111100_1;
      patterns[50618] = 25'b11000101_10111000_01111101_1;
      patterns[50619] = 25'b11000101_10111001_01111110_1;
      patterns[50620] = 25'b11000101_10111010_01111111_1;
      patterns[50621] = 25'b11000101_10111011_10000000_1;
      patterns[50622] = 25'b11000101_10111100_10000001_1;
      patterns[50623] = 25'b11000101_10111101_10000010_1;
      patterns[50624] = 25'b11000101_10111110_10000011_1;
      patterns[50625] = 25'b11000101_10111111_10000100_1;
      patterns[50626] = 25'b11000101_11000000_10000101_1;
      patterns[50627] = 25'b11000101_11000001_10000110_1;
      patterns[50628] = 25'b11000101_11000010_10000111_1;
      patterns[50629] = 25'b11000101_11000011_10001000_1;
      patterns[50630] = 25'b11000101_11000100_10001001_1;
      patterns[50631] = 25'b11000101_11000101_10001010_1;
      patterns[50632] = 25'b11000101_11000110_10001011_1;
      patterns[50633] = 25'b11000101_11000111_10001100_1;
      patterns[50634] = 25'b11000101_11001000_10001101_1;
      patterns[50635] = 25'b11000101_11001001_10001110_1;
      patterns[50636] = 25'b11000101_11001010_10001111_1;
      patterns[50637] = 25'b11000101_11001011_10010000_1;
      patterns[50638] = 25'b11000101_11001100_10010001_1;
      patterns[50639] = 25'b11000101_11001101_10010010_1;
      patterns[50640] = 25'b11000101_11001110_10010011_1;
      patterns[50641] = 25'b11000101_11001111_10010100_1;
      patterns[50642] = 25'b11000101_11010000_10010101_1;
      patterns[50643] = 25'b11000101_11010001_10010110_1;
      patterns[50644] = 25'b11000101_11010010_10010111_1;
      patterns[50645] = 25'b11000101_11010011_10011000_1;
      patterns[50646] = 25'b11000101_11010100_10011001_1;
      patterns[50647] = 25'b11000101_11010101_10011010_1;
      patterns[50648] = 25'b11000101_11010110_10011011_1;
      patterns[50649] = 25'b11000101_11010111_10011100_1;
      patterns[50650] = 25'b11000101_11011000_10011101_1;
      patterns[50651] = 25'b11000101_11011001_10011110_1;
      patterns[50652] = 25'b11000101_11011010_10011111_1;
      patterns[50653] = 25'b11000101_11011011_10100000_1;
      patterns[50654] = 25'b11000101_11011100_10100001_1;
      patterns[50655] = 25'b11000101_11011101_10100010_1;
      patterns[50656] = 25'b11000101_11011110_10100011_1;
      patterns[50657] = 25'b11000101_11011111_10100100_1;
      patterns[50658] = 25'b11000101_11100000_10100101_1;
      patterns[50659] = 25'b11000101_11100001_10100110_1;
      patterns[50660] = 25'b11000101_11100010_10100111_1;
      patterns[50661] = 25'b11000101_11100011_10101000_1;
      patterns[50662] = 25'b11000101_11100100_10101001_1;
      patterns[50663] = 25'b11000101_11100101_10101010_1;
      patterns[50664] = 25'b11000101_11100110_10101011_1;
      patterns[50665] = 25'b11000101_11100111_10101100_1;
      patterns[50666] = 25'b11000101_11101000_10101101_1;
      patterns[50667] = 25'b11000101_11101001_10101110_1;
      patterns[50668] = 25'b11000101_11101010_10101111_1;
      patterns[50669] = 25'b11000101_11101011_10110000_1;
      patterns[50670] = 25'b11000101_11101100_10110001_1;
      patterns[50671] = 25'b11000101_11101101_10110010_1;
      patterns[50672] = 25'b11000101_11101110_10110011_1;
      patterns[50673] = 25'b11000101_11101111_10110100_1;
      patterns[50674] = 25'b11000101_11110000_10110101_1;
      patterns[50675] = 25'b11000101_11110001_10110110_1;
      patterns[50676] = 25'b11000101_11110010_10110111_1;
      patterns[50677] = 25'b11000101_11110011_10111000_1;
      patterns[50678] = 25'b11000101_11110100_10111001_1;
      patterns[50679] = 25'b11000101_11110101_10111010_1;
      patterns[50680] = 25'b11000101_11110110_10111011_1;
      patterns[50681] = 25'b11000101_11110111_10111100_1;
      patterns[50682] = 25'b11000101_11111000_10111101_1;
      patterns[50683] = 25'b11000101_11111001_10111110_1;
      patterns[50684] = 25'b11000101_11111010_10111111_1;
      patterns[50685] = 25'b11000101_11111011_11000000_1;
      patterns[50686] = 25'b11000101_11111100_11000001_1;
      patterns[50687] = 25'b11000101_11111101_11000010_1;
      patterns[50688] = 25'b11000101_11111110_11000011_1;
      patterns[50689] = 25'b11000101_11111111_11000100_1;
      patterns[50690] = 25'b11000110_00000000_11000110_0;
      patterns[50691] = 25'b11000110_00000001_11000111_0;
      patterns[50692] = 25'b11000110_00000010_11001000_0;
      patterns[50693] = 25'b11000110_00000011_11001001_0;
      patterns[50694] = 25'b11000110_00000100_11001010_0;
      patterns[50695] = 25'b11000110_00000101_11001011_0;
      patterns[50696] = 25'b11000110_00000110_11001100_0;
      patterns[50697] = 25'b11000110_00000111_11001101_0;
      patterns[50698] = 25'b11000110_00001000_11001110_0;
      patterns[50699] = 25'b11000110_00001001_11001111_0;
      patterns[50700] = 25'b11000110_00001010_11010000_0;
      patterns[50701] = 25'b11000110_00001011_11010001_0;
      patterns[50702] = 25'b11000110_00001100_11010010_0;
      patterns[50703] = 25'b11000110_00001101_11010011_0;
      patterns[50704] = 25'b11000110_00001110_11010100_0;
      patterns[50705] = 25'b11000110_00001111_11010101_0;
      patterns[50706] = 25'b11000110_00010000_11010110_0;
      patterns[50707] = 25'b11000110_00010001_11010111_0;
      patterns[50708] = 25'b11000110_00010010_11011000_0;
      patterns[50709] = 25'b11000110_00010011_11011001_0;
      patterns[50710] = 25'b11000110_00010100_11011010_0;
      patterns[50711] = 25'b11000110_00010101_11011011_0;
      patterns[50712] = 25'b11000110_00010110_11011100_0;
      patterns[50713] = 25'b11000110_00010111_11011101_0;
      patterns[50714] = 25'b11000110_00011000_11011110_0;
      patterns[50715] = 25'b11000110_00011001_11011111_0;
      patterns[50716] = 25'b11000110_00011010_11100000_0;
      patterns[50717] = 25'b11000110_00011011_11100001_0;
      patterns[50718] = 25'b11000110_00011100_11100010_0;
      patterns[50719] = 25'b11000110_00011101_11100011_0;
      patterns[50720] = 25'b11000110_00011110_11100100_0;
      patterns[50721] = 25'b11000110_00011111_11100101_0;
      patterns[50722] = 25'b11000110_00100000_11100110_0;
      patterns[50723] = 25'b11000110_00100001_11100111_0;
      patterns[50724] = 25'b11000110_00100010_11101000_0;
      patterns[50725] = 25'b11000110_00100011_11101001_0;
      patterns[50726] = 25'b11000110_00100100_11101010_0;
      patterns[50727] = 25'b11000110_00100101_11101011_0;
      patterns[50728] = 25'b11000110_00100110_11101100_0;
      patterns[50729] = 25'b11000110_00100111_11101101_0;
      patterns[50730] = 25'b11000110_00101000_11101110_0;
      patterns[50731] = 25'b11000110_00101001_11101111_0;
      patterns[50732] = 25'b11000110_00101010_11110000_0;
      patterns[50733] = 25'b11000110_00101011_11110001_0;
      patterns[50734] = 25'b11000110_00101100_11110010_0;
      patterns[50735] = 25'b11000110_00101101_11110011_0;
      patterns[50736] = 25'b11000110_00101110_11110100_0;
      patterns[50737] = 25'b11000110_00101111_11110101_0;
      patterns[50738] = 25'b11000110_00110000_11110110_0;
      patterns[50739] = 25'b11000110_00110001_11110111_0;
      patterns[50740] = 25'b11000110_00110010_11111000_0;
      patterns[50741] = 25'b11000110_00110011_11111001_0;
      patterns[50742] = 25'b11000110_00110100_11111010_0;
      patterns[50743] = 25'b11000110_00110101_11111011_0;
      patterns[50744] = 25'b11000110_00110110_11111100_0;
      patterns[50745] = 25'b11000110_00110111_11111101_0;
      patterns[50746] = 25'b11000110_00111000_11111110_0;
      patterns[50747] = 25'b11000110_00111001_11111111_0;
      patterns[50748] = 25'b11000110_00111010_00000000_1;
      patterns[50749] = 25'b11000110_00111011_00000001_1;
      patterns[50750] = 25'b11000110_00111100_00000010_1;
      patterns[50751] = 25'b11000110_00111101_00000011_1;
      patterns[50752] = 25'b11000110_00111110_00000100_1;
      patterns[50753] = 25'b11000110_00111111_00000101_1;
      patterns[50754] = 25'b11000110_01000000_00000110_1;
      patterns[50755] = 25'b11000110_01000001_00000111_1;
      patterns[50756] = 25'b11000110_01000010_00001000_1;
      patterns[50757] = 25'b11000110_01000011_00001001_1;
      patterns[50758] = 25'b11000110_01000100_00001010_1;
      patterns[50759] = 25'b11000110_01000101_00001011_1;
      patterns[50760] = 25'b11000110_01000110_00001100_1;
      patterns[50761] = 25'b11000110_01000111_00001101_1;
      patterns[50762] = 25'b11000110_01001000_00001110_1;
      patterns[50763] = 25'b11000110_01001001_00001111_1;
      patterns[50764] = 25'b11000110_01001010_00010000_1;
      patterns[50765] = 25'b11000110_01001011_00010001_1;
      patterns[50766] = 25'b11000110_01001100_00010010_1;
      patterns[50767] = 25'b11000110_01001101_00010011_1;
      patterns[50768] = 25'b11000110_01001110_00010100_1;
      patterns[50769] = 25'b11000110_01001111_00010101_1;
      patterns[50770] = 25'b11000110_01010000_00010110_1;
      patterns[50771] = 25'b11000110_01010001_00010111_1;
      patterns[50772] = 25'b11000110_01010010_00011000_1;
      patterns[50773] = 25'b11000110_01010011_00011001_1;
      patterns[50774] = 25'b11000110_01010100_00011010_1;
      patterns[50775] = 25'b11000110_01010101_00011011_1;
      patterns[50776] = 25'b11000110_01010110_00011100_1;
      patterns[50777] = 25'b11000110_01010111_00011101_1;
      patterns[50778] = 25'b11000110_01011000_00011110_1;
      patterns[50779] = 25'b11000110_01011001_00011111_1;
      patterns[50780] = 25'b11000110_01011010_00100000_1;
      patterns[50781] = 25'b11000110_01011011_00100001_1;
      patterns[50782] = 25'b11000110_01011100_00100010_1;
      patterns[50783] = 25'b11000110_01011101_00100011_1;
      patterns[50784] = 25'b11000110_01011110_00100100_1;
      patterns[50785] = 25'b11000110_01011111_00100101_1;
      patterns[50786] = 25'b11000110_01100000_00100110_1;
      patterns[50787] = 25'b11000110_01100001_00100111_1;
      patterns[50788] = 25'b11000110_01100010_00101000_1;
      patterns[50789] = 25'b11000110_01100011_00101001_1;
      patterns[50790] = 25'b11000110_01100100_00101010_1;
      patterns[50791] = 25'b11000110_01100101_00101011_1;
      patterns[50792] = 25'b11000110_01100110_00101100_1;
      patterns[50793] = 25'b11000110_01100111_00101101_1;
      patterns[50794] = 25'b11000110_01101000_00101110_1;
      patterns[50795] = 25'b11000110_01101001_00101111_1;
      patterns[50796] = 25'b11000110_01101010_00110000_1;
      patterns[50797] = 25'b11000110_01101011_00110001_1;
      patterns[50798] = 25'b11000110_01101100_00110010_1;
      patterns[50799] = 25'b11000110_01101101_00110011_1;
      patterns[50800] = 25'b11000110_01101110_00110100_1;
      patterns[50801] = 25'b11000110_01101111_00110101_1;
      patterns[50802] = 25'b11000110_01110000_00110110_1;
      patterns[50803] = 25'b11000110_01110001_00110111_1;
      patterns[50804] = 25'b11000110_01110010_00111000_1;
      patterns[50805] = 25'b11000110_01110011_00111001_1;
      patterns[50806] = 25'b11000110_01110100_00111010_1;
      patterns[50807] = 25'b11000110_01110101_00111011_1;
      patterns[50808] = 25'b11000110_01110110_00111100_1;
      patterns[50809] = 25'b11000110_01110111_00111101_1;
      patterns[50810] = 25'b11000110_01111000_00111110_1;
      patterns[50811] = 25'b11000110_01111001_00111111_1;
      patterns[50812] = 25'b11000110_01111010_01000000_1;
      patterns[50813] = 25'b11000110_01111011_01000001_1;
      patterns[50814] = 25'b11000110_01111100_01000010_1;
      patterns[50815] = 25'b11000110_01111101_01000011_1;
      patterns[50816] = 25'b11000110_01111110_01000100_1;
      patterns[50817] = 25'b11000110_01111111_01000101_1;
      patterns[50818] = 25'b11000110_10000000_01000110_1;
      patterns[50819] = 25'b11000110_10000001_01000111_1;
      patterns[50820] = 25'b11000110_10000010_01001000_1;
      patterns[50821] = 25'b11000110_10000011_01001001_1;
      patterns[50822] = 25'b11000110_10000100_01001010_1;
      patterns[50823] = 25'b11000110_10000101_01001011_1;
      patterns[50824] = 25'b11000110_10000110_01001100_1;
      patterns[50825] = 25'b11000110_10000111_01001101_1;
      patterns[50826] = 25'b11000110_10001000_01001110_1;
      patterns[50827] = 25'b11000110_10001001_01001111_1;
      patterns[50828] = 25'b11000110_10001010_01010000_1;
      patterns[50829] = 25'b11000110_10001011_01010001_1;
      patterns[50830] = 25'b11000110_10001100_01010010_1;
      patterns[50831] = 25'b11000110_10001101_01010011_1;
      patterns[50832] = 25'b11000110_10001110_01010100_1;
      patterns[50833] = 25'b11000110_10001111_01010101_1;
      patterns[50834] = 25'b11000110_10010000_01010110_1;
      patterns[50835] = 25'b11000110_10010001_01010111_1;
      patterns[50836] = 25'b11000110_10010010_01011000_1;
      patterns[50837] = 25'b11000110_10010011_01011001_1;
      patterns[50838] = 25'b11000110_10010100_01011010_1;
      patterns[50839] = 25'b11000110_10010101_01011011_1;
      patterns[50840] = 25'b11000110_10010110_01011100_1;
      patterns[50841] = 25'b11000110_10010111_01011101_1;
      patterns[50842] = 25'b11000110_10011000_01011110_1;
      patterns[50843] = 25'b11000110_10011001_01011111_1;
      patterns[50844] = 25'b11000110_10011010_01100000_1;
      patterns[50845] = 25'b11000110_10011011_01100001_1;
      patterns[50846] = 25'b11000110_10011100_01100010_1;
      patterns[50847] = 25'b11000110_10011101_01100011_1;
      patterns[50848] = 25'b11000110_10011110_01100100_1;
      patterns[50849] = 25'b11000110_10011111_01100101_1;
      patterns[50850] = 25'b11000110_10100000_01100110_1;
      patterns[50851] = 25'b11000110_10100001_01100111_1;
      patterns[50852] = 25'b11000110_10100010_01101000_1;
      patterns[50853] = 25'b11000110_10100011_01101001_1;
      patterns[50854] = 25'b11000110_10100100_01101010_1;
      patterns[50855] = 25'b11000110_10100101_01101011_1;
      patterns[50856] = 25'b11000110_10100110_01101100_1;
      patterns[50857] = 25'b11000110_10100111_01101101_1;
      patterns[50858] = 25'b11000110_10101000_01101110_1;
      patterns[50859] = 25'b11000110_10101001_01101111_1;
      patterns[50860] = 25'b11000110_10101010_01110000_1;
      patterns[50861] = 25'b11000110_10101011_01110001_1;
      patterns[50862] = 25'b11000110_10101100_01110010_1;
      patterns[50863] = 25'b11000110_10101101_01110011_1;
      patterns[50864] = 25'b11000110_10101110_01110100_1;
      patterns[50865] = 25'b11000110_10101111_01110101_1;
      patterns[50866] = 25'b11000110_10110000_01110110_1;
      patterns[50867] = 25'b11000110_10110001_01110111_1;
      patterns[50868] = 25'b11000110_10110010_01111000_1;
      patterns[50869] = 25'b11000110_10110011_01111001_1;
      patterns[50870] = 25'b11000110_10110100_01111010_1;
      patterns[50871] = 25'b11000110_10110101_01111011_1;
      patterns[50872] = 25'b11000110_10110110_01111100_1;
      patterns[50873] = 25'b11000110_10110111_01111101_1;
      patterns[50874] = 25'b11000110_10111000_01111110_1;
      patterns[50875] = 25'b11000110_10111001_01111111_1;
      patterns[50876] = 25'b11000110_10111010_10000000_1;
      patterns[50877] = 25'b11000110_10111011_10000001_1;
      patterns[50878] = 25'b11000110_10111100_10000010_1;
      patterns[50879] = 25'b11000110_10111101_10000011_1;
      patterns[50880] = 25'b11000110_10111110_10000100_1;
      patterns[50881] = 25'b11000110_10111111_10000101_1;
      patterns[50882] = 25'b11000110_11000000_10000110_1;
      patterns[50883] = 25'b11000110_11000001_10000111_1;
      patterns[50884] = 25'b11000110_11000010_10001000_1;
      patterns[50885] = 25'b11000110_11000011_10001001_1;
      patterns[50886] = 25'b11000110_11000100_10001010_1;
      patterns[50887] = 25'b11000110_11000101_10001011_1;
      patterns[50888] = 25'b11000110_11000110_10001100_1;
      patterns[50889] = 25'b11000110_11000111_10001101_1;
      patterns[50890] = 25'b11000110_11001000_10001110_1;
      patterns[50891] = 25'b11000110_11001001_10001111_1;
      patterns[50892] = 25'b11000110_11001010_10010000_1;
      patterns[50893] = 25'b11000110_11001011_10010001_1;
      patterns[50894] = 25'b11000110_11001100_10010010_1;
      patterns[50895] = 25'b11000110_11001101_10010011_1;
      patterns[50896] = 25'b11000110_11001110_10010100_1;
      patterns[50897] = 25'b11000110_11001111_10010101_1;
      patterns[50898] = 25'b11000110_11010000_10010110_1;
      patterns[50899] = 25'b11000110_11010001_10010111_1;
      patterns[50900] = 25'b11000110_11010010_10011000_1;
      patterns[50901] = 25'b11000110_11010011_10011001_1;
      patterns[50902] = 25'b11000110_11010100_10011010_1;
      patterns[50903] = 25'b11000110_11010101_10011011_1;
      patterns[50904] = 25'b11000110_11010110_10011100_1;
      patterns[50905] = 25'b11000110_11010111_10011101_1;
      patterns[50906] = 25'b11000110_11011000_10011110_1;
      patterns[50907] = 25'b11000110_11011001_10011111_1;
      patterns[50908] = 25'b11000110_11011010_10100000_1;
      patterns[50909] = 25'b11000110_11011011_10100001_1;
      patterns[50910] = 25'b11000110_11011100_10100010_1;
      patterns[50911] = 25'b11000110_11011101_10100011_1;
      patterns[50912] = 25'b11000110_11011110_10100100_1;
      patterns[50913] = 25'b11000110_11011111_10100101_1;
      patterns[50914] = 25'b11000110_11100000_10100110_1;
      patterns[50915] = 25'b11000110_11100001_10100111_1;
      patterns[50916] = 25'b11000110_11100010_10101000_1;
      patterns[50917] = 25'b11000110_11100011_10101001_1;
      patterns[50918] = 25'b11000110_11100100_10101010_1;
      patterns[50919] = 25'b11000110_11100101_10101011_1;
      patterns[50920] = 25'b11000110_11100110_10101100_1;
      patterns[50921] = 25'b11000110_11100111_10101101_1;
      patterns[50922] = 25'b11000110_11101000_10101110_1;
      patterns[50923] = 25'b11000110_11101001_10101111_1;
      patterns[50924] = 25'b11000110_11101010_10110000_1;
      patterns[50925] = 25'b11000110_11101011_10110001_1;
      patterns[50926] = 25'b11000110_11101100_10110010_1;
      patterns[50927] = 25'b11000110_11101101_10110011_1;
      patterns[50928] = 25'b11000110_11101110_10110100_1;
      patterns[50929] = 25'b11000110_11101111_10110101_1;
      patterns[50930] = 25'b11000110_11110000_10110110_1;
      patterns[50931] = 25'b11000110_11110001_10110111_1;
      patterns[50932] = 25'b11000110_11110010_10111000_1;
      patterns[50933] = 25'b11000110_11110011_10111001_1;
      patterns[50934] = 25'b11000110_11110100_10111010_1;
      patterns[50935] = 25'b11000110_11110101_10111011_1;
      patterns[50936] = 25'b11000110_11110110_10111100_1;
      patterns[50937] = 25'b11000110_11110111_10111101_1;
      patterns[50938] = 25'b11000110_11111000_10111110_1;
      patterns[50939] = 25'b11000110_11111001_10111111_1;
      patterns[50940] = 25'b11000110_11111010_11000000_1;
      patterns[50941] = 25'b11000110_11111011_11000001_1;
      patterns[50942] = 25'b11000110_11111100_11000010_1;
      patterns[50943] = 25'b11000110_11111101_11000011_1;
      patterns[50944] = 25'b11000110_11111110_11000100_1;
      patterns[50945] = 25'b11000110_11111111_11000101_1;
      patterns[50946] = 25'b11000111_00000000_11000111_0;
      patterns[50947] = 25'b11000111_00000001_11001000_0;
      patterns[50948] = 25'b11000111_00000010_11001001_0;
      patterns[50949] = 25'b11000111_00000011_11001010_0;
      patterns[50950] = 25'b11000111_00000100_11001011_0;
      patterns[50951] = 25'b11000111_00000101_11001100_0;
      patterns[50952] = 25'b11000111_00000110_11001101_0;
      patterns[50953] = 25'b11000111_00000111_11001110_0;
      patterns[50954] = 25'b11000111_00001000_11001111_0;
      patterns[50955] = 25'b11000111_00001001_11010000_0;
      patterns[50956] = 25'b11000111_00001010_11010001_0;
      patterns[50957] = 25'b11000111_00001011_11010010_0;
      patterns[50958] = 25'b11000111_00001100_11010011_0;
      patterns[50959] = 25'b11000111_00001101_11010100_0;
      patterns[50960] = 25'b11000111_00001110_11010101_0;
      patterns[50961] = 25'b11000111_00001111_11010110_0;
      patterns[50962] = 25'b11000111_00010000_11010111_0;
      patterns[50963] = 25'b11000111_00010001_11011000_0;
      patterns[50964] = 25'b11000111_00010010_11011001_0;
      patterns[50965] = 25'b11000111_00010011_11011010_0;
      patterns[50966] = 25'b11000111_00010100_11011011_0;
      patterns[50967] = 25'b11000111_00010101_11011100_0;
      patterns[50968] = 25'b11000111_00010110_11011101_0;
      patterns[50969] = 25'b11000111_00010111_11011110_0;
      patterns[50970] = 25'b11000111_00011000_11011111_0;
      patterns[50971] = 25'b11000111_00011001_11100000_0;
      patterns[50972] = 25'b11000111_00011010_11100001_0;
      patterns[50973] = 25'b11000111_00011011_11100010_0;
      patterns[50974] = 25'b11000111_00011100_11100011_0;
      patterns[50975] = 25'b11000111_00011101_11100100_0;
      patterns[50976] = 25'b11000111_00011110_11100101_0;
      patterns[50977] = 25'b11000111_00011111_11100110_0;
      patterns[50978] = 25'b11000111_00100000_11100111_0;
      patterns[50979] = 25'b11000111_00100001_11101000_0;
      patterns[50980] = 25'b11000111_00100010_11101001_0;
      patterns[50981] = 25'b11000111_00100011_11101010_0;
      patterns[50982] = 25'b11000111_00100100_11101011_0;
      patterns[50983] = 25'b11000111_00100101_11101100_0;
      patterns[50984] = 25'b11000111_00100110_11101101_0;
      patterns[50985] = 25'b11000111_00100111_11101110_0;
      patterns[50986] = 25'b11000111_00101000_11101111_0;
      patterns[50987] = 25'b11000111_00101001_11110000_0;
      patterns[50988] = 25'b11000111_00101010_11110001_0;
      patterns[50989] = 25'b11000111_00101011_11110010_0;
      patterns[50990] = 25'b11000111_00101100_11110011_0;
      patterns[50991] = 25'b11000111_00101101_11110100_0;
      patterns[50992] = 25'b11000111_00101110_11110101_0;
      patterns[50993] = 25'b11000111_00101111_11110110_0;
      patterns[50994] = 25'b11000111_00110000_11110111_0;
      patterns[50995] = 25'b11000111_00110001_11111000_0;
      patterns[50996] = 25'b11000111_00110010_11111001_0;
      patterns[50997] = 25'b11000111_00110011_11111010_0;
      patterns[50998] = 25'b11000111_00110100_11111011_0;
      patterns[50999] = 25'b11000111_00110101_11111100_0;
      patterns[51000] = 25'b11000111_00110110_11111101_0;
      patterns[51001] = 25'b11000111_00110111_11111110_0;
      patterns[51002] = 25'b11000111_00111000_11111111_0;
      patterns[51003] = 25'b11000111_00111001_00000000_1;
      patterns[51004] = 25'b11000111_00111010_00000001_1;
      patterns[51005] = 25'b11000111_00111011_00000010_1;
      patterns[51006] = 25'b11000111_00111100_00000011_1;
      patterns[51007] = 25'b11000111_00111101_00000100_1;
      patterns[51008] = 25'b11000111_00111110_00000101_1;
      patterns[51009] = 25'b11000111_00111111_00000110_1;
      patterns[51010] = 25'b11000111_01000000_00000111_1;
      patterns[51011] = 25'b11000111_01000001_00001000_1;
      patterns[51012] = 25'b11000111_01000010_00001001_1;
      patterns[51013] = 25'b11000111_01000011_00001010_1;
      patterns[51014] = 25'b11000111_01000100_00001011_1;
      patterns[51015] = 25'b11000111_01000101_00001100_1;
      patterns[51016] = 25'b11000111_01000110_00001101_1;
      patterns[51017] = 25'b11000111_01000111_00001110_1;
      patterns[51018] = 25'b11000111_01001000_00001111_1;
      patterns[51019] = 25'b11000111_01001001_00010000_1;
      patterns[51020] = 25'b11000111_01001010_00010001_1;
      patterns[51021] = 25'b11000111_01001011_00010010_1;
      patterns[51022] = 25'b11000111_01001100_00010011_1;
      patterns[51023] = 25'b11000111_01001101_00010100_1;
      patterns[51024] = 25'b11000111_01001110_00010101_1;
      patterns[51025] = 25'b11000111_01001111_00010110_1;
      patterns[51026] = 25'b11000111_01010000_00010111_1;
      patterns[51027] = 25'b11000111_01010001_00011000_1;
      patterns[51028] = 25'b11000111_01010010_00011001_1;
      patterns[51029] = 25'b11000111_01010011_00011010_1;
      patterns[51030] = 25'b11000111_01010100_00011011_1;
      patterns[51031] = 25'b11000111_01010101_00011100_1;
      patterns[51032] = 25'b11000111_01010110_00011101_1;
      patterns[51033] = 25'b11000111_01010111_00011110_1;
      patterns[51034] = 25'b11000111_01011000_00011111_1;
      patterns[51035] = 25'b11000111_01011001_00100000_1;
      patterns[51036] = 25'b11000111_01011010_00100001_1;
      patterns[51037] = 25'b11000111_01011011_00100010_1;
      patterns[51038] = 25'b11000111_01011100_00100011_1;
      patterns[51039] = 25'b11000111_01011101_00100100_1;
      patterns[51040] = 25'b11000111_01011110_00100101_1;
      patterns[51041] = 25'b11000111_01011111_00100110_1;
      patterns[51042] = 25'b11000111_01100000_00100111_1;
      patterns[51043] = 25'b11000111_01100001_00101000_1;
      patterns[51044] = 25'b11000111_01100010_00101001_1;
      patterns[51045] = 25'b11000111_01100011_00101010_1;
      patterns[51046] = 25'b11000111_01100100_00101011_1;
      patterns[51047] = 25'b11000111_01100101_00101100_1;
      patterns[51048] = 25'b11000111_01100110_00101101_1;
      patterns[51049] = 25'b11000111_01100111_00101110_1;
      patterns[51050] = 25'b11000111_01101000_00101111_1;
      patterns[51051] = 25'b11000111_01101001_00110000_1;
      patterns[51052] = 25'b11000111_01101010_00110001_1;
      patterns[51053] = 25'b11000111_01101011_00110010_1;
      patterns[51054] = 25'b11000111_01101100_00110011_1;
      patterns[51055] = 25'b11000111_01101101_00110100_1;
      patterns[51056] = 25'b11000111_01101110_00110101_1;
      patterns[51057] = 25'b11000111_01101111_00110110_1;
      patterns[51058] = 25'b11000111_01110000_00110111_1;
      patterns[51059] = 25'b11000111_01110001_00111000_1;
      patterns[51060] = 25'b11000111_01110010_00111001_1;
      patterns[51061] = 25'b11000111_01110011_00111010_1;
      patterns[51062] = 25'b11000111_01110100_00111011_1;
      patterns[51063] = 25'b11000111_01110101_00111100_1;
      patterns[51064] = 25'b11000111_01110110_00111101_1;
      patterns[51065] = 25'b11000111_01110111_00111110_1;
      patterns[51066] = 25'b11000111_01111000_00111111_1;
      patterns[51067] = 25'b11000111_01111001_01000000_1;
      patterns[51068] = 25'b11000111_01111010_01000001_1;
      patterns[51069] = 25'b11000111_01111011_01000010_1;
      patterns[51070] = 25'b11000111_01111100_01000011_1;
      patterns[51071] = 25'b11000111_01111101_01000100_1;
      patterns[51072] = 25'b11000111_01111110_01000101_1;
      patterns[51073] = 25'b11000111_01111111_01000110_1;
      patterns[51074] = 25'b11000111_10000000_01000111_1;
      patterns[51075] = 25'b11000111_10000001_01001000_1;
      patterns[51076] = 25'b11000111_10000010_01001001_1;
      patterns[51077] = 25'b11000111_10000011_01001010_1;
      patterns[51078] = 25'b11000111_10000100_01001011_1;
      patterns[51079] = 25'b11000111_10000101_01001100_1;
      patterns[51080] = 25'b11000111_10000110_01001101_1;
      patterns[51081] = 25'b11000111_10000111_01001110_1;
      patterns[51082] = 25'b11000111_10001000_01001111_1;
      patterns[51083] = 25'b11000111_10001001_01010000_1;
      patterns[51084] = 25'b11000111_10001010_01010001_1;
      patterns[51085] = 25'b11000111_10001011_01010010_1;
      patterns[51086] = 25'b11000111_10001100_01010011_1;
      patterns[51087] = 25'b11000111_10001101_01010100_1;
      patterns[51088] = 25'b11000111_10001110_01010101_1;
      patterns[51089] = 25'b11000111_10001111_01010110_1;
      patterns[51090] = 25'b11000111_10010000_01010111_1;
      patterns[51091] = 25'b11000111_10010001_01011000_1;
      patterns[51092] = 25'b11000111_10010010_01011001_1;
      patterns[51093] = 25'b11000111_10010011_01011010_1;
      patterns[51094] = 25'b11000111_10010100_01011011_1;
      patterns[51095] = 25'b11000111_10010101_01011100_1;
      patterns[51096] = 25'b11000111_10010110_01011101_1;
      patterns[51097] = 25'b11000111_10010111_01011110_1;
      patterns[51098] = 25'b11000111_10011000_01011111_1;
      patterns[51099] = 25'b11000111_10011001_01100000_1;
      patterns[51100] = 25'b11000111_10011010_01100001_1;
      patterns[51101] = 25'b11000111_10011011_01100010_1;
      patterns[51102] = 25'b11000111_10011100_01100011_1;
      patterns[51103] = 25'b11000111_10011101_01100100_1;
      patterns[51104] = 25'b11000111_10011110_01100101_1;
      patterns[51105] = 25'b11000111_10011111_01100110_1;
      patterns[51106] = 25'b11000111_10100000_01100111_1;
      patterns[51107] = 25'b11000111_10100001_01101000_1;
      patterns[51108] = 25'b11000111_10100010_01101001_1;
      patterns[51109] = 25'b11000111_10100011_01101010_1;
      patterns[51110] = 25'b11000111_10100100_01101011_1;
      patterns[51111] = 25'b11000111_10100101_01101100_1;
      patterns[51112] = 25'b11000111_10100110_01101101_1;
      patterns[51113] = 25'b11000111_10100111_01101110_1;
      patterns[51114] = 25'b11000111_10101000_01101111_1;
      patterns[51115] = 25'b11000111_10101001_01110000_1;
      patterns[51116] = 25'b11000111_10101010_01110001_1;
      patterns[51117] = 25'b11000111_10101011_01110010_1;
      patterns[51118] = 25'b11000111_10101100_01110011_1;
      patterns[51119] = 25'b11000111_10101101_01110100_1;
      patterns[51120] = 25'b11000111_10101110_01110101_1;
      patterns[51121] = 25'b11000111_10101111_01110110_1;
      patterns[51122] = 25'b11000111_10110000_01110111_1;
      patterns[51123] = 25'b11000111_10110001_01111000_1;
      patterns[51124] = 25'b11000111_10110010_01111001_1;
      patterns[51125] = 25'b11000111_10110011_01111010_1;
      patterns[51126] = 25'b11000111_10110100_01111011_1;
      patterns[51127] = 25'b11000111_10110101_01111100_1;
      patterns[51128] = 25'b11000111_10110110_01111101_1;
      patterns[51129] = 25'b11000111_10110111_01111110_1;
      patterns[51130] = 25'b11000111_10111000_01111111_1;
      patterns[51131] = 25'b11000111_10111001_10000000_1;
      patterns[51132] = 25'b11000111_10111010_10000001_1;
      patterns[51133] = 25'b11000111_10111011_10000010_1;
      patterns[51134] = 25'b11000111_10111100_10000011_1;
      patterns[51135] = 25'b11000111_10111101_10000100_1;
      patterns[51136] = 25'b11000111_10111110_10000101_1;
      patterns[51137] = 25'b11000111_10111111_10000110_1;
      patterns[51138] = 25'b11000111_11000000_10000111_1;
      patterns[51139] = 25'b11000111_11000001_10001000_1;
      patterns[51140] = 25'b11000111_11000010_10001001_1;
      patterns[51141] = 25'b11000111_11000011_10001010_1;
      patterns[51142] = 25'b11000111_11000100_10001011_1;
      patterns[51143] = 25'b11000111_11000101_10001100_1;
      patterns[51144] = 25'b11000111_11000110_10001101_1;
      patterns[51145] = 25'b11000111_11000111_10001110_1;
      patterns[51146] = 25'b11000111_11001000_10001111_1;
      patterns[51147] = 25'b11000111_11001001_10010000_1;
      patterns[51148] = 25'b11000111_11001010_10010001_1;
      patterns[51149] = 25'b11000111_11001011_10010010_1;
      patterns[51150] = 25'b11000111_11001100_10010011_1;
      patterns[51151] = 25'b11000111_11001101_10010100_1;
      patterns[51152] = 25'b11000111_11001110_10010101_1;
      patterns[51153] = 25'b11000111_11001111_10010110_1;
      patterns[51154] = 25'b11000111_11010000_10010111_1;
      patterns[51155] = 25'b11000111_11010001_10011000_1;
      patterns[51156] = 25'b11000111_11010010_10011001_1;
      patterns[51157] = 25'b11000111_11010011_10011010_1;
      patterns[51158] = 25'b11000111_11010100_10011011_1;
      patterns[51159] = 25'b11000111_11010101_10011100_1;
      patterns[51160] = 25'b11000111_11010110_10011101_1;
      patterns[51161] = 25'b11000111_11010111_10011110_1;
      patterns[51162] = 25'b11000111_11011000_10011111_1;
      patterns[51163] = 25'b11000111_11011001_10100000_1;
      patterns[51164] = 25'b11000111_11011010_10100001_1;
      patterns[51165] = 25'b11000111_11011011_10100010_1;
      patterns[51166] = 25'b11000111_11011100_10100011_1;
      patterns[51167] = 25'b11000111_11011101_10100100_1;
      patterns[51168] = 25'b11000111_11011110_10100101_1;
      patterns[51169] = 25'b11000111_11011111_10100110_1;
      patterns[51170] = 25'b11000111_11100000_10100111_1;
      patterns[51171] = 25'b11000111_11100001_10101000_1;
      patterns[51172] = 25'b11000111_11100010_10101001_1;
      patterns[51173] = 25'b11000111_11100011_10101010_1;
      patterns[51174] = 25'b11000111_11100100_10101011_1;
      patterns[51175] = 25'b11000111_11100101_10101100_1;
      patterns[51176] = 25'b11000111_11100110_10101101_1;
      patterns[51177] = 25'b11000111_11100111_10101110_1;
      patterns[51178] = 25'b11000111_11101000_10101111_1;
      patterns[51179] = 25'b11000111_11101001_10110000_1;
      patterns[51180] = 25'b11000111_11101010_10110001_1;
      patterns[51181] = 25'b11000111_11101011_10110010_1;
      patterns[51182] = 25'b11000111_11101100_10110011_1;
      patterns[51183] = 25'b11000111_11101101_10110100_1;
      patterns[51184] = 25'b11000111_11101110_10110101_1;
      patterns[51185] = 25'b11000111_11101111_10110110_1;
      patterns[51186] = 25'b11000111_11110000_10110111_1;
      patterns[51187] = 25'b11000111_11110001_10111000_1;
      patterns[51188] = 25'b11000111_11110010_10111001_1;
      patterns[51189] = 25'b11000111_11110011_10111010_1;
      patterns[51190] = 25'b11000111_11110100_10111011_1;
      patterns[51191] = 25'b11000111_11110101_10111100_1;
      patterns[51192] = 25'b11000111_11110110_10111101_1;
      patterns[51193] = 25'b11000111_11110111_10111110_1;
      patterns[51194] = 25'b11000111_11111000_10111111_1;
      patterns[51195] = 25'b11000111_11111001_11000000_1;
      patterns[51196] = 25'b11000111_11111010_11000001_1;
      patterns[51197] = 25'b11000111_11111011_11000010_1;
      patterns[51198] = 25'b11000111_11111100_11000011_1;
      patterns[51199] = 25'b11000111_11111101_11000100_1;
      patterns[51200] = 25'b11000111_11111110_11000101_1;
      patterns[51201] = 25'b11000111_11111111_11000110_1;
      patterns[51202] = 25'b11001000_00000000_11001000_0;
      patterns[51203] = 25'b11001000_00000001_11001001_0;
      patterns[51204] = 25'b11001000_00000010_11001010_0;
      patterns[51205] = 25'b11001000_00000011_11001011_0;
      patterns[51206] = 25'b11001000_00000100_11001100_0;
      patterns[51207] = 25'b11001000_00000101_11001101_0;
      patterns[51208] = 25'b11001000_00000110_11001110_0;
      patterns[51209] = 25'b11001000_00000111_11001111_0;
      patterns[51210] = 25'b11001000_00001000_11010000_0;
      patterns[51211] = 25'b11001000_00001001_11010001_0;
      patterns[51212] = 25'b11001000_00001010_11010010_0;
      patterns[51213] = 25'b11001000_00001011_11010011_0;
      patterns[51214] = 25'b11001000_00001100_11010100_0;
      patterns[51215] = 25'b11001000_00001101_11010101_0;
      patterns[51216] = 25'b11001000_00001110_11010110_0;
      patterns[51217] = 25'b11001000_00001111_11010111_0;
      patterns[51218] = 25'b11001000_00010000_11011000_0;
      patterns[51219] = 25'b11001000_00010001_11011001_0;
      patterns[51220] = 25'b11001000_00010010_11011010_0;
      patterns[51221] = 25'b11001000_00010011_11011011_0;
      patterns[51222] = 25'b11001000_00010100_11011100_0;
      patterns[51223] = 25'b11001000_00010101_11011101_0;
      patterns[51224] = 25'b11001000_00010110_11011110_0;
      patterns[51225] = 25'b11001000_00010111_11011111_0;
      patterns[51226] = 25'b11001000_00011000_11100000_0;
      patterns[51227] = 25'b11001000_00011001_11100001_0;
      patterns[51228] = 25'b11001000_00011010_11100010_0;
      patterns[51229] = 25'b11001000_00011011_11100011_0;
      patterns[51230] = 25'b11001000_00011100_11100100_0;
      patterns[51231] = 25'b11001000_00011101_11100101_0;
      patterns[51232] = 25'b11001000_00011110_11100110_0;
      patterns[51233] = 25'b11001000_00011111_11100111_0;
      patterns[51234] = 25'b11001000_00100000_11101000_0;
      patterns[51235] = 25'b11001000_00100001_11101001_0;
      patterns[51236] = 25'b11001000_00100010_11101010_0;
      patterns[51237] = 25'b11001000_00100011_11101011_0;
      patterns[51238] = 25'b11001000_00100100_11101100_0;
      patterns[51239] = 25'b11001000_00100101_11101101_0;
      patterns[51240] = 25'b11001000_00100110_11101110_0;
      patterns[51241] = 25'b11001000_00100111_11101111_0;
      patterns[51242] = 25'b11001000_00101000_11110000_0;
      patterns[51243] = 25'b11001000_00101001_11110001_0;
      patterns[51244] = 25'b11001000_00101010_11110010_0;
      patterns[51245] = 25'b11001000_00101011_11110011_0;
      patterns[51246] = 25'b11001000_00101100_11110100_0;
      patterns[51247] = 25'b11001000_00101101_11110101_0;
      patterns[51248] = 25'b11001000_00101110_11110110_0;
      patterns[51249] = 25'b11001000_00101111_11110111_0;
      patterns[51250] = 25'b11001000_00110000_11111000_0;
      patterns[51251] = 25'b11001000_00110001_11111001_0;
      patterns[51252] = 25'b11001000_00110010_11111010_0;
      patterns[51253] = 25'b11001000_00110011_11111011_0;
      patterns[51254] = 25'b11001000_00110100_11111100_0;
      patterns[51255] = 25'b11001000_00110101_11111101_0;
      patterns[51256] = 25'b11001000_00110110_11111110_0;
      patterns[51257] = 25'b11001000_00110111_11111111_0;
      patterns[51258] = 25'b11001000_00111000_00000000_1;
      patterns[51259] = 25'b11001000_00111001_00000001_1;
      patterns[51260] = 25'b11001000_00111010_00000010_1;
      patterns[51261] = 25'b11001000_00111011_00000011_1;
      patterns[51262] = 25'b11001000_00111100_00000100_1;
      patterns[51263] = 25'b11001000_00111101_00000101_1;
      patterns[51264] = 25'b11001000_00111110_00000110_1;
      patterns[51265] = 25'b11001000_00111111_00000111_1;
      patterns[51266] = 25'b11001000_01000000_00001000_1;
      patterns[51267] = 25'b11001000_01000001_00001001_1;
      patterns[51268] = 25'b11001000_01000010_00001010_1;
      patterns[51269] = 25'b11001000_01000011_00001011_1;
      patterns[51270] = 25'b11001000_01000100_00001100_1;
      patterns[51271] = 25'b11001000_01000101_00001101_1;
      patterns[51272] = 25'b11001000_01000110_00001110_1;
      patterns[51273] = 25'b11001000_01000111_00001111_1;
      patterns[51274] = 25'b11001000_01001000_00010000_1;
      patterns[51275] = 25'b11001000_01001001_00010001_1;
      patterns[51276] = 25'b11001000_01001010_00010010_1;
      patterns[51277] = 25'b11001000_01001011_00010011_1;
      patterns[51278] = 25'b11001000_01001100_00010100_1;
      patterns[51279] = 25'b11001000_01001101_00010101_1;
      patterns[51280] = 25'b11001000_01001110_00010110_1;
      patterns[51281] = 25'b11001000_01001111_00010111_1;
      patterns[51282] = 25'b11001000_01010000_00011000_1;
      patterns[51283] = 25'b11001000_01010001_00011001_1;
      patterns[51284] = 25'b11001000_01010010_00011010_1;
      patterns[51285] = 25'b11001000_01010011_00011011_1;
      patterns[51286] = 25'b11001000_01010100_00011100_1;
      patterns[51287] = 25'b11001000_01010101_00011101_1;
      patterns[51288] = 25'b11001000_01010110_00011110_1;
      patterns[51289] = 25'b11001000_01010111_00011111_1;
      patterns[51290] = 25'b11001000_01011000_00100000_1;
      patterns[51291] = 25'b11001000_01011001_00100001_1;
      patterns[51292] = 25'b11001000_01011010_00100010_1;
      patterns[51293] = 25'b11001000_01011011_00100011_1;
      patterns[51294] = 25'b11001000_01011100_00100100_1;
      patterns[51295] = 25'b11001000_01011101_00100101_1;
      patterns[51296] = 25'b11001000_01011110_00100110_1;
      patterns[51297] = 25'b11001000_01011111_00100111_1;
      patterns[51298] = 25'b11001000_01100000_00101000_1;
      patterns[51299] = 25'b11001000_01100001_00101001_1;
      patterns[51300] = 25'b11001000_01100010_00101010_1;
      patterns[51301] = 25'b11001000_01100011_00101011_1;
      patterns[51302] = 25'b11001000_01100100_00101100_1;
      patterns[51303] = 25'b11001000_01100101_00101101_1;
      patterns[51304] = 25'b11001000_01100110_00101110_1;
      patterns[51305] = 25'b11001000_01100111_00101111_1;
      patterns[51306] = 25'b11001000_01101000_00110000_1;
      patterns[51307] = 25'b11001000_01101001_00110001_1;
      patterns[51308] = 25'b11001000_01101010_00110010_1;
      patterns[51309] = 25'b11001000_01101011_00110011_1;
      patterns[51310] = 25'b11001000_01101100_00110100_1;
      patterns[51311] = 25'b11001000_01101101_00110101_1;
      patterns[51312] = 25'b11001000_01101110_00110110_1;
      patterns[51313] = 25'b11001000_01101111_00110111_1;
      patterns[51314] = 25'b11001000_01110000_00111000_1;
      patterns[51315] = 25'b11001000_01110001_00111001_1;
      patterns[51316] = 25'b11001000_01110010_00111010_1;
      patterns[51317] = 25'b11001000_01110011_00111011_1;
      patterns[51318] = 25'b11001000_01110100_00111100_1;
      patterns[51319] = 25'b11001000_01110101_00111101_1;
      patterns[51320] = 25'b11001000_01110110_00111110_1;
      patterns[51321] = 25'b11001000_01110111_00111111_1;
      patterns[51322] = 25'b11001000_01111000_01000000_1;
      patterns[51323] = 25'b11001000_01111001_01000001_1;
      patterns[51324] = 25'b11001000_01111010_01000010_1;
      patterns[51325] = 25'b11001000_01111011_01000011_1;
      patterns[51326] = 25'b11001000_01111100_01000100_1;
      patterns[51327] = 25'b11001000_01111101_01000101_1;
      patterns[51328] = 25'b11001000_01111110_01000110_1;
      patterns[51329] = 25'b11001000_01111111_01000111_1;
      patterns[51330] = 25'b11001000_10000000_01001000_1;
      patterns[51331] = 25'b11001000_10000001_01001001_1;
      patterns[51332] = 25'b11001000_10000010_01001010_1;
      patterns[51333] = 25'b11001000_10000011_01001011_1;
      patterns[51334] = 25'b11001000_10000100_01001100_1;
      patterns[51335] = 25'b11001000_10000101_01001101_1;
      patterns[51336] = 25'b11001000_10000110_01001110_1;
      patterns[51337] = 25'b11001000_10000111_01001111_1;
      patterns[51338] = 25'b11001000_10001000_01010000_1;
      patterns[51339] = 25'b11001000_10001001_01010001_1;
      patterns[51340] = 25'b11001000_10001010_01010010_1;
      patterns[51341] = 25'b11001000_10001011_01010011_1;
      patterns[51342] = 25'b11001000_10001100_01010100_1;
      patterns[51343] = 25'b11001000_10001101_01010101_1;
      patterns[51344] = 25'b11001000_10001110_01010110_1;
      patterns[51345] = 25'b11001000_10001111_01010111_1;
      patterns[51346] = 25'b11001000_10010000_01011000_1;
      patterns[51347] = 25'b11001000_10010001_01011001_1;
      patterns[51348] = 25'b11001000_10010010_01011010_1;
      patterns[51349] = 25'b11001000_10010011_01011011_1;
      patterns[51350] = 25'b11001000_10010100_01011100_1;
      patterns[51351] = 25'b11001000_10010101_01011101_1;
      patterns[51352] = 25'b11001000_10010110_01011110_1;
      patterns[51353] = 25'b11001000_10010111_01011111_1;
      patterns[51354] = 25'b11001000_10011000_01100000_1;
      patterns[51355] = 25'b11001000_10011001_01100001_1;
      patterns[51356] = 25'b11001000_10011010_01100010_1;
      patterns[51357] = 25'b11001000_10011011_01100011_1;
      patterns[51358] = 25'b11001000_10011100_01100100_1;
      patterns[51359] = 25'b11001000_10011101_01100101_1;
      patterns[51360] = 25'b11001000_10011110_01100110_1;
      patterns[51361] = 25'b11001000_10011111_01100111_1;
      patterns[51362] = 25'b11001000_10100000_01101000_1;
      patterns[51363] = 25'b11001000_10100001_01101001_1;
      patterns[51364] = 25'b11001000_10100010_01101010_1;
      patterns[51365] = 25'b11001000_10100011_01101011_1;
      patterns[51366] = 25'b11001000_10100100_01101100_1;
      patterns[51367] = 25'b11001000_10100101_01101101_1;
      patterns[51368] = 25'b11001000_10100110_01101110_1;
      patterns[51369] = 25'b11001000_10100111_01101111_1;
      patterns[51370] = 25'b11001000_10101000_01110000_1;
      patterns[51371] = 25'b11001000_10101001_01110001_1;
      patterns[51372] = 25'b11001000_10101010_01110010_1;
      patterns[51373] = 25'b11001000_10101011_01110011_1;
      patterns[51374] = 25'b11001000_10101100_01110100_1;
      patterns[51375] = 25'b11001000_10101101_01110101_1;
      patterns[51376] = 25'b11001000_10101110_01110110_1;
      patterns[51377] = 25'b11001000_10101111_01110111_1;
      patterns[51378] = 25'b11001000_10110000_01111000_1;
      patterns[51379] = 25'b11001000_10110001_01111001_1;
      patterns[51380] = 25'b11001000_10110010_01111010_1;
      patterns[51381] = 25'b11001000_10110011_01111011_1;
      patterns[51382] = 25'b11001000_10110100_01111100_1;
      patterns[51383] = 25'b11001000_10110101_01111101_1;
      patterns[51384] = 25'b11001000_10110110_01111110_1;
      patterns[51385] = 25'b11001000_10110111_01111111_1;
      patterns[51386] = 25'b11001000_10111000_10000000_1;
      patterns[51387] = 25'b11001000_10111001_10000001_1;
      patterns[51388] = 25'b11001000_10111010_10000010_1;
      patterns[51389] = 25'b11001000_10111011_10000011_1;
      patterns[51390] = 25'b11001000_10111100_10000100_1;
      patterns[51391] = 25'b11001000_10111101_10000101_1;
      patterns[51392] = 25'b11001000_10111110_10000110_1;
      patterns[51393] = 25'b11001000_10111111_10000111_1;
      patterns[51394] = 25'b11001000_11000000_10001000_1;
      patterns[51395] = 25'b11001000_11000001_10001001_1;
      patterns[51396] = 25'b11001000_11000010_10001010_1;
      patterns[51397] = 25'b11001000_11000011_10001011_1;
      patterns[51398] = 25'b11001000_11000100_10001100_1;
      patterns[51399] = 25'b11001000_11000101_10001101_1;
      patterns[51400] = 25'b11001000_11000110_10001110_1;
      patterns[51401] = 25'b11001000_11000111_10001111_1;
      patterns[51402] = 25'b11001000_11001000_10010000_1;
      patterns[51403] = 25'b11001000_11001001_10010001_1;
      patterns[51404] = 25'b11001000_11001010_10010010_1;
      patterns[51405] = 25'b11001000_11001011_10010011_1;
      patterns[51406] = 25'b11001000_11001100_10010100_1;
      patterns[51407] = 25'b11001000_11001101_10010101_1;
      patterns[51408] = 25'b11001000_11001110_10010110_1;
      patterns[51409] = 25'b11001000_11001111_10010111_1;
      patterns[51410] = 25'b11001000_11010000_10011000_1;
      patterns[51411] = 25'b11001000_11010001_10011001_1;
      patterns[51412] = 25'b11001000_11010010_10011010_1;
      patterns[51413] = 25'b11001000_11010011_10011011_1;
      patterns[51414] = 25'b11001000_11010100_10011100_1;
      patterns[51415] = 25'b11001000_11010101_10011101_1;
      patterns[51416] = 25'b11001000_11010110_10011110_1;
      patterns[51417] = 25'b11001000_11010111_10011111_1;
      patterns[51418] = 25'b11001000_11011000_10100000_1;
      patterns[51419] = 25'b11001000_11011001_10100001_1;
      patterns[51420] = 25'b11001000_11011010_10100010_1;
      patterns[51421] = 25'b11001000_11011011_10100011_1;
      patterns[51422] = 25'b11001000_11011100_10100100_1;
      patterns[51423] = 25'b11001000_11011101_10100101_1;
      patterns[51424] = 25'b11001000_11011110_10100110_1;
      patterns[51425] = 25'b11001000_11011111_10100111_1;
      patterns[51426] = 25'b11001000_11100000_10101000_1;
      patterns[51427] = 25'b11001000_11100001_10101001_1;
      patterns[51428] = 25'b11001000_11100010_10101010_1;
      patterns[51429] = 25'b11001000_11100011_10101011_1;
      patterns[51430] = 25'b11001000_11100100_10101100_1;
      patterns[51431] = 25'b11001000_11100101_10101101_1;
      patterns[51432] = 25'b11001000_11100110_10101110_1;
      patterns[51433] = 25'b11001000_11100111_10101111_1;
      patterns[51434] = 25'b11001000_11101000_10110000_1;
      patterns[51435] = 25'b11001000_11101001_10110001_1;
      patterns[51436] = 25'b11001000_11101010_10110010_1;
      patterns[51437] = 25'b11001000_11101011_10110011_1;
      patterns[51438] = 25'b11001000_11101100_10110100_1;
      patterns[51439] = 25'b11001000_11101101_10110101_1;
      patterns[51440] = 25'b11001000_11101110_10110110_1;
      patterns[51441] = 25'b11001000_11101111_10110111_1;
      patterns[51442] = 25'b11001000_11110000_10111000_1;
      patterns[51443] = 25'b11001000_11110001_10111001_1;
      patterns[51444] = 25'b11001000_11110010_10111010_1;
      patterns[51445] = 25'b11001000_11110011_10111011_1;
      patterns[51446] = 25'b11001000_11110100_10111100_1;
      patterns[51447] = 25'b11001000_11110101_10111101_1;
      patterns[51448] = 25'b11001000_11110110_10111110_1;
      patterns[51449] = 25'b11001000_11110111_10111111_1;
      patterns[51450] = 25'b11001000_11111000_11000000_1;
      patterns[51451] = 25'b11001000_11111001_11000001_1;
      patterns[51452] = 25'b11001000_11111010_11000010_1;
      patterns[51453] = 25'b11001000_11111011_11000011_1;
      patterns[51454] = 25'b11001000_11111100_11000100_1;
      patterns[51455] = 25'b11001000_11111101_11000101_1;
      patterns[51456] = 25'b11001000_11111110_11000110_1;
      patterns[51457] = 25'b11001000_11111111_11000111_1;
      patterns[51458] = 25'b11001001_00000000_11001001_0;
      patterns[51459] = 25'b11001001_00000001_11001010_0;
      patterns[51460] = 25'b11001001_00000010_11001011_0;
      patterns[51461] = 25'b11001001_00000011_11001100_0;
      patterns[51462] = 25'b11001001_00000100_11001101_0;
      patterns[51463] = 25'b11001001_00000101_11001110_0;
      patterns[51464] = 25'b11001001_00000110_11001111_0;
      patterns[51465] = 25'b11001001_00000111_11010000_0;
      patterns[51466] = 25'b11001001_00001000_11010001_0;
      patterns[51467] = 25'b11001001_00001001_11010010_0;
      patterns[51468] = 25'b11001001_00001010_11010011_0;
      patterns[51469] = 25'b11001001_00001011_11010100_0;
      patterns[51470] = 25'b11001001_00001100_11010101_0;
      patterns[51471] = 25'b11001001_00001101_11010110_0;
      patterns[51472] = 25'b11001001_00001110_11010111_0;
      patterns[51473] = 25'b11001001_00001111_11011000_0;
      patterns[51474] = 25'b11001001_00010000_11011001_0;
      patterns[51475] = 25'b11001001_00010001_11011010_0;
      patterns[51476] = 25'b11001001_00010010_11011011_0;
      patterns[51477] = 25'b11001001_00010011_11011100_0;
      patterns[51478] = 25'b11001001_00010100_11011101_0;
      patterns[51479] = 25'b11001001_00010101_11011110_0;
      patterns[51480] = 25'b11001001_00010110_11011111_0;
      patterns[51481] = 25'b11001001_00010111_11100000_0;
      patterns[51482] = 25'b11001001_00011000_11100001_0;
      patterns[51483] = 25'b11001001_00011001_11100010_0;
      patterns[51484] = 25'b11001001_00011010_11100011_0;
      patterns[51485] = 25'b11001001_00011011_11100100_0;
      patterns[51486] = 25'b11001001_00011100_11100101_0;
      patterns[51487] = 25'b11001001_00011101_11100110_0;
      patterns[51488] = 25'b11001001_00011110_11100111_0;
      patterns[51489] = 25'b11001001_00011111_11101000_0;
      patterns[51490] = 25'b11001001_00100000_11101001_0;
      patterns[51491] = 25'b11001001_00100001_11101010_0;
      patterns[51492] = 25'b11001001_00100010_11101011_0;
      patterns[51493] = 25'b11001001_00100011_11101100_0;
      patterns[51494] = 25'b11001001_00100100_11101101_0;
      patterns[51495] = 25'b11001001_00100101_11101110_0;
      patterns[51496] = 25'b11001001_00100110_11101111_0;
      patterns[51497] = 25'b11001001_00100111_11110000_0;
      patterns[51498] = 25'b11001001_00101000_11110001_0;
      patterns[51499] = 25'b11001001_00101001_11110010_0;
      patterns[51500] = 25'b11001001_00101010_11110011_0;
      patterns[51501] = 25'b11001001_00101011_11110100_0;
      patterns[51502] = 25'b11001001_00101100_11110101_0;
      patterns[51503] = 25'b11001001_00101101_11110110_0;
      patterns[51504] = 25'b11001001_00101110_11110111_0;
      patterns[51505] = 25'b11001001_00101111_11111000_0;
      patterns[51506] = 25'b11001001_00110000_11111001_0;
      patterns[51507] = 25'b11001001_00110001_11111010_0;
      patterns[51508] = 25'b11001001_00110010_11111011_0;
      patterns[51509] = 25'b11001001_00110011_11111100_0;
      patterns[51510] = 25'b11001001_00110100_11111101_0;
      patterns[51511] = 25'b11001001_00110101_11111110_0;
      patterns[51512] = 25'b11001001_00110110_11111111_0;
      patterns[51513] = 25'b11001001_00110111_00000000_1;
      patterns[51514] = 25'b11001001_00111000_00000001_1;
      patterns[51515] = 25'b11001001_00111001_00000010_1;
      patterns[51516] = 25'b11001001_00111010_00000011_1;
      patterns[51517] = 25'b11001001_00111011_00000100_1;
      patterns[51518] = 25'b11001001_00111100_00000101_1;
      patterns[51519] = 25'b11001001_00111101_00000110_1;
      patterns[51520] = 25'b11001001_00111110_00000111_1;
      patterns[51521] = 25'b11001001_00111111_00001000_1;
      patterns[51522] = 25'b11001001_01000000_00001001_1;
      patterns[51523] = 25'b11001001_01000001_00001010_1;
      patterns[51524] = 25'b11001001_01000010_00001011_1;
      patterns[51525] = 25'b11001001_01000011_00001100_1;
      patterns[51526] = 25'b11001001_01000100_00001101_1;
      patterns[51527] = 25'b11001001_01000101_00001110_1;
      patterns[51528] = 25'b11001001_01000110_00001111_1;
      patterns[51529] = 25'b11001001_01000111_00010000_1;
      patterns[51530] = 25'b11001001_01001000_00010001_1;
      patterns[51531] = 25'b11001001_01001001_00010010_1;
      patterns[51532] = 25'b11001001_01001010_00010011_1;
      patterns[51533] = 25'b11001001_01001011_00010100_1;
      patterns[51534] = 25'b11001001_01001100_00010101_1;
      patterns[51535] = 25'b11001001_01001101_00010110_1;
      patterns[51536] = 25'b11001001_01001110_00010111_1;
      patterns[51537] = 25'b11001001_01001111_00011000_1;
      patterns[51538] = 25'b11001001_01010000_00011001_1;
      patterns[51539] = 25'b11001001_01010001_00011010_1;
      patterns[51540] = 25'b11001001_01010010_00011011_1;
      patterns[51541] = 25'b11001001_01010011_00011100_1;
      patterns[51542] = 25'b11001001_01010100_00011101_1;
      patterns[51543] = 25'b11001001_01010101_00011110_1;
      patterns[51544] = 25'b11001001_01010110_00011111_1;
      patterns[51545] = 25'b11001001_01010111_00100000_1;
      patterns[51546] = 25'b11001001_01011000_00100001_1;
      patterns[51547] = 25'b11001001_01011001_00100010_1;
      patterns[51548] = 25'b11001001_01011010_00100011_1;
      patterns[51549] = 25'b11001001_01011011_00100100_1;
      patterns[51550] = 25'b11001001_01011100_00100101_1;
      patterns[51551] = 25'b11001001_01011101_00100110_1;
      patterns[51552] = 25'b11001001_01011110_00100111_1;
      patterns[51553] = 25'b11001001_01011111_00101000_1;
      patterns[51554] = 25'b11001001_01100000_00101001_1;
      patterns[51555] = 25'b11001001_01100001_00101010_1;
      patterns[51556] = 25'b11001001_01100010_00101011_1;
      patterns[51557] = 25'b11001001_01100011_00101100_1;
      patterns[51558] = 25'b11001001_01100100_00101101_1;
      patterns[51559] = 25'b11001001_01100101_00101110_1;
      patterns[51560] = 25'b11001001_01100110_00101111_1;
      patterns[51561] = 25'b11001001_01100111_00110000_1;
      patterns[51562] = 25'b11001001_01101000_00110001_1;
      patterns[51563] = 25'b11001001_01101001_00110010_1;
      patterns[51564] = 25'b11001001_01101010_00110011_1;
      patterns[51565] = 25'b11001001_01101011_00110100_1;
      patterns[51566] = 25'b11001001_01101100_00110101_1;
      patterns[51567] = 25'b11001001_01101101_00110110_1;
      patterns[51568] = 25'b11001001_01101110_00110111_1;
      patterns[51569] = 25'b11001001_01101111_00111000_1;
      patterns[51570] = 25'b11001001_01110000_00111001_1;
      patterns[51571] = 25'b11001001_01110001_00111010_1;
      patterns[51572] = 25'b11001001_01110010_00111011_1;
      patterns[51573] = 25'b11001001_01110011_00111100_1;
      patterns[51574] = 25'b11001001_01110100_00111101_1;
      patterns[51575] = 25'b11001001_01110101_00111110_1;
      patterns[51576] = 25'b11001001_01110110_00111111_1;
      patterns[51577] = 25'b11001001_01110111_01000000_1;
      patterns[51578] = 25'b11001001_01111000_01000001_1;
      patterns[51579] = 25'b11001001_01111001_01000010_1;
      patterns[51580] = 25'b11001001_01111010_01000011_1;
      patterns[51581] = 25'b11001001_01111011_01000100_1;
      patterns[51582] = 25'b11001001_01111100_01000101_1;
      patterns[51583] = 25'b11001001_01111101_01000110_1;
      patterns[51584] = 25'b11001001_01111110_01000111_1;
      patterns[51585] = 25'b11001001_01111111_01001000_1;
      patterns[51586] = 25'b11001001_10000000_01001001_1;
      patterns[51587] = 25'b11001001_10000001_01001010_1;
      patterns[51588] = 25'b11001001_10000010_01001011_1;
      patterns[51589] = 25'b11001001_10000011_01001100_1;
      patterns[51590] = 25'b11001001_10000100_01001101_1;
      patterns[51591] = 25'b11001001_10000101_01001110_1;
      patterns[51592] = 25'b11001001_10000110_01001111_1;
      patterns[51593] = 25'b11001001_10000111_01010000_1;
      patterns[51594] = 25'b11001001_10001000_01010001_1;
      patterns[51595] = 25'b11001001_10001001_01010010_1;
      patterns[51596] = 25'b11001001_10001010_01010011_1;
      patterns[51597] = 25'b11001001_10001011_01010100_1;
      patterns[51598] = 25'b11001001_10001100_01010101_1;
      patterns[51599] = 25'b11001001_10001101_01010110_1;
      patterns[51600] = 25'b11001001_10001110_01010111_1;
      patterns[51601] = 25'b11001001_10001111_01011000_1;
      patterns[51602] = 25'b11001001_10010000_01011001_1;
      patterns[51603] = 25'b11001001_10010001_01011010_1;
      patterns[51604] = 25'b11001001_10010010_01011011_1;
      patterns[51605] = 25'b11001001_10010011_01011100_1;
      patterns[51606] = 25'b11001001_10010100_01011101_1;
      patterns[51607] = 25'b11001001_10010101_01011110_1;
      patterns[51608] = 25'b11001001_10010110_01011111_1;
      patterns[51609] = 25'b11001001_10010111_01100000_1;
      patterns[51610] = 25'b11001001_10011000_01100001_1;
      patterns[51611] = 25'b11001001_10011001_01100010_1;
      patterns[51612] = 25'b11001001_10011010_01100011_1;
      patterns[51613] = 25'b11001001_10011011_01100100_1;
      patterns[51614] = 25'b11001001_10011100_01100101_1;
      patterns[51615] = 25'b11001001_10011101_01100110_1;
      patterns[51616] = 25'b11001001_10011110_01100111_1;
      patterns[51617] = 25'b11001001_10011111_01101000_1;
      patterns[51618] = 25'b11001001_10100000_01101001_1;
      patterns[51619] = 25'b11001001_10100001_01101010_1;
      patterns[51620] = 25'b11001001_10100010_01101011_1;
      patterns[51621] = 25'b11001001_10100011_01101100_1;
      patterns[51622] = 25'b11001001_10100100_01101101_1;
      patterns[51623] = 25'b11001001_10100101_01101110_1;
      patterns[51624] = 25'b11001001_10100110_01101111_1;
      patterns[51625] = 25'b11001001_10100111_01110000_1;
      patterns[51626] = 25'b11001001_10101000_01110001_1;
      patterns[51627] = 25'b11001001_10101001_01110010_1;
      patterns[51628] = 25'b11001001_10101010_01110011_1;
      patterns[51629] = 25'b11001001_10101011_01110100_1;
      patterns[51630] = 25'b11001001_10101100_01110101_1;
      patterns[51631] = 25'b11001001_10101101_01110110_1;
      patterns[51632] = 25'b11001001_10101110_01110111_1;
      patterns[51633] = 25'b11001001_10101111_01111000_1;
      patterns[51634] = 25'b11001001_10110000_01111001_1;
      patterns[51635] = 25'b11001001_10110001_01111010_1;
      patterns[51636] = 25'b11001001_10110010_01111011_1;
      patterns[51637] = 25'b11001001_10110011_01111100_1;
      patterns[51638] = 25'b11001001_10110100_01111101_1;
      patterns[51639] = 25'b11001001_10110101_01111110_1;
      patterns[51640] = 25'b11001001_10110110_01111111_1;
      patterns[51641] = 25'b11001001_10110111_10000000_1;
      patterns[51642] = 25'b11001001_10111000_10000001_1;
      patterns[51643] = 25'b11001001_10111001_10000010_1;
      patterns[51644] = 25'b11001001_10111010_10000011_1;
      patterns[51645] = 25'b11001001_10111011_10000100_1;
      patterns[51646] = 25'b11001001_10111100_10000101_1;
      patterns[51647] = 25'b11001001_10111101_10000110_1;
      patterns[51648] = 25'b11001001_10111110_10000111_1;
      patterns[51649] = 25'b11001001_10111111_10001000_1;
      patterns[51650] = 25'b11001001_11000000_10001001_1;
      patterns[51651] = 25'b11001001_11000001_10001010_1;
      patterns[51652] = 25'b11001001_11000010_10001011_1;
      patterns[51653] = 25'b11001001_11000011_10001100_1;
      patterns[51654] = 25'b11001001_11000100_10001101_1;
      patterns[51655] = 25'b11001001_11000101_10001110_1;
      patterns[51656] = 25'b11001001_11000110_10001111_1;
      patterns[51657] = 25'b11001001_11000111_10010000_1;
      patterns[51658] = 25'b11001001_11001000_10010001_1;
      patterns[51659] = 25'b11001001_11001001_10010010_1;
      patterns[51660] = 25'b11001001_11001010_10010011_1;
      patterns[51661] = 25'b11001001_11001011_10010100_1;
      patterns[51662] = 25'b11001001_11001100_10010101_1;
      patterns[51663] = 25'b11001001_11001101_10010110_1;
      patterns[51664] = 25'b11001001_11001110_10010111_1;
      patterns[51665] = 25'b11001001_11001111_10011000_1;
      patterns[51666] = 25'b11001001_11010000_10011001_1;
      patterns[51667] = 25'b11001001_11010001_10011010_1;
      patterns[51668] = 25'b11001001_11010010_10011011_1;
      patterns[51669] = 25'b11001001_11010011_10011100_1;
      patterns[51670] = 25'b11001001_11010100_10011101_1;
      patterns[51671] = 25'b11001001_11010101_10011110_1;
      patterns[51672] = 25'b11001001_11010110_10011111_1;
      patterns[51673] = 25'b11001001_11010111_10100000_1;
      patterns[51674] = 25'b11001001_11011000_10100001_1;
      patterns[51675] = 25'b11001001_11011001_10100010_1;
      patterns[51676] = 25'b11001001_11011010_10100011_1;
      patterns[51677] = 25'b11001001_11011011_10100100_1;
      patterns[51678] = 25'b11001001_11011100_10100101_1;
      patterns[51679] = 25'b11001001_11011101_10100110_1;
      patterns[51680] = 25'b11001001_11011110_10100111_1;
      patterns[51681] = 25'b11001001_11011111_10101000_1;
      patterns[51682] = 25'b11001001_11100000_10101001_1;
      patterns[51683] = 25'b11001001_11100001_10101010_1;
      patterns[51684] = 25'b11001001_11100010_10101011_1;
      patterns[51685] = 25'b11001001_11100011_10101100_1;
      patterns[51686] = 25'b11001001_11100100_10101101_1;
      patterns[51687] = 25'b11001001_11100101_10101110_1;
      patterns[51688] = 25'b11001001_11100110_10101111_1;
      patterns[51689] = 25'b11001001_11100111_10110000_1;
      patterns[51690] = 25'b11001001_11101000_10110001_1;
      patterns[51691] = 25'b11001001_11101001_10110010_1;
      patterns[51692] = 25'b11001001_11101010_10110011_1;
      patterns[51693] = 25'b11001001_11101011_10110100_1;
      patterns[51694] = 25'b11001001_11101100_10110101_1;
      patterns[51695] = 25'b11001001_11101101_10110110_1;
      patterns[51696] = 25'b11001001_11101110_10110111_1;
      patterns[51697] = 25'b11001001_11101111_10111000_1;
      patterns[51698] = 25'b11001001_11110000_10111001_1;
      patterns[51699] = 25'b11001001_11110001_10111010_1;
      patterns[51700] = 25'b11001001_11110010_10111011_1;
      patterns[51701] = 25'b11001001_11110011_10111100_1;
      patterns[51702] = 25'b11001001_11110100_10111101_1;
      patterns[51703] = 25'b11001001_11110101_10111110_1;
      patterns[51704] = 25'b11001001_11110110_10111111_1;
      patterns[51705] = 25'b11001001_11110111_11000000_1;
      patterns[51706] = 25'b11001001_11111000_11000001_1;
      patterns[51707] = 25'b11001001_11111001_11000010_1;
      patterns[51708] = 25'b11001001_11111010_11000011_1;
      patterns[51709] = 25'b11001001_11111011_11000100_1;
      patterns[51710] = 25'b11001001_11111100_11000101_1;
      patterns[51711] = 25'b11001001_11111101_11000110_1;
      patterns[51712] = 25'b11001001_11111110_11000111_1;
      patterns[51713] = 25'b11001001_11111111_11001000_1;
      patterns[51714] = 25'b11001010_00000000_11001010_0;
      patterns[51715] = 25'b11001010_00000001_11001011_0;
      patterns[51716] = 25'b11001010_00000010_11001100_0;
      patterns[51717] = 25'b11001010_00000011_11001101_0;
      patterns[51718] = 25'b11001010_00000100_11001110_0;
      patterns[51719] = 25'b11001010_00000101_11001111_0;
      patterns[51720] = 25'b11001010_00000110_11010000_0;
      patterns[51721] = 25'b11001010_00000111_11010001_0;
      patterns[51722] = 25'b11001010_00001000_11010010_0;
      patterns[51723] = 25'b11001010_00001001_11010011_0;
      patterns[51724] = 25'b11001010_00001010_11010100_0;
      patterns[51725] = 25'b11001010_00001011_11010101_0;
      patterns[51726] = 25'b11001010_00001100_11010110_0;
      patterns[51727] = 25'b11001010_00001101_11010111_0;
      patterns[51728] = 25'b11001010_00001110_11011000_0;
      patterns[51729] = 25'b11001010_00001111_11011001_0;
      patterns[51730] = 25'b11001010_00010000_11011010_0;
      patterns[51731] = 25'b11001010_00010001_11011011_0;
      patterns[51732] = 25'b11001010_00010010_11011100_0;
      patterns[51733] = 25'b11001010_00010011_11011101_0;
      patterns[51734] = 25'b11001010_00010100_11011110_0;
      patterns[51735] = 25'b11001010_00010101_11011111_0;
      patterns[51736] = 25'b11001010_00010110_11100000_0;
      patterns[51737] = 25'b11001010_00010111_11100001_0;
      patterns[51738] = 25'b11001010_00011000_11100010_0;
      patterns[51739] = 25'b11001010_00011001_11100011_0;
      patterns[51740] = 25'b11001010_00011010_11100100_0;
      patterns[51741] = 25'b11001010_00011011_11100101_0;
      patterns[51742] = 25'b11001010_00011100_11100110_0;
      patterns[51743] = 25'b11001010_00011101_11100111_0;
      patterns[51744] = 25'b11001010_00011110_11101000_0;
      patterns[51745] = 25'b11001010_00011111_11101001_0;
      patterns[51746] = 25'b11001010_00100000_11101010_0;
      patterns[51747] = 25'b11001010_00100001_11101011_0;
      patterns[51748] = 25'b11001010_00100010_11101100_0;
      patterns[51749] = 25'b11001010_00100011_11101101_0;
      patterns[51750] = 25'b11001010_00100100_11101110_0;
      patterns[51751] = 25'b11001010_00100101_11101111_0;
      patterns[51752] = 25'b11001010_00100110_11110000_0;
      patterns[51753] = 25'b11001010_00100111_11110001_0;
      patterns[51754] = 25'b11001010_00101000_11110010_0;
      patterns[51755] = 25'b11001010_00101001_11110011_0;
      patterns[51756] = 25'b11001010_00101010_11110100_0;
      patterns[51757] = 25'b11001010_00101011_11110101_0;
      patterns[51758] = 25'b11001010_00101100_11110110_0;
      patterns[51759] = 25'b11001010_00101101_11110111_0;
      patterns[51760] = 25'b11001010_00101110_11111000_0;
      patterns[51761] = 25'b11001010_00101111_11111001_0;
      patterns[51762] = 25'b11001010_00110000_11111010_0;
      patterns[51763] = 25'b11001010_00110001_11111011_0;
      patterns[51764] = 25'b11001010_00110010_11111100_0;
      patterns[51765] = 25'b11001010_00110011_11111101_0;
      patterns[51766] = 25'b11001010_00110100_11111110_0;
      patterns[51767] = 25'b11001010_00110101_11111111_0;
      patterns[51768] = 25'b11001010_00110110_00000000_1;
      patterns[51769] = 25'b11001010_00110111_00000001_1;
      patterns[51770] = 25'b11001010_00111000_00000010_1;
      patterns[51771] = 25'b11001010_00111001_00000011_1;
      patterns[51772] = 25'b11001010_00111010_00000100_1;
      patterns[51773] = 25'b11001010_00111011_00000101_1;
      patterns[51774] = 25'b11001010_00111100_00000110_1;
      patterns[51775] = 25'b11001010_00111101_00000111_1;
      patterns[51776] = 25'b11001010_00111110_00001000_1;
      patterns[51777] = 25'b11001010_00111111_00001001_1;
      patterns[51778] = 25'b11001010_01000000_00001010_1;
      patterns[51779] = 25'b11001010_01000001_00001011_1;
      patterns[51780] = 25'b11001010_01000010_00001100_1;
      patterns[51781] = 25'b11001010_01000011_00001101_1;
      patterns[51782] = 25'b11001010_01000100_00001110_1;
      patterns[51783] = 25'b11001010_01000101_00001111_1;
      patterns[51784] = 25'b11001010_01000110_00010000_1;
      patterns[51785] = 25'b11001010_01000111_00010001_1;
      patterns[51786] = 25'b11001010_01001000_00010010_1;
      patterns[51787] = 25'b11001010_01001001_00010011_1;
      patterns[51788] = 25'b11001010_01001010_00010100_1;
      patterns[51789] = 25'b11001010_01001011_00010101_1;
      patterns[51790] = 25'b11001010_01001100_00010110_1;
      patterns[51791] = 25'b11001010_01001101_00010111_1;
      patterns[51792] = 25'b11001010_01001110_00011000_1;
      patterns[51793] = 25'b11001010_01001111_00011001_1;
      patterns[51794] = 25'b11001010_01010000_00011010_1;
      patterns[51795] = 25'b11001010_01010001_00011011_1;
      patterns[51796] = 25'b11001010_01010010_00011100_1;
      patterns[51797] = 25'b11001010_01010011_00011101_1;
      patterns[51798] = 25'b11001010_01010100_00011110_1;
      patterns[51799] = 25'b11001010_01010101_00011111_1;
      patterns[51800] = 25'b11001010_01010110_00100000_1;
      patterns[51801] = 25'b11001010_01010111_00100001_1;
      patterns[51802] = 25'b11001010_01011000_00100010_1;
      patterns[51803] = 25'b11001010_01011001_00100011_1;
      patterns[51804] = 25'b11001010_01011010_00100100_1;
      patterns[51805] = 25'b11001010_01011011_00100101_1;
      patterns[51806] = 25'b11001010_01011100_00100110_1;
      patterns[51807] = 25'b11001010_01011101_00100111_1;
      patterns[51808] = 25'b11001010_01011110_00101000_1;
      patterns[51809] = 25'b11001010_01011111_00101001_1;
      patterns[51810] = 25'b11001010_01100000_00101010_1;
      patterns[51811] = 25'b11001010_01100001_00101011_1;
      patterns[51812] = 25'b11001010_01100010_00101100_1;
      patterns[51813] = 25'b11001010_01100011_00101101_1;
      patterns[51814] = 25'b11001010_01100100_00101110_1;
      patterns[51815] = 25'b11001010_01100101_00101111_1;
      patterns[51816] = 25'b11001010_01100110_00110000_1;
      patterns[51817] = 25'b11001010_01100111_00110001_1;
      patterns[51818] = 25'b11001010_01101000_00110010_1;
      patterns[51819] = 25'b11001010_01101001_00110011_1;
      patterns[51820] = 25'b11001010_01101010_00110100_1;
      patterns[51821] = 25'b11001010_01101011_00110101_1;
      patterns[51822] = 25'b11001010_01101100_00110110_1;
      patterns[51823] = 25'b11001010_01101101_00110111_1;
      patterns[51824] = 25'b11001010_01101110_00111000_1;
      patterns[51825] = 25'b11001010_01101111_00111001_1;
      patterns[51826] = 25'b11001010_01110000_00111010_1;
      patterns[51827] = 25'b11001010_01110001_00111011_1;
      patterns[51828] = 25'b11001010_01110010_00111100_1;
      patterns[51829] = 25'b11001010_01110011_00111101_1;
      patterns[51830] = 25'b11001010_01110100_00111110_1;
      patterns[51831] = 25'b11001010_01110101_00111111_1;
      patterns[51832] = 25'b11001010_01110110_01000000_1;
      patterns[51833] = 25'b11001010_01110111_01000001_1;
      patterns[51834] = 25'b11001010_01111000_01000010_1;
      patterns[51835] = 25'b11001010_01111001_01000011_1;
      patterns[51836] = 25'b11001010_01111010_01000100_1;
      patterns[51837] = 25'b11001010_01111011_01000101_1;
      patterns[51838] = 25'b11001010_01111100_01000110_1;
      patterns[51839] = 25'b11001010_01111101_01000111_1;
      patterns[51840] = 25'b11001010_01111110_01001000_1;
      patterns[51841] = 25'b11001010_01111111_01001001_1;
      patterns[51842] = 25'b11001010_10000000_01001010_1;
      patterns[51843] = 25'b11001010_10000001_01001011_1;
      patterns[51844] = 25'b11001010_10000010_01001100_1;
      patterns[51845] = 25'b11001010_10000011_01001101_1;
      patterns[51846] = 25'b11001010_10000100_01001110_1;
      patterns[51847] = 25'b11001010_10000101_01001111_1;
      patterns[51848] = 25'b11001010_10000110_01010000_1;
      patterns[51849] = 25'b11001010_10000111_01010001_1;
      patterns[51850] = 25'b11001010_10001000_01010010_1;
      patterns[51851] = 25'b11001010_10001001_01010011_1;
      patterns[51852] = 25'b11001010_10001010_01010100_1;
      patterns[51853] = 25'b11001010_10001011_01010101_1;
      patterns[51854] = 25'b11001010_10001100_01010110_1;
      patterns[51855] = 25'b11001010_10001101_01010111_1;
      patterns[51856] = 25'b11001010_10001110_01011000_1;
      patterns[51857] = 25'b11001010_10001111_01011001_1;
      patterns[51858] = 25'b11001010_10010000_01011010_1;
      patterns[51859] = 25'b11001010_10010001_01011011_1;
      patterns[51860] = 25'b11001010_10010010_01011100_1;
      patterns[51861] = 25'b11001010_10010011_01011101_1;
      patterns[51862] = 25'b11001010_10010100_01011110_1;
      patterns[51863] = 25'b11001010_10010101_01011111_1;
      patterns[51864] = 25'b11001010_10010110_01100000_1;
      patterns[51865] = 25'b11001010_10010111_01100001_1;
      patterns[51866] = 25'b11001010_10011000_01100010_1;
      patterns[51867] = 25'b11001010_10011001_01100011_1;
      patterns[51868] = 25'b11001010_10011010_01100100_1;
      patterns[51869] = 25'b11001010_10011011_01100101_1;
      patterns[51870] = 25'b11001010_10011100_01100110_1;
      patterns[51871] = 25'b11001010_10011101_01100111_1;
      patterns[51872] = 25'b11001010_10011110_01101000_1;
      patterns[51873] = 25'b11001010_10011111_01101001_1;
      patterns[51874] = 25'b11001010_10100000_01101010_1;
      patterns[51875] = 25'b11001010_10100001_01101011_1;
      patterns[51876] = 25'b11001010_10100010_01101100_1;
      patterns[51877] = 25'b11001010_10100011_01101101_1;
      patterns[51878] = 25'b11001010_10100100_01101110_1;
      patterns[51879] = 25'b11001010_10100101_01101111_1;
      patterns[51880] = 25'b11001010_10100110_01110000_1;
      patterns[51881] = 25'b11001010_10100111_01110001_1;
      patterns[51882] = 25'b11001010_10101000_01110010_1;
      patterns[51883] = 25'b11001010_10101001_01110011_1;
      patterns[51884] = 25'b11001010_10101010_01110100_1;
      patterns[51885] = 25'b11001010_10101011_01110101_1;
      patterns[51886] = 25'b11001010_10101100_01110110_1;
      patterns[51887] = 25'b11001010_10101101_01110111_1;
      patterns[51888] = 25'b11001010_10101110_01111000_1;
      patterns[51889] = 25'b11001010_10101111_01111001_1;
      patterns[51890] = 25'b11001010_10110000_01111010_1;
      patterns[51891] = 25'b11001010_10110001_01111011_1;
      patterns[51892] = 25'b11001010_10110010_01111100_1;
      patterns[51893] = 25'b11001010_10110011_01111101_1;
      patterns[51894] = 25'b11001010_10110100_01111110_1;
      patterns[51895] = 25'b11001010_10110101_01111111_1;
      patterns[51896] = 25'b11001010_10110110_10000000_1;
      patterns[51897] = 25'b11001010_10110111_10000001_1;
      patterns[51898] = 25'b11001010_10111000_10000010_1;
      patterns[51899] = 25'b11001010_10111001_10000011_1;
      patterns[51900] = 25'b11001010_10111010_10000100_1;
      patterns[51901] = 25'b11001010_10111011_10000101_1;
      patterns[51902] = 25'b11001010_10111100_10000110_1;
      patterns[51903] = 25'b11001010_10111101_10000111_1;
      patterns[51904] = 25'b11001010_10111110_10001000_1;
      patterns[51905] = 25'b11001010_10111111_10001001_1;
      patterns[51906] = 25'b11001010_11000000_10001010_1;
      patterns[51907] = 25'b11001010_11000001_10001011_1;
      patterns[51908] = 25'b11001010_11000010_10001100_1;
      patterns[51909] = 25'b11001010_11000011_10001101_1;
      patterns[51910] = 25'b11001010_11000100_10001110_1;
      patterns[51911] = 25'b11001010_11000101_10001111_1;
      patterns[51912] = 25'b11001010_11000110_10010000_1;
      patterns[51913] = 25'b11001010_11000111_10010001_1;
      patterns[51914] = 25'b11001010_11001000_10010010_1;
      patterns[51915] = 25'b11001010_11001001_10010011_1;
      patterns[51916] = 25'b11001010_11001010_10010100_1;
      patterns[51917] = 25'b11001010_11001011_10010101_1;
      patterns[51918] = 25'b11001010_11001100_10010110_1;
      patterns[51919] = 25'b11001010_11001101_10010111_1;
      patterns[51920] = 25'b11001010_11001110_10011000_1;
      patterns[51921] = 25'b11001010_11001111_10011001_1;
      patterns[51922] = 25'b11001010_11010000_10011010_1;
      patterns[51923] = 25'b11001010_11010001_10011011_1;
      patterns[51924] = 25'b11001010_11010010_10011100_1;
      patterns[51925] = 25'b11001010_11010011_10011101_1;
      patterns[51926] = 25'b11001010_11010100_10011110_1;
      patterns[51927] = 25'b11001010_11010101_10011111_1;
      patterns[51928] = 25'b11001010_11010110_10100000_1;
      patterns[51929] = 25'b11001010_11010111_10100001_1;
      patterns[51930] = 25'b11001010_11011000_10100010_1;
      patterns[51931] = 25'b11001010_11011001_10100011_1;
      patterns[51932] = 25'b11001010_11011010_10100100_1;
      patterns[51933] = 25'b11001010_11011011_10100101_1;
      patterns[51934] = 25'b11001010_11011100_10100110_1;
      patterns[51935] = 25'b11001010_11011101_10100111_1;
      patterns[51936] = 25'b11001010_11011110_10101000_1;
      patterns[51937] = 25'b11001010_11011111_10101001_1;
      patterns[51938] = 25'b11001010_11100000_10101010_1;
      patterns[51939] = 25'b11001010_11100001_10101011_1;
      patterns[51940] = 25'b11001010_11100010_10101100_1;
      patterns[51941] = 25'b11001010_11100011_10101101_1;
      patterns[51942] = 25'b11001010_11100100_10101110_1;
      patterns[51943] = 25'b11001010_11100101_10101111_1;
      patterns[51944] = 25'b11001010_11100110_10110000_1;
      patterns[51945] = 25'b11001010_11100111_10110001_1;
      patterns[51946] = 25'b11001010_11101000_10110010_1;
      patterns[51947] = 25'b11001010_11101001_10110011_1;
      patterns[51948] = 25'b11001010_11101010_10110100_1;
      patterns[51949] = 25'b11001010_11101011_10110101_1;
      patterns[51950] = 25'b11001010_11101100_10110110_1;
      patterns[51951] = 25'b11001010_11101101_10110111_1;
      patterns[51952] = 25'b11001010_11101110_10111000_1;
      patterns[51953] = 25'b11001010_11101111_10111001_1;
      patterns[51954] = 25'b11001010_11110000_10111010_1;
      patterns[51955] = 25'b11001010_11110001_10111011_1;
      patterns[51956] = 25'b11001010_11110010_10111100_1;
      patterns[51957] = 25'b11001010_11110011_10111101_1;
      patterns[51958] = 25'b11001010_11110100_10111110_1;
      patterns[51959] = 25'b11001010_11110101_10111111_1;
      patterns[51960] = 25'b11001010_11110110_11000000_1;
      patterns[51961] = 25'b11001010_11110111_11000001_1;
      patterns[51962] = 25'b11001010_11111000_11000010_1;
      patterns[51963] = 25'b11001010_11111001_11000011_1;
      patterns[51964] = 25'b11001010_11111010_11000100_1;
      patterns[51965] = 25'b11001010_11111011_11000101_1;
      patterns[51966] = 25'b11001010_11111100_11000110_1;
      patterns[51967] = 25'b11001010_11111101_11000111_1;
      patterns[51968] = 25'b11001010_11111110_11001000_1;
      patterns[51969] = 25'b11001010_11111111_11001001_1;
      patterns[51970] = 25'b11001011_00000000_11001011_0;
      patterns[51971] = 25'b11001011_00000001_11001100_0;
      patterns[51972] = 25'b11001011_00000010_11001101_0;
      patterns[51973] = 25'b11001011_00000011_11001110_0;
      patterns[51974] = 25'b11001011_00000100_11001111_0;
      patterns[51975] = 25'b11001011_00000101_11010000_0;
      patterns[51976] = 25'b11001011_00000110_11010001_0;
      patterns[51977] = 25'b11001011_00000111_11010010_0;
      patterns[51978] = 25'b11001011_00001000_11010011_0;
      patterns[51979] = 25'b11001011_00001001_11010100_0;
      patterns[51980] = 25'b11001011_00001010_11010101_0;
      patterns[51981] = 25'b11001011_00001011_11010110_0;
      patterns[51982] = 25'b11001011_00001100_11010111_0;
      patterns[51983] = 25'b11001011_00001101_11011000_0;
      patterns[51984] = 25'b11001011_00001110_11011001_0;
      patterns[51985] = 25'b11001011_00001111_11011010_0;
      patterns[51986] = 25'b11001011_00010000_11011011_0;
      patterns[51987] = 25'b11001011_00010001_11011100_0;
      patterns[51988] = 25'b11001011_00010010_11011101_0;
      patterns[51989] = 25'b11001011_00010011_11011110_0;
      patterns[51990] = 25'b11001011_00010100_11011111_0;
      patterns[51991] = 25'b11001011_00010101_11100000_0;
      patterns[51992] = 25'b11001011_00010110_11100001_0;
      patterns[51993] = 25'b11001011_00010111_11100010_0;
      patterns[51994] = 25'b11001011_00011000_11100011_0;
      patterns[51995] = 25'b11001011_00011001_11100100_0;
      patterns[51996] = 25'b11001011_00011010_11100101_0;
      patterns[51997] = 25'b11001011_00011011_11100110_0;
      patterns[51998] = 25'b11001011_00011100_11100111_0;
      patterns[51999] = 25'b11001011_00011101_11101000_0;
      patterns[52000] = 25'b11001011_00011110_11101001_0;
      patterns[52001] = 25'b11001011_00011111_11101010_0;
      patterns[52002] = 25'b11001011_00100000_11101011_0;
      patterns[52003] = 25'b11001011_00100001_11101100_0;
      patterns[52004] = 25'b11001011_00100010_11101101_0;
      patterns[52005] = 25'b11001011_00100011_11101110_0;
      patterns[52006] = 25'b11001011_00100100_11101111_0;
      patterns[52007] = 25'b11001011_00100101_11110000_0;
      patterns[52008] = 25'b11001011_00100110_11110001_0;
      patterns[52009] = 25'b11001011_00100111_11110010_0;
      patterns[52010] = 25'b11001011_00101000_11110011_0;
      patterns[52011] = 25'b11001011_00101001_11110100_0;
      patterns[52012] = 25'b11001011_00101010_11110101_0;
      patterns[52013] = 25'b11001011_00101011_11110110_0;
      patterns[52014] = 25'b11001011_00101100_11110111_0;
      patterns[52015] = 25'b11001011_00101101_11111000_0;
      patterns[52016] = 25'b11001011_00101110_11111001_0;
      patterns[52017] = 25'b11001011_00101111_11111010_0;
      patterns[52018] = 25'b11001011_00110000_11111011_0;
      patterns[52019] = 25'b11001011_00110001_11111100_0;
      patterns[52020] = 25'b11001011_00110010_11111101_0;
      patterns[52021] = 25'b11001011_00110011_11111110_0;
      patterns[52022] = 25'b11001011_00110100_11111111_0;
      patterns[52023] = 25'b11001011_00110101_00000000_1;
      patterns[52024] = 25'b11001011_00110110_00000001_1;
      patterns[52025] = 25'b11001011_00110111_00000010_1;
      patterns[52026] = 25'b11001011_00111000_00000011_1;
      patterns[52027] = 25'b11001011_00111001_00000100_1;
      patterns[52028] = 25'b11001011_00111010_00000101_1;
      patterns[52029] = 25'b11001011_00111011_00000110_1;
      patterns[52030] = 25'b11001011_00111100_00000111_1;
      patterns[52031] = 25'b11001011_00111101_00001000_1;
      patterns[52032] = 25'b11001011_00111110_00001001_1;
      patterns[52033] = 25'b11001011_00111111_00001010_1;
      patterns[52034] = 25'b11001011_01000000_00001011_1;
      patterns[52035] = 25'b11001011_01000001_00001100_1;
      patterns[52036] = 25'b11001011_01000010_00001101_1;
      patterns[52037] = 25'b11001011_01000011_00001110_1;
      patterns[52038] = 25'b11001011_01000100_00001111_1;
      patterns[52039] = 25'b11001011_01000101_00010000_1;
      patterns[52040] = 25'b11001011_01000110_00010001_1;
      patterns[52041] = 25'b11001011_01000111_00010010_1;
      patterns[52042] = 25'b11001011_01001000_00010011_1;
      patterns[52043] = 25'b11001011_01001001_00010100_1;
      patterns[52044] = 25'b11001011_01001010_00010101_1;
      patterns[52045] = 25'b11001011_01001011_00010110_1;
      patterns[52046] = 25'b11001011_01001100_00010111_1;
      patterns[52047] = 25'b11001011_01001101_00011000_1;
      patterns[52048] = 25'b11001011_01001110_00011001_1;
      patterns[52049] = 25'b11001011_01001111_00011010_1;
      patterns[52050] = 25'b11001011_01010000_00011011_1;
      patterns[52051] = 25'b11001011_01010001_00011100_1;
      patterns[52052] = 25'b11001011_01010010_00011101_1;
      patterns[52053] = 25'b11001011_01010011_00011110_1;
      patterns[52054] = 25'b11001011_01010100_00011111_1;
      patterns[52055] = 25'b11001011_01010101_00100000_1;
      patterns[52056] = 25'b11001011_01010110_00100001_1;
      patterns[52057] = 25'b11001011_01010111_00100010_1;
      patterns[52058] = 25'b11001011_01011000_00100011_1;
      patterns[52059] = 25'b11001011_01011001_00100100_1;
      patterns[52060] = 25'b11001011_01011010_00100101_1;
      patterns[52061] = 25'b11001011_01011011_00100110_1;
      patterns[52062] = 25'b11001011_01011100_00100111_1;
      patterns[52063] = 25'b11001011_01011101_00101000_1;
      patterns[52064] = 25'b11001011_01011110_00101001_1;
      patterns[52065] = 25'b11001011_01011111_00101010_1;
      patterns[52066] = 25'b11001011_01100000_00101011_1;
      patterns[52067] = 25'b11001011_01100001_00101100_1;
      patterns[52068] = 25'b11001011_01100010_00101101_1;
      patterns[52069] = 25'b11001011_01100011_00101110_1;
      patterns[52070] = 25'b11001011_01100100_00101111_1;
      patterns[52071] = 25'b11001011_01100101_00110000_1;
      patterns[52072] = 25'b11001011_01100110_00110001_1;
      patterns[52073] = 25'b11001011_01100111_00110010_1;
      patterns[52074] = 25'b11001011_01101000_00110011_1;
      patterns[52075] = 25'b11001011_01101001_00110100_1;
      patterns[52076] = 25'b11001011_01101010_00110101_1;
      patterns[52077] = 25'b11001011_01101011_00110110_1;
      patterns[52078] = 25'b11001011_01101100_00110111_1;
      patterns[52079] = 25'b11001011_01101101_00111000_1;
      patterns[52080] = 25'b11001011_01101110_00111001_1;
      patterns[52081] = 25'b11001011_01101111_00111010_1;
      patterns[52082] = 25'b11001011_01110000_00111011_1;
      patterns[52083] = 25'b11001011_01110001_00111100_1;
      patterns[52084] = 25'b11001011_01110010_00111101_1;
      patterns[52085] = 25'b11001011_01110011_00111110_1;
      patterns[52086] = 25'b11001011_01110100_00111111_1;
      patterns[52087] = 25'b11001011_01110101_01000000_1;
      patterns[52088] = 25'b11001011_01110110_01000001_1;
      patterns[52089] = 25'b11001011_01110111_01000010_1;
      patterns[52090] = 25'b11001011_01111000_01000011_1;
      patterns[52091] = 25'b11001011_01111001_01000100_1;
      patterns[52092] = 25'b11001011_01111010_01000101_1;
      patterns[52093] = 25'b11001011_01111011_01000110_1;
      patterns[52094] = 25'b11001011_01111100_01000111_1;
      patterns[52095] = 25'b11001011_01111101_01001000_1;
      patterns[52096] = 25'b11001011_01111110_01001001_1;
      patterns[52097] = 25'b11001011_01111111_01001010_1;
      patterns[52098] = 25'b11001011_10000000_01001011_1;
      patterns[52099] = 25'b11001011_10000001_01001100_1;
      patterns[52100] = 25'b11001011_10000010_01001101_1;
      patterns[52101] = 25'b11001011_10000011_01001110_1;
      patterns[52102] = 25'b11001011_10000100_01001111_1;
      patterns[52103] = 25'b11001011_10000101_01010000_1;
      patterns[52104] = 25'b11001011_10000110_01010001_1;
      patterns[52105] = 25'b11001011_10000111_01010010_1;
      patterns[52106] = 25'b11001011_10001000_01010011_1;
      patterns[52107] = 25'b11001011_10001001_01010100_1;
      patterns[52108] = 25'b11001011_10001010_01010101_1;
      patterns[52109] = 25'b11001011_10001011_01010110_1;
      patterns[52110] = 25'b11001011_10001100_01010111_1;
      patterns[52111] = 25'b11001011_10001101_01011000_1;
      patterns[52112] = 25'b11001011_10001110_01011001_1;
      patterns[52113] = 25'b11001011_10001111_01011010_1;
      patterns[52114] = 25'b11001011_10010000_01011011_1;
      patterns[52115] = 25'b11001011_10010001_01011100_1;
      patterns[52116] = 25'b11001011_10010010_01011101_1;
      patterns[52117] = 25'b11001011_10010011_01011110_1;
      patterns[52118] = 25'b11001011_10010100_01011111_1;
      patterns[52119] = 25'b11001011_10010101_01100000_1;
      patterns[52120] = 25'b11001011_10010110_01100001_1;
      patterns[52121] = 25'b11001011_10010111_01100010_1;
      patterns[52122] = 25'b11001011_10011000_01100011_1;
      patterns[52123] = 25'b11001011_10011001_01100100_1;
      patterns[52124] = 25'b11001011_10011010_01100101_1;
      patterns[52125] = 25'b11001011_10011011_01100110_1;
      patterns[52126] = 25'b11001011_10011100_01100111_1;
      patterns[52127] = 25'b11001011_10011101_01101000_1;
      patterns[52128] = 25'b11001011_10011110_01101001_1;
      patterns[52129] = 25'b11001011_10011111_01101010_1;
      patterns[52130] = 25'b11001011_10100000_01101011_1;
      patterns[52131] = 25'b11001011_10100001_01101100_1;
      patterns[52132] = 25'b11001011_10100010_01101101_1;
      patterns[52133] = 25'b11001011_10100011_01101110_1;
      patterns[52134] = 25'b11001011_10100100_01101111_1;
      patterns[52135] = 25'b11001011_10100101_01110000_1;
      patterns[52136] = 25'b11001011_10100110_01110001_1;
      patterns[52137] = 25'b11001011_10100111_01110010_1;
      patterns[52138] = 25'b11001011_10101000_01110011_1;
      patterns[52139] = 25'b11001011_10101001_01110100_1;
      patterns[52140] = 25'b11001011_10101010_01110101_1;
      patterns[52141] = 25'b11001011_10101011_01110110_1;
      patterns[52142] = 25'b11001011_10101100_01110111_1;
      patterns[52143] = 25'b11001011_10101101_01111000_1;
      patterns[52144] = 25'b11001011_10101110_01111001_1;
      patterns[52145] = 25'b11001011_10101111_01111010_1;
      patterns[52146] = 25'b11001011_10110000_01111011_1;
      patterns[52147] = 25'b11001011_10110001_01111100_1;
      patterns[52148] = 25'b11001011_10110010_01111101_1;
      patterns[52149] = 25'b11001011_10110011_01111110_1;
      patterns[52150] = 25'b11001011_10110100_01111111_1;
      patterns[52151] = 25'b11001011_10110101_10000000_1;
      patterns[52152] = 25'b11001011_10110110_10000001_1;
      patterns[52153] = 25'b11001011_10110111_10000010_1;
      patterns[52154] = 25'b11001011_10111000_10000011_1;
      patterns[52155] = 25'b11001011_10111001_10000100_1;
      patterns[52156] = 25'b11001011_10111010_10000101_1;
      patterns[52157] = 25'b11001011_10111011_10000110_1;
      patterns[52158] = 25'b11001011_10111100_10000111_1;
      patterns[52159] = 25'b11001011_10111101_10001000_1;
      patterns[52160] = 25'b11001011_10111110_10001001_1;
      patterns[52161] = 25'b11001011_10111111_10001010_1;
      patterns[52162] = 25'b11001011_11000000_10001011_1;
      patterns[52163] = 25'b11001011_11000001_10001100_1;
      patterns[52164] = 25'b11001011_11000010_10001101_1;
      patterns[52165] = 25'b11001011_11000011_10001110_1;
      patterns[52166] = 25'b11001011_11000100_10001111_1;
      patterns[52167] = 25'b11001011_11000101_10010000_1;
      patterns[52168] = 25'b11001011_11000110_10010001_1;
      patterns[52169] = 25'b11001011_11000111_10010010_1;
      patterns[52170] = 25'b11001011_11001000_10010011_1;
      patterns[52171] = 25'b11001011_11001001_10010100_1;
      patterns[52172] = 25'b11001011_11001010_10010101_1;
      patterns[52173] = 25'b11001011_11001011_10010110_1;
      patterns[52174] = 25'b11001011_11001100_10010111_1;
      patterns[52175] = 25'b11001011_11001101_10011000_1;
      patterns[52176] = 25'b11001011_11001110_10011001_1;
      patterns[52177] = 25'b11001011_11001111_10011010_1;
      patterns[52178] = 25'b11001011_11010000_10011011_1;
      patterns[52179] = 25'b11001011_11010001_10011100_1;
      patterns[52180] = 25'b11001011_11010010_10011101_1;
      patterns[52181] = 25'b11001011_11010011_10011110_1;
      patterns[52182] = 25'b11001011_11010100_10011111_1;
      patterns[52183] = 25'b11001011_11010101_10100000_1;
      patterns[52184] = 25'b11001011_11010110_10100001_1;
      patterns[52185] = 25'b11001011_11010111_10100010_1;
      patterns[52186] = 25'b11001011_11011000_10100011_1;
      patterns[52187] = 25'b11001011_11011001_10100100_1;
      patterns[52188] = 25'b11001011_11011010_10100101_1;
      patterns[52189] = 25'b11001011_11011011_10100110_1;
      patterns[52190] = 25'b11001011_11011100_10100111_1;
      patterns[52191] = 25'b11001011_11011101_10101000_1;
      patterns[52192] = 25'b11001011_11011110_10101001_1;
      patterns[52193] = 25'b11001011_11011111_10101010_1;
      patterns[52194] = 25'b11001011_11100000_10101011_1;
      patterns[52195] = 25'b11001011_11100001_10101100_1;
      patterns[52196] = 25'b11001011_11100010_10101101_1;
      patterns[52197] = 25'b11001011_11100011_10101110_1;
      patterns[52198] = 25'b11001011_11100100_10101111_1;
      patterns[52199] = 25'b11001011_11100101_10110000_1;
      patterns[52200] = 25'b11001011_11100110_10110001_1;
      patterns[52201] = 25'b11001011_11100111_10110010_1;
      patterns[52202] = 25'b11001011_11101000_10110011_1;
      patterns[52203] = 25'b11001011_11101001_10110100_1;
      patterns[52204] = 25'b11001011_11101010_10110101_1;
      patterns[52205] = 25'b11001011_11101011_10110110_1;
      patterns[52206] = 25'b11001011_11101100_10110111_1;
      patterns[52207] = 25'b11001011_11101101_10111000_1;
      patterns[52208] = 25'b11001011_11101110_10111001_1;
      patterns[52209] = 25'b11001011_11101111_10111010_1;
      patterns[52210] = 25'b11001011_11110000_10111011_1;
      patterns[52211] = 25'b11001011_11110001_10111100_1;
      patterns[52212] = 25'b11001011_11110010_10111101_1;
      patterns[52213] = 25'b11001011_11110011_10111110_1;
      patterns[52214] = 25'b11001011_11110100_10111111_1;
      patterns[52215] = 25'b11001011_11110101_11000000_1;
      patterns[52216] = 25'b11001011_11110110_11000001_1;
      patterns[52217] = 25'b11001011_11110111_11000010_1;
      patterns[52218] = 25'b11001011_11111000_11000011_1;
      patterns[52219] = 25'b11001011_11111001_11000100_1;
      patterns[52220] = 25'b11001011_11111010_11000101_1;
      patterns[52221] = 25'b11001011_11111011_11000110_1;
      patterns[52222] = 25'b11001011_11111100_11000111_1;
      patterns[52223] = 25'b11001011_11111101_11001000_1;
      patterns[52224] = 25'b11001011_11111110_11001001_1;
      patterns[52225] = 25'b11001011_11111111_11001010_1;
      patterns[52226] = 25'b11001100_00000000_11001100_0;
      patterns[52227] = 25'b11001100_00000001_11001101_0;
      patterns[52228] = 25'b11001100_00000010_11001110_0;
      patterns[52229] = 25'b11001100_00000011_11001111_0;
      patterns[52230] = 25'b11001100_00000100_11010000_0;
      patterns[52231] = 25'b11001100_00000101_11010001_0;
      patterns[52232] = 25'b11001100_00000110_11010010_0;
      patterns[52233] = 25'b11001100_00000111_11010011_0;
      patterns[52234] = 25'b11001100_00001000_11010100_0;
      patterns[52235] = 25'b11001100_00001001_11010101_0;
      patterns[52236] = 25'b11001100_00001010_11010110_0;
      patterns[52237] = 25'b11001100_00001011_11010111_0;
      patterns[52238] = 25'b11001100_00001100_11011000_0;
      patterns[52239] = 25'b11001100_00001101_11011001_0;
      patterns[52240] = 25'b11001100_00001110_11011010_0;
      patterns[52241] = 25'b11001100_00001111_11011011_0;
      patterns[52242] = 25'b11001100_00010000_11011100_0;
      patterns[52243] = 25'b11001100_00010001_11011101_0;
      patterns[52244] = 25'b11001100_00010010_11011110_0;
      patterns[52245] = 25'b11001100_00010011_11011111_0;
      patterns[52246] = 25'b11001100_00010100_11100000_0;
      patterns[52247] = 25'b11001100_00010101_11100001_0;
      patterns[52248] = 25'b11001100_00010110_11100010_0;
      patterns[52249] = 25'b11001100_00010111_11100011_0;
      patterns[52250] = 25'b11001100_00011000_11100100_0;
      patterns[52251] = 25'b11001100_00011001_11100101_0;
      patterns[52252] = 25'b11001100_00011010_11100110_0;
      patterns[52253] = 25'b11001100_00011011_11100111_0;
      patterns[52254] = 25'b11001100_00011100_11101000_0;
      patterns[52255] = 25'b11001100_00011101_11101001_0;
      patterns[52256] = 25'b11001100_00011110_11101010_0;
      patterns[52257] = 25'b11001100_00011111_11101011_0;
      patterns[52258] = 25'b11001100_00100000_11101100_0;
      patterns[52259] = 25'b11001100_00100001_11101101_0;
      patterns[52260] = 25'b11001100_00100010_11101110_0;
      patterns[52261] = 25'b11001100_00100011_11101111_0;
      patterns[52262] = 25'b11001100_00100100_11110000_0;
      patterns[52263] = 25'b11001100_00100101_11110001_0;
      patterns[52264] = 25'b11001100_00100110_11110010_0;
      patterns[52265] = 25'b11001100_00100111_11110011_0;
      patterns[52266] = 25'b11001100_00101000_11110100_0;
      patterns[52267] = 25'b11001100_00101001_11110101_0;
      patterns[52268] = 25'b11001100_00101010_11110110_0;
      patterns[52269] = 25'b11001100_00101011_11110111_0;
      patterns[52270] = 25'b11001100_00101100_11111000_0;
      patterns[52271] = 25'b11001100_00101101_11111001_0;
      patterns[52272] = 25'b11001100_00101110_11111010_0;
      patterns[52273] = 25'b11001100_00101111_11111011_0;
      patterns[52274] = 25'b11001100_00110000_11111100_0;
      patterns[52275] = 25'b11001100_00110001_11111101_0;
      patterns[52276] = 25'b11001100_00110010_11111110_0;
      patterns[52277] = 25'b11001100_00110011_11111111_0;
      patterns[52278] = 25'b11001100_00110100_00000000_1;
      patterns[52279] = 25'b11001100_00110101_00000001_1;
      patterns[52280] = 25'b11001100_00110110_00000010_1;
      patterns[52281] = 25'b11001100_00110111_00000011_1;
      patterns[52282] = 25'b11001100_00111000_00000100_1;
      patterns[52283] = 25'b11001100_00111001_00000101_1;
      patterns[52284] = 25'b11001100_00111010_00000110_1;
      patterns[52285] = 25'b11001100_00111011_00000111_1;
      patterns[52286] = 25'b11001100_00111100_00001000_1;
      patterns[52287] = 25'b11001100_00111101_00001001_1;
      patterns[52288] = 25'b11001100_00111110_00001010_1;
      patterns[52289] = 25'b11001100_00111111_00001011_1;
      patterns[52290] = 25'b11001100_01000000_00001100_1;
      patterns[52291] = 25'b11001100_01000001_00001101_1;
      patterns[52292] = 25'b11001100_01000010_00001110_1;
      patterns[52293] = 25'b11001100_01000011_00001111_1;
      patterns[52294] = 25'b11001100_01000100_00010000_1;
      patterns[52295] = 25'b11001100_01000101_00010001_1;
      patterns[52296] = 25'b11001100_01000110_00010010_1;
      patterns[52297] = 25'b11001100_01000111_00010011_1;
      patterns[52298] = 25'b11001100_01001000_00010100_1;
      patterns[52299] = 25'b11001100_01001001_00010101_1;
      patterns[52300] = 25'b11001100_01001010_00010110_1;
      patterns[52301] = 25'b11001100_01001011_00010111_1;
      patterns[52302] = 25'b11001100_01001100_00011000_1;
      patterns[52303] = 25'b11001100_01001101_00011001_1;
      patterns[52304] = 25'b11001100_01001110_00011010_1;
      patterns[52305] = 25'b11001100_01001111_00011011_1;
      patterns[52306] = 25'b11001100_01010000_00011100_1;
      patterns[52307] = 25'b11001100_01010001_00011101_1;
      patterns[52308] = 25'b11001100_01010010_00011110_1;
      patterns[52309] = 25'b11001100_01010011_00011111_1;
      patterns[52310] = 25'b11001100_01010100_00100000_1;
      patterns[52311] = 25'b11001100_01010101_00100001_1;
      patterns[52312] = 25'b11001100_01010110_00100010_1;
      patterns[52313] = 25'b11001100_01010111_00100011_1;
      patterns[52314] = 25'b11001100_01011000_00100100_1;
      patterns[52315] = 25'b11001100_01011001_00100101_1;
      patterns[52316] = 25'b11001100_01011010_00100110_1;
      patterns[52317] = 25'b11001100_01011011_00100111_1;
      patterns[52318] = 25'b11001100_01011100_00101000_1;
      patterns[52319] = 25'b11001100_01011101_00101001_1;
      patterns[52320] = 25'b11001100_01011110_00101010_1;
      patterns[52321] = 25'b11001100_01011111_00101011_1;
      patterns[52322] = 25'b11001100_01100000_00101100_1;
      patterns[52323] = 25'b11001100_01100001_00101101_1;
      patterns[52324] = 25'b11001100_01100010_00101110_1;
      patterns[52325] = 25'b11001100_01100011_00101111_1;
      patterns[52326] = 25'b11001100_01100100_00110000_1;
      patterns[52327] = 25'b11001100_01100101_00110001_1;
      patterns[52328] = 25'b11001100_01100110_00110010_1;
      patterns[52329] = 25'b11001100_01100111_00110011_1;
      patterns[52330] = 25'b11001100_01101000_00110100_1;
      patterns[52331] = 25'b11001100_01101001_00110101_1;
      patterns[52332] = 25'b11001100_01101010_00110110_1;
      patterns[52333] = 25'b11001100_01101011_00110111_1;
      patterns[52334] = 25'b11001100_01101100_00111000_1;
      patterns[52335] = 25'b11001100_01101101_00111001_1;
      patterns[52336] = 25'b11001100_01101110_00111010_1;
      patterns[52337] = 25'b11001100_01101111_00111011_1;
      patterns[52338] = 25'b11001100_01110000_00111100_1;
      patterns[52339] = 25'b11001100_01110001_00111101_1;
      patterns[52340] = 25'b11001100_01110010_00111110_1;
      patterns[52341] = 25'b11001100_01110011_00111111_1;
      patterns[52342] = 25'b11001100_01110100_01000000_1;
      patterns[52343] = 25'b11001100_01110101_01000001_1;
      patterns[52344] = 25'b11001100_01110110_01000010_1;
      patterns[52345] = 25'b11001100_01110111_01000011_1;
      patterns[52346] = 25'b11001100_01111000_01000100_1;
      patterns[52347] = 25'b11001100_01111001_01000101_1;
      patterns[52348] = 25'b11001100_01111010_01000110_1;
      patterns[52349] = 25'b11001100_01111011_01000111_1;
      patterns[52350] = 25'b11001100_01111100_01001000_1;
      patterns[52351] = 25'b11001100_01111101_01001001_1;
      patterns[52352] = 25'b11001100_01111110_01001010_1;
      patterns[52353] = 25'b11001100_01111111_01001011_1;
      patterns[52354] = 25'b11001100_10000000_01001100_1;
      patterns[52355] = 25'b11001100_10000001_01001101_1;
      patterns[52356] = 25'b11001100_10000010_01001110_1;
      patterns[52357] = 25'b11001100_10000011_01001111_1;
      patterns[52358] = 25'b11001100_10000100_01010000_1;
      patterns[52359] = 25'b11001100_10000101_01010001_1;
      patterns[52360] = 25'b11001100_10000110_01010010_1;
      patterns[52361] = 25'b11001100_10000111_01010011_1;
      patterns[52362] = 25'b11001100_10001000_01010100_1;
      patterns[52363] = 25'b11001100_10001001_01010101_1;
      patterns[52364] = 25'b11001100_10001010_01010110_1;
      patterns[52365] = 25'b11001100_10001011_01010111_1;
      patterns[52366] = 25'b11001100_10001100_01011000_1;
      patterns[52367] = 25'b11001100_10001101_01011001_1;
      patterns[52368] = 25'b11001100_10001110_01011010_1;
      patterns[52369] = 25'b11001100_10001111_01011011_1;
      patterns[52370] = 25'b11001100_10010000_01011100_1;
      patterns[52371] = 25'b11001100_10010001_01011101_1;
      patterns[52372] = 25'b11001100_10010010_01011110_1;
      patterns[52373] = 25'b11001100_10010011_01011111_1;
      patterns[52374] = 25'b11001100_10010100_01100000_1;
      patterns[52375] = 25'b11001100_10010101_01100001_1;
      patterns[52376] = 25'b11001100_10010110_01100010_1;
      patterns[52377] = 25'b11001100_10010111_01100011_1;
      patterns[52378] = 25'b11001100_10011000_01100100_1;
      patterns[52379] = 25'b11001100_10011001_01100101_1;
      patterns[52380] = 25'b11001100_10011010_01100110_1;
      patterns[52381] = 25'b11001100_10011011_01100111_1;
      patterns[52382] = 25'b11001100_10011100_01101000_1;
      patterns[52383] = 25'b11001100_10011101_01101001_1;
      patterns[52384] = 25'b11001100_10011110_01101010_1;
      patterns[52385] = 25'b11001100_10011111_01101011_1;
      patterns[52386] = 25'b11001100_10100000_01101100_1;
      patterns[52387] = 25'b11001100_10100001_01101101_1;
      patterns[52388] = 25'b11001100_10100010_01101110_1;
      patterns[52389] = 25'b11001100_10100011_01101111_1;
      patterns[52390] = 25'b11001100_10100100_01110000_1;
      patterns[52391] = 25'b11001100_10100101_01110001_1;
      patterns[52392] = 25'b11001100_10100110_01110010_1;
      patterns[52393] = 25'b11001100_10100111_01110011_1;
      patterns[52394] = 25'b11001100_10101000_01110100_1;
      patterns[52395] = 25'b11001100_10101001_01110101_1;
      patterns[52396] = 25'b11001100_10101010_01110110_1;
      patterns[52397] = 25'b11001100_10101011_01110111_1;
      patterns[52398] = 25'b11001100_10101100_01111000_1;
      patterns[52399] = 25'b11001100_10101101_01111001_1;
      patterns[52400] = 25'b11001100_10101110_01111010_1;
      patterns[52401] = 25'b11001100_10101111_01111011_1;
      patterns[52402] = 25'b11001100_10110000_01111100_1;
      patterns[52403] = 25'b11001100_10110001_01111101_1;
      patterns[52404] = 25'b11001100_10110010_01111110_1;
      patterns[52405] = 25'b11001100_10110011_01111111_1;
      patterns[52406] = 25'b11001100_10110100_10000000_1;
      patterns[52407] = 25'b11001100_10110101_10000001_1;
      patterns[52408] = 25'b11001100_10110110_10000010_1;
      patterns[52409] = 25'b11001100_10110111_10000011_1;
      patterns[52410] = 25'b11001100_10111000_10000100_1;
      patterns[52411] = 25'b11001100_10111001_10000101_1;
      patterns[52412] = 25'b11001100_10111010_10000110_1;
      patterns[52413] = 25'b11001100_10111011_10000111_1;
      patterns[52414] = 25'b11001100_10111100_10001000_1;
      patterns[52415] = 25'b11001100_10111101_10001001_1;
      patterns[52416] = 25'b11001100_10111110_10001010_1;
      patterns[52417] = 25'b11001100_10111111_10001011_1;
      patterns[52418] = 25'b11001100_11000000_10001100_1;
      patterns[52419] = 25'b11001100_11000001_10001101_1;
      patterns[52420] = 25'b11001100_11000010_10001110_1;
      patterns[52421] = 25'b11001100_11000011_10001111_1;
      patterns[52422] = 25'b11001100_11000100_10010000_1;
      patterns[52423] = 25'b11001100_11000101_10010001_1;
      patterns[52424] = 25'b11001100_11000110_10010010_1;
      patterns[52425] = 25'b11001100_11000111_10010011_1;
      patterns[52426] = 25'b11001100_11001000_10010100_1;
      patterns[52427] = 25'b11001100_11001001_10010101_1;
      patterns[52428] = 25'b11001100_11001010_10010110_1;
      patterns[52429] = 25'b11001100_11001011_10010111_1;
      patterns[52430] = 25'b11001100_11001100_10011000_1;
      patterns[52431] = 25'b11001100_11001101_10011001_1;
      patterns[52432] = 25'b11001100_11001110_10011010_1;
      patterns[52433] = 25'b11001100_11001111_10011011_1;
      patterns[52434] = 25'b11001100_11010000_10011100_1;
      patterns[52435] = 25'b11001100_11010001_10011101_1;
      patterns[52436] = 25'b11001100_11010010_10011110_1;
      patterns[52437] = 25'b11001100_11010011_10011111_1;
      patterns[52438] = 25'b11001100_11010100_10100000_1;
      patterns[52439] = 25'b11001100_11010101_10100001_1;
      patterns[52440] = 25'b11001100_11010110_10100010_1;
      patterns[52441] = 25'b11001100_11010111_10100011_1;
      patterns[52442] = 25'b11001100_11011000_10100100_1;
      patterns[52443] = 25'b11001100_11011001_10100101_1;
      patterns[52444] = 25'b11001100_11011010_10100110_1;
      patterns[52445] = 25'b11001100_11011011_10100111_1;
      patterns[52446] = 25'b11001100_11011100_10101000_1;
      patterns[52447] = 25'b11001100_11011101_10101001_1;
      patterns[52448] = 25'b11001100_11011110_10101010_1;
      patterns[52449] = 25'b11001100_11011111_10101011_1;
      patterns[52450] = 25'b11001100_11100000_10101100_1;
      patterns[52451] = 25'b11001100_11100001_10101101_1;
      patterns[52452] = 25'b11001100_11100010_10101110_1;
      patterns[52453] = 25'b11001100_11100011_10101111_1;
      patterns[52454] = 25'b11001100_11100100_10110000_1;
      patterns[52455] = 25'b11001100_11100101_10110001_1;
      patterns[52456] = 25'b11001100_11100110_10110010_1;
      patterns[52457] = 25'b11001100_11100111_10110011_1;
      patterns[52458] = 25'b11001100_11101000_10110100_1;
      patterns[52459] = 25'b11001100_11101001_10110101_1;
      patterns[52460] = 25'b11001100_11101010_10110110_1;
      patterns[52461] = 25'b11001100_11101011_10110111_1;
      patterns[52462] = 25'b11001100_11101100_10111000_1;
      patterns[52463] = 25'b11001100_11101101_10111001_1;
      patterns[52464] = 25'b11001100_11101110_10111010_1;
      patterns[52465] = 25'b11001100_11101111_10111011_1;
      patterns[52466] = 25'b11001100_11110000_10111100_1;
      patterns[52467] = 25'b11001100_11110001_10111101_1;
      patterns[52468] = 25'b11001100_11110010_10111110_1;
      patterns[52469] = 25'b11001100_11110011_10111111_1;
      patterns[52470] = 25'b11001100_11110100_11000000_1;
      patterns[52471] = 25'b11001100_11110101_11000001_1;
      patterns[52472] = 25'b11001100_11110110_11000010_1;
      patterns[52473] = 25'b11001100_11110111_11000011_1;
      patterns[52474] = 25'b11001100_11111000_11000100_1;
      patterns[52475] = 25'b11001100_11111001_11000101_1;
      patterns[52476] = 25'b11001100_11111010_11000110_1;
      patterns[52477] = 25'b11001100_11111011_11000111_1;
      patterns[52478] = 25'b11001100_11111100_11001000_1;
      patterns[52479] = 25'b11001100_11111101_11001001_1;
      patterns[52480] = 25'b11001100_11111110_11001010_1;
      patterns[52481] = 25'b11001100_11111111_11001011_1;
      patterns[52482] = 25'b11001101_00000000_11001101_0;
      patterns[52483] = 25'b11001101_00000001_11001110_0;
      patterns[52484] = 25'b11001101_00000010_11001111_0;
      patterns[52485] = 25'b11001101_00000011_11010000_0;
      patterns[52486] = 25'b11001101_00000100_11010001_0;
      patterns[52487] = 25'b11001101_00000101_11010010_0;
      patterns[52488] = 25'b11001101_00000110_11010011_0;
      patterns[52489] = 25'b11001101_00000111_11010100_0;
      patterns[52490] = 25'b11001101_00001000_11010101_0;
      patterns[52491] = 25'b11001101_00001001_11010110_0;
      patterns[52492] = 25'b11001101_00001010_11010111_0;
      patterns[52493] = 25'b11001101_00001011_11011000_0;
      patterns[52494] = 25'b11001101_00001100_11011001_0;
      patterns[52495] = 25'b11001101_00001101_11011010_0;
      patterns[52496] = 25'b11001101_00001110_11011011_0;
      patterns[52497] = 25'b11001101_00001111_11011100_0;
      patterns[52498] = 25'b11001101_00010000_11011101_0;
      patterns[52499] = 25'b11001101_00010001_11011110_0;
      patterns[52500] = 25'b11001101_00010010_11011111_0;
      patterns[52501] = 25'b11001101_00010011_11100000_0;
      patterns[52502] = 25'b11001101_00010100_11100001_0;
      patterns[52503] = 25'b11001101_00010101_11100010_0;
      patterns[52504] = 25'b11001101_00010110_11100011_0;
      patterns[52505] = 25'b11001101_00010111_11100100_0;
      patterns[52506] = 25'b11001101_00011000_11100101_0;
      patterns[52507] = 25'b11001101_00011001_11100110_0;
      patterns[52508] = 25'b11001101_00011010_11100111_0;
      patterns[52509] = 25'b11001101_00011011_11101000_0;
      patterns[52510] = 25'b11001101_00011100_11101001_0;
      patterns[52511] = 25'b11001101_00011101_11101010_0;
      patterns[52512] = 25'b11001101_00011110_11101011_0;
      patterns[52513] = 25'b11001101_00011111_11101100_0;
      patterns[52514] = 25'b11001101_00100000_11101101_0;
      patterns[52515] = 25'b11001101_00100001_11101110_0;
      patterns[52516] = 25'b11001101_00100010_11101111_0;
      patterns[52517] = 25'b11001101_00100011_11110000_0;
      patterns[52518] = 25'b11001101_00100100_11110001_0;
      patterns[52519] = 25'b11001101_00100101_11110010_0;
      patterns[52520] = 25'b11001101_00100110_11110011_0;
      patterns[52521] = 25'b11001101_00100111_11110100_0;
      patterns[52522] = 25'b11001101_00101000_11110101_0;
      patterns[52523] = 25'b11001101_00101001_11110110_0;
      patterns[52524] = 25'b11001101_00101010_11110111_0;
      patterns[52525] = 25'b11001101_00101011_11111000_0;
      patterns[52526] = 25'b11001101_00101100_11111001_0;
      patterns[52527] = 25'b11001101_00101101_11111010_0;
      patterns[52528] = 25'b11001101_00101110_11111011_0;
      patterns[52529] = 25'b11001101_00101111_11111100_0;
      patterns[52530] = 25'b11001101_00110000_11111101_0;
      patterns[52531] = 25'b11001101_00110001_11111110_0;
      patterns[52532] = 25'b11001101_00110010_11111111_0;
      patterns[52533] = 25'b11001101_00110011_00000000_1;
      patterns[52534] = 25'b11001101_00110100_00000001_1;
      patterns[52535] = 25'b11001101_00110101_00000010_1;
      patterns[52536] = 25'b11001101_00110110_00000011_1;
      patterns[52537] = 25'b11001101_00110111_00000100_1;
      patterns[52538] = 25'b11001101_00111000_00000101_1;
      patterns[52539] = 25'b11001101_00111001_00000110_1;
      patterns[52540] = 25'b11001101_00111010_00000111_1;
      patterns[52541] = 25'b11001101_00111011_00001000_1;
      patterns[52542] = 25'b11001101_00111100_00001001_1;
      patterns[52543] = 25'b11001101_00111101_00001010_1;
      patterns[52544] = 25'b11001101_00111110_00001011_1;
      patterns[52545] = 25'b11001101_00111111_00001100_1;
      patterns[52546] = 25'b11001101_01000000_00001101_1;
      patterns[52547] = 25'b11001101_01000001_00001110_1;
      patterns[52548] = 25'b11001101_01000010_00001111_1;
      patterns[52549] = 25'b11001101_01000011_00010000_1;
      patterns[52550] = 25'b11001101_01000100_00010001_1;
      patterns[52551] = 25'b11001101_01000101_00010010_1;
      patterns[52552] = 25'b11001101_01000110_00010011_1;
      patterns[52553] = 25'b11001101_01000111_00010100_1;
      patterns[52554] = 25'b11001101_01001000_00010101_1;
      patterns[52555] = 25'b11001101_01001001_00010110_1;
      patterns[52556] = 25'b11001101_01001010_00010111_1;
      patterns[52557] = 25'b11001101_01001011_00011000_1;
      patterns[52558] = 25'b11001101_01001100_00011001_1;
      patterns[52559] = 25'b11001101_01001101_00011010_1;
      patterns[52560] = 25'b11001101_01001110_00011011_1;
      patterns[52561] = 25'b11001101_01001111_00011100_1;
      patterns[52562] = 25'b11001101_01010000_00011101_1;
      patterns[52563] = 25'b11001101_01010001_00011110_1;
      patterns[52564] = 25'b11001101_01010010_00011111_1;
      patterns[52565] = 25'b11001101_01010011_00100000_1;
      patterns[52566] = 25'b11001101_01010100_00100001_1;
      patterns[52567] = 25'b11001101_01010101_00100010_1;
      patterns[52568] = 25'b11001101_01010110_00100011_1;
      patterns[52569] = 25'b11001101_01010111_00100100_1;
      patterns[52570] = 25'b11001101_01011000_00100101_1;
      patterns[52571] = 25'b11001101_01011001_00100110_1;
      patterns[52572] = 25'b11001101_01011010_00100111_1;
      patterns[52573] = 25'b11001101_01011011_00101000_1;
      patterns[52574] = 25'b11001101_01011100_00101001_1;
      patterns[52575] = 25'b11001101_01011101_00101010_1;
      patterns[52576] = 25'b11001101_01011110_00101011_1;
      patterns[52577] = 25'b11001101_01011111_00101100_1;
      patterns[52578] = 25'b11001101_01100000_00101101_1;
      patterns[52579] = 25'b11001101_01100001_00101110_1;
      patterns[52580] = 25'b11001101_01100010_00101111_1;
      patterns[52581] = 25'b11001101_01100011_00110000_1;
      patterns[52582] = 25'b11001101_01100100_00110001_1;
      patterns[52583] = 25'b11001101_01100101_00110010_1;
      patterns[52584] = 25'b11001101_01100110_00110011_1;
      patterns[52585] = 25'b11001101_01100111_00110100_1;
      patterns[52586] = 25'b11001101_01101000_00110101_1;
      patterns[52587] = 25'b11001101_01101001_00110110_1;
      patterns[52588] = 25'b11001101_01101010_00110111_1;
      patterns[52589] = 25'b11001101_01101011_00111000_1;
      patterns[52590] = 25'b11001101_01101100_00111001_1;
      patterns[52591] = 25'b11001101_01101101_00111010_1;
      patterns[52592] = 25'b11001101_01101110_00111011_1;
      patterns[52593] = 25'b11001101_01101111_00111100_1;
      patterns[52594] = 25'b11001101_01110000_00111101_1;
      patterns[52595] = 25'b11001101_01110001_00111110_1;
      patterns[52596] = 25'b11001101_01110010_00111111_1;
      patterns[52597] = 25'b11001101_01110011_01000000_1;
      patterns[52598] = 25'b11001101_01110100_01000001_1;
      patterns[52599] = 25'b11001101_01110101_01000010_1;
      patterns[52600] = 25'b11001101_01110110_01000011_1;
      patterns[52601] = 25'b11001101_01110111_01000100_1;
      patterns[52602] = 25'b11001101_01111000_01000101_1;
      patterns[52603] = 25'b11001101_01111001_01000110_1;
      patterns[52604] = 25'b11001101_01111010_01000111_1;
      patterns[52605] = 25'b11001101_01111011_01001000_1;
      patterns[52606] = 25'b11001101_01111100_01001001_1;
      patterns[52607] = 25'b11001101_01111101_01001010_1;
      patterns[52608] = 25'b11001101_01111110_01001011_1;
      patterns[52609] = 25'b11001101_01111111_01001100_1;
      patterns[52610] = 25'b11001101_10000000_01001101_1;
      patterns[52611] = 25'b11001101_10000001_01001110_1;
      patterns[52612] = 25'b11001101_10000010_01001111_1;
      patterns[52613] = 25'b11001101_10000011_01010000_1;
      patterns[52614] = 25'b11001101_10000100_01010001_1;
      patterns[52615] = 25'b11001101_10000101_01010010_1;
      patterns[52616] = 25'b11001101_10000110_01010011_1;
      patterns[52617] = 25'b11001101_10000111_01010100_1;
      patterns[52618] = 25'b11001101_10001000_01010101_1;
      patterns[52619] = 25'b11001101_10001001_01010110_1;
      patterns[52620] = 25'b11001101_10001010_01010111_1;
      patterns[52621] = 25'b11001101_10001011_01011000_1;
      patterns[52622] = 25'b11001101_10001100_01011001_1;
      patterns[52623] = 25'b11001101_10001101_01011010_1;
      patterns[52624] = 25'b11001101_10001110_01011011_1;
      patterns[52625] = 25'b11001101_10001111_01011100_1;
      patterns[52626] = 25'b11001101_10010000_01011101_1;
      patterns[52627] = 25'b11001101_10010001_01011110_1;
      patterns[52628] = 25'b11001101_10010010_01011111_1;
      patterns[52629] = 25'b11001101_10010011_01100000_1;
      patterns[52630] = 25'b11001101_10010100_01100001_1;
      patterns[52631] = 25'b11001101_10010101_01100010_1;
      patterns[52632] = 25'b11001101_10010110_01100011_1;
      patterns[52633] = 25'b11001101_10010111_01100100_1;
      patterns[52634] = 25'b11001101_10011000_01100101_1;
      patterns[52635] = 25'b11001101_10011001_01100110_1;
      patterns[52636] = 25'b11001101_10011010_01100111_1;
      patterns[52637] = 25'b11001101_10011011_01101000_1;
      patterns[52638] = 25'b11001101_10011100_01101001_1;
      patterns[52639] = 25'b11001101_10011101_01101010_1;
      patterns[52640] = 25'b11001101_10011110_01101011_1;
      patterns[52641] = 25'b11001101_10011111_01101100_1;
      patterns[52642] = 25'b11001101_10100000_01101101_1;
      patterns[52643] = 25'b11001101_10100001_01101110_1;
      patterns[52644] = 25'b11001101_10100010_01101111_1;
      patterns[52645] = 25'b11001101_10100011_01110000_1;
      patterns[52646] = 25'b11001101_10100100_01110001_1;
      patterns[52647] = 25'b11001101_10100101_01110010_1;
      patterns[52648] = 25'b11001101_10100110_01110011_1;
      patterns[52649] = 25'b11001101_10100111_01110100_1;
      patterns[52650] = 25'b11001101_10101000_01110101_1;
      patterns[52651] = 25'b11001101_10101001_01110110_1;
      patterns[52652] = 25'b11001101_10101010_01110111_1;
      patterns[52653] = 25'b11001101_10101011_01111000_1;
      patterns[52654] = 25'b11001101_10101100_01111001_1;
      patterns[52655] = 25'b11001101_10101101_01111010_1;
      patterns[52656] = 25'b11001101_10101110_01111011_1;
      patterns[52657] = 25'b11001101_10101111_01111100_1;
      patterns[52658] = 25'b11001101_10110000_01111101_1;
      patterns[52659] = 25'b11001101_10110001_01111110_1;
      patterns[52660] = 25'b11001101_10110010_01111111_1;
      patterns[52661] = 25'b11001101_10110011_10000000_1;
      patterns[52662] = 25'b11001101_10110100_10000001_1;
      patterns[52663] = 25'b11001101_10110101_10000010_1;
      patterns[52664] = 25'b11001101_10110110_10000011_1;
      patterns[52665] = 25'b11001101_10110111_10000100_1;
      patterns[52666] = 25'b11001101_10111000_10000101_1;
      patterns[52667] = 25'b11001101_10111001_10000110_1;
      patterns[52668] = 25'b11001101_10111010_10000111_1;
      patterns[52669] = 25'b11001101_10111011_10001000_1;
      patterns[52670] = 25'b11001101_10111100_10001001_1;
      patterns[52671] = 25'b11001101_10111101_10001010_1;
      patterns[52672] = 25'b11001101_10111110_10001011_1;
      patterns[52673] = 25'b11001101_10111111_10001100_1;
      patterns[52674] = 25'b11001101_11000000_10001101_1;
      patterns[52675] = 25'b11001101_11000001_10001110_1;
      patterns[52676] = 25'b11001101_11000010_10001111_1;
      patterns[52677] = 25'b11001101_11000011_10010000_1;
      patterns[52678] = 25'b11001101_11000100_10010001_1;
      patterns[52679] = 25'b11001101_11000101_10010010_1;
      patterns[52680] = 25'b11001101_11000110_10010011_1;
      patterns[52681] = 25'b11001101_11000111_10010100_1;
      patterns[52682] = 25'b11001101_11001000_10010101_1;
      patterns[52683] = 25'b11001101_11001001_10010110_1;
      patterns[52684] = 25'b11001101_11001010_10010111_1;
      patterns[52685] = 25'b11001101_11001011_10011000_1;
      patterns[52686] = 25'b11001101_11001100_10011001_1;
      patterns[52687] = 25'b11001101_11001101_10011010_1;
      patterns[52688] = 25'b11001101_11001110_10011011_1;
      patterns[52689] = 25'b11001101_11001111_10011100_1;
      patterns[52690] = 25'b11001101_11010000_10011101_1;
      patterns[52691] = 25'b11001101_11010001_10011110_1;
      patterns[52692] = 25'b11001101_11010010_10011111_1;
      patterns[52693] = 25'b11001101_11010011_10100000_1;
      patterns[52694] = 25'b11001101_11010100_10100001_1;
      patterns[52695] = 25'b11001101_11010101_10100010_1;
      patterns[52696] = 25'b11001101_11010110_10100011_1;
      patterns[52697] = 25'b11001101_11010111_10100100_1;
      patterns[52698] = 25'b11001101_11011000_10100101_1;
      patterns[52699] = 25'b11001101_11011001_10100110_1;
      patterns[52700] = 25'b11001101_11011010_10100111_1;
      patterns[52701] = 25'b11001101_11011011_10101000_1;
      patterns[52702] = 25'b11001101_11011100_10101001_1;
      patterns[52703] = 25'b11001101_11011101_10101010_1;
      patterns[52704] = 25'b11001101_11011110_10101011_1;
      patterns[52705] = 25'b11001101_11011111_10101100_1;
      patterns[52706] = 25'b11001101_11100000_10101101_1;
      patterns[52707] = 25'b11001101_11100001_10101110_1;
      patterns[52708] = 25'b11001101_11100010_10101111_1;
      patterns[52709] = 25'b11001101_11100011_10110000_1;
      patterns[52710] = 25'b11001101_11100100_10110001_1;
      patterns[52711] = 25'b11001101_11100101_10110010_1;
      patterns[52712] = 25'b11001101_11100110_10110011_1;
      patterns[52713] = 25'b11001101_11100111_10110100_1;
      patterns[52714] = 25'b11001101_11101000_10110101_1;
      patterns[52715] = 25'b11001101_11101001_10110110_1;
      patterns[52716] = 25'b11001101_11101010_10110111_1;
      patterns[52717] = 25'b11001101_11101011_10111000_1;
      patterns[52718] = 25'b11001101_11101100_10111001_1;
      patterns[52719] = 25'b11001101_11101101_10111010_1;
      patterns[52720] = 25'b11001101_11101110_10111011_1;
      patterns[52721] = 25'b11001101_11101111_10111100_1;
      patterns[52722] = 25'b11001101_11110000_10111101_1;
      patterns[52723] = 25'b11001101_11110001_10111110_1;
      patterns[52724] = 25'b11001101_11110010_10111111_1;
      patterns[52725] = 25'b11001101_11110011_11000000_1;
      patterns[52726] = 25'b11001101_11110100_11000001_1;
      patterns[52727] = 25'b11001101_11110101_11000010_1;
      patterns[52728] = 25'b11001101_11110110_11000011_1;
      patterns[52729] = 25'b11001101_11110111_11000100_1;
      patterns[52730] = 25'b11001101_11111000_11000101_1;
      patterns[52731] = 25'b11001101_11111001_11000110_1;
      patterns[52732] = 25'b11001101_11111010_11000111_1;
      patterns[52733] = 25'b11001101_11111011_11001000_1;
      patterns[52734] = 25'b11001101_11111100_11001001_1;
      patterns[52735] = 25'b11001101_11111101_11001010_1;
      patterns[52736] = 25'b11001101_11111110_11001011_1;
      patterns[52737] = 25'b11001101_11111111_11001100_1;
      patterns[52738] = 25'b11001110_00000000_11001110_0;
      patterns[52739] = 25'b11001110_00000001_11001111_0;
      patterns[52740] = 25'b11001110_00000010_11010000_0;
      patterns[52741] = 25'b11001110_00000011_11010001_0;
      patterns[52742] = 25'b11001110_00000100_11010010_0;
      patterns[52743] = 25'b11001110_00000101_11010011_0;
      patterns[52744] = 25'b11001110_00000110_11010100_0;
      patterns[52745] = 25'b11001110_00000111_11010101_0;
      patterns[52746] = 25'b11001110_00001000_11010110_0;
      patterns[52747] = 25'b11001110_00001001_11010111_0;
      patterns[52748] = 25'b11001110_00001010_11011000_0;
      patterns[52749] = 25'b11001110_00001011_11011001_0;
      patterns[52750] = 25'b11001110_00001100_11011010_0;
      patterns[52751] = 25'b11001110_00001101_11011011_0;
      patterns[52752] = 25'b11001110_00001110_11011100_0;
      patterns[52753] = 25'b11001110_00001111_11011101_0;
      patterns[52754] = 25'b11001110_00010000_11011110_0;
      patterns[52755] = 25'b11001110_00010001_11011111_0;
      patterns[52756] = 25'b11001110_00010010_11100000_0;
      patterns[52757] = 25'b11001110_00010011_11100001_0;
      patterns[52758] = 25'b11001110_00010100_11100010_0;
      patterns[52759] = 25'b11001110_00010101_11100011_0;
      patterns[52760] = 25'b11001110_00010110_11100100_0;
      patterns[52761] = 25'b11001110_00010111_11100101_0;
      patterns[52762] = 25'b11001110_00011000_11100110_0;
      patterns[52763] = 25'b11001110_00011001_11100111_0;
      patterns[52764] = 25'b11001110_00011010_11101000_0;
      patterns[52765] = 25'b11001110_00011011_11101001_0;
      patterns[52766] = 25'b11001110_00011100_11101010_0;
      patterns[52767] = 25'b11001110_00011101_11101011_0;
      patterns[52768] = 25'b11001110_00011110_11101100_0;
      patterns[52769] = 25'b11001110_00011111_11101101_0;
      patterns[52770] = 25'b11001110_00100000_11101110_0;
      patterns[52771] = 25'b11001110_00100001_11101111_0;
      patterns[52772] = 25'b11001110_00100010_11110000_0;
      patterns[52773] = 25'b11001110_00100011_11110001_0;
      patterns[52774] = 25'b11001110_00100100_11110010_0;
      patterns[52775] = 25'b11001110_00100101_11110011_0;
      patterns[52776] = 25'b11001110_00100110_11110100_0;
      patterns[52777] = 25'b11001110_00100111_11110101_0;
      patterns[52778] = 25'b11001110_00101000_11110110_0;
      patterns[52779] = 25'b11001110_00101001_11110111_0;
      patterns[52780] = 25'b11001110_00101010_11111000_0;
      patterns[52781] = 25'b11001110_00101011_11111001_0;
      patterns[52782] = 25'b11001110_00101100_11111010_0;
      patterns[52783] = 25'b11001110_00101101_11111011_0;
      patterns[52784] = 25'b11001110_00101110_11111100_0;
      patterns[52785] = 25'b11001110_00101111_11111101_0;
      patterns[52786] = 25'b11001110_00110000_11111110_0;
      patterns[52787] = 25'b11001110_00110001_11111111_0;
      patterns[52788] = 25'b11001110_00110010_00000000_1;
      patterns[52789] = 25'b11001110_00110011_00000001_1;
      patterns[52790] = 25'b11001110_00110100_00000010_1;
      patterns[52791] = 25'b11001110_00110101_00000011_1;
      patterns[52792] = 25'b11001110_00110110_00000100_1;
      patterns[52793] = 25'b11001110_00110111_00000101_1;
      patterns[52794] = 25'b11001110_00111000_00000110_1;
      patterns[52795] = 25'b11001110_00111001_00000111_1;
      patterns[52796] = 25'b11001110_00111010_00001000_1;
      patterns[52797] = 25'b11001110_00111011_00001001_1;
      patterns[52798] = 25'b11001110_00111100_00001010_1;
      patterns[52799] = 25'b11001110_00111101_00001011_1;
      patterns[52800] = 25'b11001110_00111110_00001100_1;
      patterns[52801] = 25'b11001110_00111111_00001101_1;
      patterns[52802] = 25'b11001110_01000000_00001110_1;
      patterns[52803] = 25'b11001110_01000001_00001111_1;
      patterns[52804] = 25'b11001110_01000010_00010000_1;
      patterns[52805] = 25'b11001110_01000011_00010001_1;
      patterns[52806] = 25'b11001110_01000100_00010010_1;
      patterns[52807] = 25'b11001110_01000101_00010011_1;
      patterns[52808] = 25'b11001110_01000110_00010100_1;
      patterns[52809] = 25'b11001110_01000111_00010101_1;
      patterns[52810] = 25'b11001110_01001000_00010110_1;
      patterns[52811] = 25'b11001110_01001001_00010111_1;
      patterns[52812] = 25'b11001110_01001010_00011000_1;
      patterns[52813] = 25'b11001110_01001011_00011001_1;
      patterns[52814] = 25'b11001110_01001100_00011010_1;
      patterns[52815] = 25'b11001110_01001101_00011011_1;
      patterns[52816] = 25'b11001110_01001110_00011100_1;
      patterns[52817] = 25'b11001110_01001111_00011101_1;
      patterns[52818] = 25'b11001110_01010000_00011110_1;
      patterns[52819] = 25'b11001110_01010001_00011111_1;
      patterns[52820] = 25'b11001110_01010010_00100000_1;
      patterns[52821] = 25'b11001110_01010011_00100001_1;
      patterns[52822] = 25'b11001110_01010100_00100010_1;
      patterns[52823] = 25'b11001110_01010101_00100011_1;
      patterns[52824] = 25'b11001110_01010110_00100100_1;
      patterns[52825] = 25'b11001110_01010111_00100101_1;
      patterns[52826] = 25'b11001110_01011000_00100110_1;
      patterns[52827] = 25'b11001110_01011001_00100111_1;
      patterns[52828] = 25'b11001110_01011010_00101000_1;
      patterns[52829] = 25'b11001110_01011011_00101001_1;
      patterns[52830] = 25'b11001110_01011100_00101010_1;
      patterns[52831] = 25'b11001110_01011101_00101011_1;
      patterns[52832] = 25'b11001110_01011110_00101100_1;
      patterns[52833] = 25'b11001110_01011111_00101101_1;
      patterns[52834] = 25'b11001110_01100000_00101110_1;
      patterns[52835] = 25'b11001110_01100001_00101111_1;
      patterns[52836] = 25'b11001110_01100010_00110000_1;
      patterns[52837] = 25'b11001110_01100011_00110001_1;
      patterns[52838] = 25'b11001110_01100100_00110010_1;
      patterns[52839] = 25'b11001110_01100101_00110011_1;
      patterns[52840] = 25'b11001110_01100110_00110100_1;
      patterns[52841] = 25'b11001110_01100111_00110101_1;
      patterns[52842] = 25'b11001110_01101000_00110110_1;
      patterns[52843] = 25'b11001110_01101001_00110111_1;
      patterns[52844] = 25'b11001110_01101010_00111000_1;
      patterns[52845] = 25'b11001110_01101011_00111001_1;
      patterns[52846] = 25'b11001110_01101100_00111010_1;
      patterns[52847] = 25'b11001110_01101101_00111011_1;
      patterns[52848] = 25'b11001110_01101110_00111100_1;
      patterns[52849] = 25'b11001110_01101111_00111101_1;
      patterns[52850] = 25'b11001110_01110000_00111110_1;
      patterns[52851] = 25'b11001110_01110001_00111111_1;
      patterns[52852] = 25'b11001110_01110010_01000000_1;
      patterns[52853] = 25'b11001110_01110011_01000001_1;
      patterns[52854] = 25'b11001110_01110100_01000010_1;
      patterns[52855] = 25'b11001110_01110101_01000011_1;
      patterns[52856] = 25'b11001110_01110110_01000100_1;
      patterns[52857] = 25'b11001110_01110111_01000101_1;
      patterns[52858] = 25'b11001110_01111000_01000110_1;
      patterns[52859] = 25'b11001110_01111001_01000111_1;
      patterns[52860] = 25'b11001110_01111010_01001000_1;
      patterns[52861] = 25'b11001110_01111011_01001001_1;
      patterns[52862] = 25'b11001110_01111100_01001010_1;
      patterns[52863] = 25'b11001110_01111101_01001011_1;
      patterns[52864] = 25'b11001110_01111110_01001100_1;
      patterns[52865] = 25'b11001110_01111111_01001101_1;
      patterns[52866] = 25'b11001110_10000000_01001110_1;
      patterns[52867] = 25'b11001110_10000001_01001111_1;
      patterns[52868] = 25'b11001110_10000010_01010000_1;
      patterns[52869] = 25'b11001110_10000011_01010001_1;
      patterns[52870] = 25'b11001110_10000100_01010010_1;
      patterns[52871] = 25'b11001110_10000101_01010011_1;
      patterns[52872] = 25'b11001110_10000110_01010100_1;
      patterns[52873] = 25'b11001110_10000111_01010101_1;
      patterns[52874] = 25'b11001110_10001000_01010110_1;
      patterns[52875] = 25'b11001110_10001001_01010111_1;
      patterns[52876] = 25'b11001110_10001010_01011000_1;
      patterns[52877] = 25'b11001110_10001011_01011001_1;
      patterns[52878] = 25'b11001110_10001100_01011010_1;
      patterns[52879] = 25'b11001110_10001101_01011011_1;
      patterns[52880] = 25'b11001110_10001110_01011100_1;
      patterns[52881] = 25'b11001110_10001111_01011101_1;
      patterns[52882] = 25'b11001110_10010000_01011110_1;
      patterns[52883] = 25'b11001110_10010001_01011111_1;
      patterns[52884] = 25'b11001110_10010010_01100000_1;
      patterns[52885] = 25'b11001110_10010011_01100001_1;
      patterns[52886] = 25'b11001110_10010100_01100010_1;
      patterns[52887] = 25'b11001110_10010101_01100011_1;
      patterns[52888] = 25'b11001110_10010110_01100100_1;
      patterns[52889] = 25'b11001110_10010111_01100101_1;
      patterns[52890] = 25'b11001110_10011000_01100110_1;
      patterns[52891] = 25'b11001110_10011001_01100111_1;
      patterns[52892] = 25'b11001110_10011010_01101000_1;
      patterns[52893] = 25'b11001110_10011011_01101001_1;
      patterns[52894] = 25'b11001110_10011100_01101010_1;
      patterns[52895] = 25'b11001110_10011101_01101011_1;
      patterns[52896] = 25'b11001110_10011110_01101100_1;
      patterns[52897] = 25'b11001110_10011111_01101101_1;
      patterns[52898] = 25'b11001110_10100000_01101110_1;
      patterns[52899] = 25'b11001110_10100001_01101111_1;
      patterns[52900] = 25'b11001110_10100010_01110000_1;
      patterns[52901] = 25'b11001110_10100011_01110001_1;
      patterns[52902] = 25'b11001110_10100100_01110010_1;
      patterns[52903] = 25'b11001110_10100101_01110011_1;
      patterns[52904] = 25'b11001110_10100110_01110100_1;
      patterns[52905] = 25'b11001110_10100111_01110101_1;
      patterns[52906] = 25'b11001110_10101000_01110110_1;
      patterns[52907] = 25'b11001110_10101001_01110111_1;
      patterns[52908] = 25'b11001110_10101010_01111000_1;
      patterns[52909] = 25'b11001110_10101011_01111001_1;
      patterns[52910] = 25'b11001110_10101100_01111010_1;
      patterns[52911] = 25'b11001110_10101101_01111011_1;
      patterns[52912] = 25'b11001110_10101110_01111100_1;
      patterns[52913] = 25'b11001110_10101111_01111101_1;
      patterns[52914] = 25'b11001110_10110000_01111110_1;
      patterns[52915] = 25'b11001110_10110001_01111111_1;
      patterns[52916] = 25'b11001110_10110010_10000000_1;
      patterns[52917] = 25'b11001110_10110011_10000001_1;
      patterns[52918] = 25'b11001110_10110100_10000010_1;
      patterns[52919] = 25'b11001110_10110101_10000011_1;
      patterns[52920] = 25'b11001110_10110110_10000100_1;
      patterns[52921] = 25'b11001110_10110111_10000101_1;
      patterns[52922] = 25'b11001110_10111000_10000110_1;
      patterns[52923] = 25'b11001110_10111001_10000111_1;
      patterns[52924] = 25'b11001110_10111010_10001000_1;
      patterns[52925] = 25'b11001110_10111011_10001001_1;
      patterns[52926] = 25'b11001110_10111100_10001010_1;
      patterns[52927] = 25'b11001110_10111101_10001011_1;
      patterns[52928] = 25'b11001110_10111110_10001100_1;
      patterns[52929] = 25'b11001110_10111111_10001101_1;
      patterns[52930] = 25'b11001110_11000000_10001110_1;
      patterns[52931] = 25'b11001110_11000001_10001111_1;
      patterns[52932] = 25'b11001110_11000010_10010000_1;
      patterns[52933] = 25'b11001110_11000011_10010001_1;
      patterns[52934] = 25'b11001110_11000100_10010010_1;
      patterns[52935] = 25'b11001110_11000101_10010011_1;
      patterns[52936] = 25'b11001110_11000110_10010100_1;
      patterns[52937] = 25'b11001110_11000111_10010101_1;
      patterns[52938] = 25'b11001110_11001000_10010110_1;
      patterns[52939] = 25'b11001110_11001001_10010111_1;
      patterns[52940] = 25'b11001110_11001010_10011000_1;
      patterns[52941] = 25'b11001110_11001011_10011001_1;
      patterns[52942] = 25'b11001110_11001100_10011010_1;
      patterns[52943] = 25'b11001110_11001101_10011011_1;
      patterns[52944] = 25'b11001110_11001110_10011100_1;
      patterns[52945] = 25'b11001110_11001111_10011101_1;
      patterns[52946] = 25'b11001110_11010000_10011110_1;
      patterns[52947] = 25'b11001110_11010001_10011111_1;
      patterns[52948] = 25'b11001110_11010010_10100000_1;
      patterns[52949] = 25'b11001110_11010011_10100001_1;
      patterns[52950] = 25'b11001110_11010100_10100010_1;
      patterns[52951] = 25'b11001110_11010101_10100011_1;
      patterns[52952] = 25'b11001110_11010110_10100100_1;
      patterns[52953] = 25'b11001110_11010111_10100101_1;
      patterns[52954] = 25'b11001110_11011000_10100110_1;
      patterns[52955] = 25'b11001110_11011001_10100111_1;
      patterns[52956] = 25'b11001110_11011010_10101000_1;
      patterns[52957] = 25'b11001110_11011011_10101001_1;
      patterns[52958] = 25'b11001110_11011100_10101010_1;
      patterns[52959] = 25'b11001110_11011101_10101011_1;
      patterns[52960] = 25'b11001110_11011110_10101100_1;
      patterns[52961] = 25'b11001110_11011111_10101101_1;
      patterns[52962] = 25'b11001110_11100000_10101110_1;
      patterns[52963] = 25'b11001110_11100001_10101111_1;
      patterns[52964] = 25'b11001110_11100010_10110000_1;
      patterns[52965] = 25'b11001110_11100011_10110001_1;
      patterns[52966] = 25'b11001110_11100100_10110010_1;
      patterns[52967] = 25'b11001110_11100101_10110011_1;
      patterns[52968] = 25'b11001110_11100110_10110100_1;
      patterns[52969] = 25'b11001110_11100111_10110101_1;
      patterns[52970] = 25'b11001110_11101000_10110110_1;
      patterns[52971] = 25'b11001110_11101001_10110111_1;
      patterns[52972] = 25'b11001110_11101010_10111000_1;
      patterns[52973] = 25'b11001110_11101011_10111001_1;
      patterns[52974] = 25'b11001110_11101100_10111010_1;
      patterns[52975] = 25'b11001110_11101101_10111011_1;
      patterns[52976] = 25'b11001110_11101110_10111100_1;
      patterns[52977] = 25'b11001110_11101111_10111101_1;
      patterns[52978] = 25'b11001110_11110000_10111110_1;
      patterns[52979] = 25'b11001110_11110001_10111111_1;
      patterns[52980] = 25'b11001110_11110010_11000000_1;
      patterns[52981] = 25'b11001110_11110011_11000001_1;
      patterns[52982] = 25'b11001110_11110100_11000010_1;
      patterns[52983] = 25'b11001110_11110101_11000011_1;
      patterns[52984] = 25'b11001110_11110110_11000100_1;
      patterns[52985] = 25'b11001110_11110111_11000101_1;
      patterns[52986] = 25'b11001110_11111000_11000110_1;
      patterns[52987] = 25'b11001110_11111001_11000111_1;
      patterns[52988] = 25'b11001110_11111010_11001000_1;
      patterns[52989] = 25'b11001110_11111011_11001001_1;
      patterns[52990] = 25'b11001110_11111100_11001010_1;
      patterns[52991] = 25'b11001110_11111101_11001011_1;
      patterns[52992] = 25'b11001110_11111110_11001100_1;
      patterns[52993] = 25'b11001110_11111111_11001101_1;
      patterns[52994] = 25'b11001111_00000000_11001111_0;
      patterns[52995] = 25'b11001111_00000001_11010000_0;
      patterns[52996] = 25'b11001111_00000010_11010001_0;
      patterns[52997] = 25'b11001111_00000011_11010010_0;
      patterns[52998] = 25'b11001111_00000100_11010011_0;
      patterns[52999] = 25'b11001111_00000101_11010100_0;
      patterns[53000] = 25'b11001111_00000110_11010101_0;
      patterns[53001] = 25'b11001111_00000111_11010110_0;
      patterns[53002] = 25'b11001111_00001000_11010111_0;
      patterns[53003] = 25'b11001111_00001001_11011000_0;
      patterns[53004] = 25'b11001111_00001010_11011001_0;
      patterns[53005] = 25'b11001111_00001011_11011010_0;
      patterns[53006] = 25'b11001111_00001100_11011011_0;
      patterns[53007] = 25'b11001111_00001101_11011100_0;
      patterns[53008] = 25'b11001111_00001110_11011101_0;
      patterns[53009] = 25'b11001111_00001111_11011110_0;
      patterns[53010] = 25'b11001111_00010000_11011111_0;
      patterns[53011] = 25'b11001111_00010001_11100000_0;
      patterns[53012] = 25'b11001111_00010010_11100001_0;
      patterns[53013] = 25'b11001111_00010011_11100010_0;
      patterns[53014] = 25'b11001111_00010100_11100011_0;
      patterns[53015] = 25'b11001111_00010101_11100100_0;
      patterns[53016] = 25'b11001111_00010110_11100101_0;
      patterns[53017] = 25'b11001111_00010111_11100110_0;
      patterns[53018] = 25'b11001111_00011000_11100111_0;
      patterns[53019] = 25'b11001111_00011001_11101000_0;
      patterns[53020] = 25'b11001111_00011010_11101001_0;
      patterns[53021] = 25'b11001111_00011011_11101010_0;
      patterns[53022] = 25'b11001111_00011100_11101011_0;
      patterns[53023] = 25'b11001111_00011101_11101100_0;
      patterns[53024] = 25'b11001111_00011110_11101101_0;
      patterns[53025] = 25'b11001111_00011111_11101110_0;
      patterns[53026] = 25'b11001111_00100000_11101111_0;
      patterns[53027] = 25'b11001111_00100001_11110000_0;
      patterns[53028] = 25'b11001111_00100010_11110001_0;
      patterns[53029] = 25'b11001111_00100011_11110010_0;
      patterns[53030] = 25'b11001111_00100100_11110011_0;
      patterns[53031] = 25'b11001111_00100101_11110100_0;
      patterns[53032] = 25'b11001111_00100110_11110101_0;
      patterns[53033] = 25'b11001111_00100111_11110110_0;
      patterns[53034] = 25'b11001111_00101000_11110111_0;
      patterns[53035] = 25'b11001111_00101001_11111000_0;
      patterns[53036] = 25'b11001111_00101010_11111001_0;
      patterns[53037] = 25'b11001111_00101011_11111010_0;
      patterns[53038] = 25'b11001111_00101100_11111011_0;
      patterns[53039] = 25'b11001111_00101101_11111100_0;
      patterns[53040] = 25'b11001111_00101110_11111101_0;
      patterns[53041] = 25'b11001111_00101111_11111110_0;
      patterns[53042] = 25'b11001111_00110000_11111111_0;
      patterns[53043] = 25'b11001111_00110001_00000000_1;
      patterns[53044] = 25'b11001111_00110010_00000001_1;
      patterns[53045] = 25'b11001111_00110011_00000010_1;
      patterns[53046] = 25'b11001111_00110100_00000011_1;
      patterns[53047] = 25'b11001111_00110101_00000100_1;
      patterns[53048] = 25'b11001111_00110110_00000101_1;
      patterns[53049] = 25'b11001111_00110111_00000110_1;
      patterns[53050] = 25'b11001111_00111000_00000111_1;
      patterns[53051] = 25'b11001111_00111001_00001000_1;
      patterns[53052] = 25'b11001111_00111010_00001001_1;
      patterns[53053] = 25'b11001111_00111011_00001010_1;
      patterns[53054] = 25'b11001111_00111100_00001011_1;
      patterns[53055] = 25'b11001111_00111101_00001100_1;
      patterns[53056] = 25'b11001111_00111110_00001101_1;
      patterns[53057] = 25'b11001111_00111111_00001110_1;
      patterns[53058] = 25'b11001111_01000000_00001111_1;
      patterns[53059] = 25'b11001111_01000001_00010000_1;
      patterns[53060] = 25'b11001111_01000010_00010001_1;
      patterns[53061] = 25'b11001111_01000011_00010010_1;
      patterns[53062] = 25'b11001111_01000100_00010011_1;
      patterns[53063] = 25'b11001111_01000101_00010100_1;
      patterns[53064] = 25'b11001111_01000110_00010101_1;
      patterns[53065] = 25'b11001111_01000111_00010110_1;
      patterns[53066] = 25'b11001111_01001000_00010111_1;
      patterns[53067] = 25'b11001111_01001001_00011000_1;
      patterns[53068] = 25'b11001111_01001010_00011001_1;
      patterns[53069] = 25'b11001111_01001011_00011010_1;
      patterns[53070] = 25'b11001111_01001100_00011011_1;
      patterns[53071] = 25'b11001111_01001101_00011100_1;
      patterns[53072] = 25'b11001111_01001110_00011101_1;
      patterns[53073] = 25'b11001111_01001111_00011110_1;
      patterns[53074] = 25'b11001111_01010000_00011111_1;
      patterns[53075] = 25'b11001111_01010001_00100000_1;
      patterns[53076] = 25'b11001111_01010010_00100001_1;
      patterns[53077] = 25'b11001111_01010011_00100010_1;
      patterns[53078] = 25'b11001111_01010100_00100011_1;
      patterns[53079] = 25'b11001111_01010101_00100100_1;
      patterns[53080] = 25'b11001111_01010110_00100101_1;
      patterns[53081] = 25'b11001111_01010111_00100110_1;
      patterns[53082] = 25'b11001111_01011000_00100111_1;
      patterns[53083] = 25'b11001111_01011001_00101000_1;
      patterns[53084] = 25'b11001111_01011010_00101001_1;
      patterns[53085] = 25'b11001111_01011011_00101010_1;
      patterns[53086] = 25'b11001111_01011100_00101011_1;
      patterns[53087] = 25'b11001111_01011101_00101100_1;
      patterns[53088] = 25'b11001111_01011110_00101101_1;
      patterns[53089] = 25'b11001111_01011111_00101110_1;
      patterns[53090] = 25'b11001111_01100000_00101111_1;
      patterns[53091] = 25'b11001111_01100001_00110000_1;
      patterns[53092] = 25'b11001111_01100010_00110001_1;
      patterns[53093] = 25'b11001111_01100011_00110010_1;
      patterns[53094] = 25'b11001111_01100100_00110011_1;
      patterns[53095] = 25'b11001111_01100101_00110100_1;
      patterns[53096] = 25'b11001111_01100110_00110101_1;
      patterns[53097] = 25'b11001111_01100111_00110110_1;
      patterns[53098] = 25'b11001111_01101000_00110111_1;
      patterns[53099] = 25'b11001111_01101001_00111000_1;
      patterns[53100] = 25'b11001111_01101010_00111001_1;
      patterns[53101] = 25'b11001111_01101011_00111010_1;
      patterns[53102] = 25'b11001111_01101100_00111011_1;
      patterns[53103] = 25'b11001111_01101101_00111100_1;
      patterns[53104] = 25'b11001111_01101110_00111101_1;
      patterns[53105] = 25'b11001111_01101111_00111110_1;
      patterns[53106] = 25'b11001111_01110000_00111111_1;
      patterns[53107] = 25'b11001111_01110001_01000000_1;
      patterns[53108] = 25'b11001111_01110010_01000001_1;
      patterns[53109] = 25'b11001111_01110011_01000010_1;
      patterns[53110] = 25'b11001111_01110100_01000011_1;
      patterns[53111] = 25'b11001111_01110101_01000100_1;
      patterns[53112] = 25'b11001111_01110110_01000101_1;
      patterns[53113] = 25'b11001111_01110111_01000110_1;
      patterns[53114] = 25'b11001111_01111000_01000111_1;
      patterns[53115] = 25'b11001111_01111001_01001000_1;
      patterns[53116] = 25'b11001111_01111010_01001001_1;
      patterns[53117] = 25'b11001111_01111011_01001010_1;
      patterns[53118] = 25'b11001111_01111100_01001011_1;
      patterns[53119] = 25'b11001111_01111101_01001100_1;
      patterns[53120] = 25'b11001111_01111110_01001101_1;
      patterns[53121] = 25'b11001111_01111111_01001110_1;
      patterns[53122] = 25'b11001111_10000000_01001111_1;
      patterns[53123] = 25'b11001111_10000001_01010000_1;
      patterns[53124] = 25'b11001111_10000010_01010001_1;
      patterns[53125] = 25'b11001111_10000011_01010010_1;
      patterns[53126] = 25'b11001111_10000100_01010011_1;
      patterns[53127] = 25'b11001111_10000101_01010100_1;
      patterns[53128] = 25'b11001111_10000110_01010101_1;
      patterns[53129] = 25'b11001111_10000111_01010110_1;
      patterns[53130] = 25'b11001111_10001000_01010111_1;
      patterns[53131] = 25'b11001111_10001001_01011000_1;
      patterns[53132] = 25'b11001111_10001010_01011001_1;
      patterns[53133] = 25'b11001111_10001011_01011010_1;
      patterns[53134] = 25'b11001111_10001100_01011011_1;
      patterns[53135] = 25'b11001111_10001101_01011100_1;
      patterns[53136] = 25'b11001111_10001110_01011101_1;
      patterns[53137] = 25'b11001111_10001111_01011110_1;
      patterns[53138] = 25'b11001111_10010000_01011111_1;
      patterns[53139] = 25'b11001111_10010001_01100000_1;
      patterns[53140] = 25'b11001111_10010010_01100001_1;
      patterns[53141] = 25'b11001111_10010011_01100010_1;
      patterns[53142] = 25'b11001111_10010100_01100011_1;
      patterns[53143] = 25'b11001111_10010101_01100100_1;
      patterns[53144] = 25'b11001111_10010110_01100101_1;
      patterns[53145] = 25'b11001111_10010111_01100110_1;
      patterns[53146] = 25'b11001111_10011000_01100111_1;
      patterns[53147] = 25'b11001111_10011001_01101000_1;
      patterns[53148] = 25'b11001111_10011010_01101001_1;
      patterns[53149] = 25'b11001111_10011011_01101010_1;
      patterns[53150] = 25'b11001111_10011100_01101011_1;
      patterns[53151] = 25'b11001111_10011101_01101100_1;
      patterns[53152] = 25'b11001111_10011110_01101101_1;
      patterns[53153] = 25'b11001111_10011111_01101110_1;
      patterns[53154] = 25'b11001111_10100000_01101111_1;
      patterns[53155] = 25'b11001111_10100001_01110000_1;
      patterns[53156] = 25'b11001111_10100010_01110001_1;
      patterns[53157] = 25'b11001111_10100011_01110010_1;
      patterns[53158] = 25'b11001111_10100100_01110011_1;
      patterns[53159] = 25'b11001111_10100101_01110100_1;
      patterns[53160] = 25'b11001111_10100110_01110101_1;
      patterns[53161] = 25'b11001111_10100111_01110110_1;
      patterns[53162] = 25'b11001111_10101000_01110111_1;
      patterns[53163] = 25'b11001111_10101001_01111000_1;
      patterns[53164] = 25'b11001111_10101010_01111001_1;
      patterns[53165] = 25'b11001111_10101011_01111010_1;
      patterns[53166] = 25'b11001111_10101100_01111011_1;
      patterns[53167] = 25'b11001111_10101101_01111100_1;
      patterns[53168] = 25'b11001111_10101110_01111101_1;
      patterns[53169] = 25'b11001111_10101111_01111110_1;
      patterns[53170] = 25'b11001111_10110000_01111111_1;
      patterns[53171] = 25'b11001111_10110001_10000000_1;
      patterns[53172] = 25'b11001111_10110010_10000001_1;
      patterns[53173] = 25'b11001111_10110011_10000010_1;
      patterns[53174] = 25'b11001111_10110100_10000011_1;
      patterns[53175] = 25'b11001111_10110101_10000100_1;
      patterns[53176] = 25'b11001111_10110110_10000101_1;
      patterns[53177] = 25'b11001111_10110111_10000110_1;
      patterns[53178] = 25'b11001111_10111000_10000111_1;
      patterns[53179] = 25'b11001111_10111001_10001000_1;
      patterns[53180] = 25'b11001111_10111010_10001001_1;
      patterns[53181] = 25'b11001111_10111011_10001010_1;
      patterns[53182] = 25'b11001111_10111100_10001011_1;
      patterns[53183] = 25'b11001111_10111101_10001100_1;
      patterns[53184] = 25'b11001111_10111110_10001101_1;
      patterns[53185] = 25'b11001111_10111111_10001110_1;
      patterns[53186] = 25'b11001111_11000000_10001111_1;
      patterns[53187] = 25'b11001111_11000001_10010000_1;
      patterns[53188] = 25'b11001111_11000010_10010001_1;
      patterns[53189] = 25'b11001111_11000011_10010010_1;
      patterns[53190] = 25'b11001111_11000100_10010011_1;
      patterns[53191] = 25'b11001111_11000101_10010100_1;
      patterns[53192] = 25'b11001111_11000110_10010101_1;
      patterns[53193] = 25'b11001111_11000111_10010110_1;
      patterns[53194] = 25'b11001111_11001000_10010111_1;
      patterns[53195] = 25'b11001111_11001001_10011000_1;
      patterns[53196] = 25'b11001111_11001010_10011001_1;
      patterns[53197] = 25'b11001111_11001011_10011010_1;
      patterns[53198] = 25'b11001111_11001100_10011011_1;
      patterns[53199] = 25'b11001111_11001101_10011100_1;
      patterns[53200] = 25'b11001111_11001110_10011101_1;
      patterns[53201] = 25'b11001111_11001111_10011110_1;
      patterns[53202] = 25'b11001111_11010000_10011111_1;
      patterns[53203] = 25'b11001111_11010001_10100000_1;
      patterns[53204] = 25'b11001111_11010010_10100001_1;
      patterns[53205] = 25'b11001111_11010011_10100010_1;
      patterns[53206] = 25'b11001111_11010100_10100011_1;
      patterns[53207] = 25'b11001111_11010101_10100100_1;
      patterns[53208] = 25'b11001111_11010110_10100101_1;
      patterns[53209] = 25'b11001111_11010111_10100110_1;
      patterns[53210] = 25'b11001111_11011000_10100111_1;
      patterns[53211] = 25'b11001111_11011001_10101000_1;
      patterns[53212] = 25'b11001111_11011010_10101001_1;
      patterns[53213] = 25'b11001111_11011011_10101010_1;
      patterns[53214] = 25'b11001111_11011100_10101011_1;
      patterns[53215] = 25'b11001111_11011101_10101100_1;
      patterns[53216] = 25'b11001111_11011110_10101101_1;
      patterns[53217] = 25'b11001111_11011111_10101110_1;
      patterns[53218] = 25'b11001111_11100000_10101111_1;
      patterns[53219] = 25'b11001111_11100001_10110000_1;
      patterns[53220] = 25'b11001111_11100010_10110001_1;
      patterns[53221] = 25'b11001111_11100011_10110010_1;
      patterns[53222] = 25'b11001111_11100100_10110011_1;
      patterns[53223] = 25'b11001111_11100101_10110100_1;
      patterns[53224] = 25'b11001111_11100110_10110101_1;
      patterns[53225] = 25'b11001111_11100111_10110110_1;
      patterns[53226] = 25'b11001111_11101000_10110111_1;
      patterns[53227] = 25'b11001111_11101001_10111000_1;
      patterns[53228] = 25'b11001111_11101010_10111001_1;
      patterns[53229] = 25'b11001111_11101011_10111010_1;
      patterns[53230] = 25'b11001111_11101100_10111011_1;
      patterns[53231] = 25'b11001111_11101101_10111100_1;
      patterns[53232] = 25'b11001111_11101110_10111101_1;
      patterns[53233] = 25'b11001111_11101111_10111110_1;
      patterns[53234] = 25'b11001111_11110000_10111111_1;
      patterns[53235] = 25'b11001111_11110001_11000000_1;
      patterns[53236] = 25'b11001111_11110010_11000001_1;
      patterns[53237] = 25'b11001111_11110011_11000010_1;
      patterns[53238] = 25'b11001111_11110100_11000011_1;
      patterns[53239] = 25'b11001111_11110101_11000100_1;
      patterns[53240] = 25'b11001111_11110110_11000101_1;
      patterns[53241] = 25'b11001111_11110111_11000110_1;
      patterns[53242] = 25'b11001111_11111000_11000111_1;
      patterns[53243] = 25'b11001111_11111001_11001000_1;
      patterns[53244] = 25'b11001111_11111010_11001001_1;
      patterns[53245] = 25'b11001111_11111011_11001010_1;
      patterns[53246] = 25'b11001111_11111100_11001011_1;
      patterns[53247] = 25'b11001111_11111101_11001100_1;
      patterns[53248] = 25'b11001111_11111110_11001101_1;
      patterns[53249] = 25'b11001111_11111111_11001110_1;
      patterns[53250] = 25'b11010000_00000000_11010000_0;
      patterns[53251] = 25'b11010000_00000001_11010001_0;
      patterns[53252] = 25'b11010000_00000010_11010010_0;
      patterns[53253] = 25'b11010000_00000011_11010011_0;
      patterns[53254] = 25'b11010000_00000100_11010100_0;
      patterns[53255] = 25'b11010000_00000101_11010101_0;
      patterns[53256] = 25'b11010000_00000110_11010110_0;
      patterns[53257] = 25'b11010000_00000111_11010111_0;
      patterns[53258] = 25'b11010000_00001000_11011000_0;
      patterns[53259] = 25'b11010000_00001001_11011001_0;
      patterns[53260] = 25'b11010000_00001010_11011010_0;
      patterns[53261] = 25'b11010000_00001011_11011011_0;
      patterns[53262] = 25'b11010000_00001100_11011100_0;
      patterns[53263] = 25'b11010000_00001101_11011101_0;
      patterns[53264] = 25'b11010000_00001110_11011110_0;
      patterns[53265] = 25'b11010000_00001111_11011111_0;
      patterns[53266] = 25'b11010000_00010000_11100000_0;
      patterns[53267] = 25'b11010000_00010001_11100001_0;
      patterns[53268] = 25'b11010000_00010010_11100010_0;
      patterns[53269] = 25'b11010000_00010011_11100011_0;
      patterns[53270] = 25'b11010000_00010100_11100100_0;
      patterns[53271] = 25'b11010000_00010101_11100101_0;
      patterns[53272] = 25'b11010000_00010110_11100110_0;
      patterns[53273] = 25'b11010000_00010111_11100111_0;
      patterns[53274] = 25'b11010000_00011000_11101000_0;
      patterns[53275] = 25'b11010000_00011001_11101001_0;
      patterns[53276] = 25'b11010000_00011010_11101010_0;
      patterns[53277] = 25'b11010000_00011011_11101011_0;
      patterns[53278] = 25'b11010000_00011100_11101100_0;
      patterns[53279] = 25'b11010000_00011101_11101101_0;
      patterns[53280] = 25'b11010000_00011110_11101110_0;
      patterns[53281] = 25'b11010000_00011111_11101111_0;
      patterns[53282] = 25'b11010000_00100000_11110000_0;
      patterns[53283] = 25'b11010000_00100001_11110001_0;
      patterns[53284] = 25'b11010000_00100010_11110010_0;
      patterns[53285] = 25'b11010000_00100011_11110011_0;
      patterns[53286] = 25'b11010000_00100100_11110100_0;
      patterns[53287] = 25'b11010000_00100101_11110101_0;
      patterns[53288] = 25'b11010000_00100110_11110110_0;
      patterns[53289] = 25'b11010000_00100111_11110111_0;
      patterns[53290] = 25'b11010000_00101000_11111000_0;
      patterns[53291] = 25'b11010000_00101001_11111001_0;
      patterns[53292] = 25'b11010000_00101010_11111010_0;
      patterns[53293] = 25'b11010000_00101011_11111011_0;
      patterns[53294] = 25'b11010000_00101100_11111100_0;
      patterns[53295] = 25'b11010000_00101101_11111101_0;
      patterns[53296] = 25'b11010000_00101110_11111110_0;
      patterns[53297] = 25'b11010000_00101111_11111111_0;
      patterns[53298] = 25'b11010000_00110000_00000000_1;
      patterns[53299] = 25'b11010000_00110001_00000001_1;
      patterns[53300] = 25'b11010000_00110010_00000010_1;
      patterns[53301] = 25'b11010000_00110011_00000011_1;
      patterns[53302] = 25'b11010000_00110100_00000100_1;
      patterns[53303] = 25'b11010000_00110101_00000101_1;
      patterns[53304] = 25'b11010000_00110110_00000110_1;
      patterns[53305] = 25'b11010000_00110111_00000111_1;
      patterns[53306] = 25'b11010000_00111000_00001000_1;
      patterns[53307] = 25'b11010000_00111001_00001001_1;
      patterns[53308] = 25'b11010000_00111010_00001010_1;
      patterns[53309] = 25'b11010000_00111011_00001011_1;
      patterns[53310] = 25'b11010000_00111100_00001100_1;
      patterns[53311] = 25'b11010000_00111101_00001101_1;
      patterns[53312] = 25'b11010000_00111110_00001110_1;
      patterns[53313] = 25'b11010000_00111111_00001111_1;
      patterns[53314] = 25'b11010000_01000000_00010000_1;
      patterns[53315] = 25'b11010000_01000001_00010001_1;
      patterns[53316] = 25'b11010000_01000010_00010010_1;
      patterns[53317] = 25'b11010000_01000011_00010011_1;
      patterns[53318] = 25'b11010000_01000100_00010100_1;
      patterns[53319] = 25'b11010000_01000101_00010101_1;
      patterns[53320] = 25'b11010000_01000110_00010110_1;
      patterns[53321] = 25'b11010000_01000111_00010111_1;
      patterns[53322] = 25'b11010000_01001000_00011000_1;
      patterns[53323] = 25'b11010000_01001001_00011001_1;
      patterns[53324] = 25'b11010000_01001010_00011010_1;
      patterns[53325] = 25'b11010000_01001011_00011011_1;
      patterns[53326] = 25'b11010000_01001100_00011100_1;
      patterns[53327] = 25'b11010000_01001101_00011101_1;
      patterns[53328] = 25'b11010000_01001110_00011110_1;
      patterns[53329] = 25'b11010000_01001111_00011111_1;
      patterns[53330] = 25'b11010000_01010000_00100000_1;
      patterns[53331] = 25'b11010000_01010001_00100001_1;
      patterns[53332] = 25'b11010000_01010010_00100010_1;
      patterns[53333] = 25'b11010000_01010011_00100011_1;
      patterns[53334] = 25'b11010000_01010100_00100100_1;
      patterns[53335] = 25'b11010000_01010101_00100101_1;
      patterns[53336] = 25'b11010000_01010110_00100110_1;
      patterns[53337] = 25'b11010000_01010111_00100111_1;
      patterns[53338] = 25'b11010000_01011000_00101000_1;
      patterns[53339] = 25'b11010000_01011001_00101001_1;
      patterns[53340] = 25'b11010000_01011010_00101010_1;
      patterns[53341] = 25'b11010000_01011011_00101011_1;
      patterns[53342] = 25'b11010000_01011100_00101100_1;
      patterns[53343] = 25'b11010000_01011101_00101101_1;
      patterns[53344] = 25'b11010000_01011110_00101110_1;
      patterns[53345] = 25'b11010000_01011111_00101111_1;
      patterns[53346] = 25'b11010000_01100000_00110000_1;
      patterns[53347] = 25'b11010000_01100001_00110001_1;
      patterns[53348] = 25'b11010000_01100010_00110010_1;
      patterns[53349] = 25'b11010000_01100011_00110011_1;
      patterns[53350] = 25'b11010000_01100100_00110100_1;
      patterns[53351] = 25'b11010000_01100101_00110101_1;
      patterns[53352] = 25'b11010000_01100110_00110110_1;
      patterns[53353] = 25'b11010000_01100111_00110111_1;
      patterns[53354] = 25'b11010000_01101000_00111000_1;
      patterns[53355] = 25'b11010000_01101001_00111001_1;
      patterns[53356] = 25'b11010000_01101010_00111010_1;
      patterns[53357] = 25'b11010000_01101011_00111011_1;
      patterns[53358] = 25'b11010000_01101100_00111100_1;
      patterns[53359] = 25'b11010000_01101101_00111101_1;
      patterns[53360] = 25'b11010000_01101110_00111110_1;
      patterns[53361] = 25'b11010000_01101111_00111111_1;
      patterns[53362] = 25'b11010000_01110000_01000000_1;
      patterns[53363] = 25'b11010000_01110001_01000001_1;
      patterns[53364] = 25'b11010000_01110010_01000010_1;
      patterns[53365] = 25'b11010000_01110011_01000011_1;
      patterns[53366] = 25'b11010000_01110100_01000100_1;
      patterns[53367] = 25'b11010000_01110101_01000101_1;
      patterns[53368] = 25'b11010000_01110110_01000110_1;
      patterns[53369] = 25'b11010000_01110111_01000111_1;
      patterns[53370] = 25'b11010000_01111000_01001000_1;
      patterns[53371] = 25'b11010000_01111001_01001001_1;
      patterns[53372] = 25'b11010000_01111010_01001010_1;
      patterns[53373] = 25'b11010000_01111011_01001011_1;
      patterns[53374] = 25'b11010000_01111100_01001100_1;
      patterns[53375] = 25'b11010000_01111101_01001101_1;
      patterns[53376] = 25'b11010000_01111110_01001110_1;
      patterns[53377] = 25'b11010000_01111111_01001111_1;
      patterns[53378] = 25'b11010000_10000000_01010000_1;
      patterns[53379] = 25'b11010000_10000001_01010001_1;
      patterns[53380] = 25'b11010000_10000010_01010010_1;
      patterns[53381] = 25'b11010000_10000011_01010011_1;
      patterns[53382] = 25'b11010000_10000100_01010100_1;
      patterns[53383] = 25'b11010000_10000101_01010101_1;
      patterns[53384] = 25'b11010000_10000110_01010110_1;
      patterns[53385] = 25'b11010000_10000111_01010111_1;
      patterns[53386] = 25'b11010000_10001000_01011000_1;
      patterns[53387] = 25'b11010000_10001001_01011001_1;
      patterns[53388] = 25'b11010000_10001010_01011010_1;
      patterns[53389] = 25'b11010000_10001011_01011011_1;
      patterns[53390] = 25'b11010000_10001100_01011100_1;
      patterns[53391] = 25'b11010000_10001101_01011101_1;
      patterns[53392] = 25'b11010000_10001110_01011110_1;
      patterns[53393] = 25'b11010000_10001111_01011111_1;
      patterns[53394] = 25'b11010000_10010000_01100000_1;
      patterns[53395] = 25'b11010000_10010001_01100001_1;
      patterns[53396] = 25'b11010000_10010010_01100010_1;
      patterns[53397] = 25'b11010000_10010011_01100011_1;
      patterns[53398] = 25'b11010000_10010100_01100100_1;
      patterns[53399] = 25'b11010000_10010101_01100101_1;
      patterns[53400] = 25'b11010000_10010110_01100110_1;
      patterns[53401] = 25'b11010000_10010111_01100111_1;
      patterns[53402] = 25'b11010000_10011000_01101000_1;
      patterns[53403] = 25'b11010000_10011001_01101001_1;
      patterns[53404] = 25'b11010000_10011010_01101010_1;
      patterns[53405] = 25'b11010000_10011011_01101011_1;
      patterns[53406] = 25'b11010000_10011100_01101100_1;
      patterns[53407] = 25'b11010000_10011101_01101101_1;
      patterns[53408] = 25'b11010000_10011110_01101110_1;
      patterns[53409] = 25'b11010000_10011111_01101111_1;
      patterns[53410] = 25'b11010000_10100000_01110000_1;
      patterns[53411] = 25'b11010000_10100001_01110001_1;
      patterns[53412] = 25'b11010000_10100010_01110010_1;
      patterns[53413] = 25'b11010000_10100011_01110011_1;
      patterns[53414] = 25'b11010000_10100100_01110100_1;
      patterns[53415] = 25'b11010000_10100101_01110101_1;
      patterns[53416] = 25'b11010000_10100110_01110110_1;
      patterns[53417] = 25'b11010000_10100111_01110111_1;
      patterns[53418] = 25'b11010000_10101000_01111000_1;
      patterns[53419] = 25'b11010000_10101001_01111001_1;
      patterns[53420] = 25'b11010000_10101010_01111010_1;
      patterns[53421] = 25'b11010000_10101011_01111011_1;
      patterns[53422] = 25'b11010000_10101100_01111100_1;
      patterns[53423] = 25'b11010000_10101101_01111101_1;
      patterns[53424] = 25'b11010000_10101110_01111110_1;
      patterns[53425] = 25'b11010000_10101111_01111111_1;
      patterns[53426] = 25'b11010000_10110000_10000000_1;
      patterns[53427] = 25'b11010000_10110001_10000001_1;
      patterns[53428] = 25'b11010000_10110010_10000010_1;
      patterns[53429] = 25'b11010000_10110011_10000011_1;
      patterns[53430] = 25'b11010000_10110100_10000100_1;
      patterns[53431] = 25'b11010000_10110101_10000101_1;
      patterns[53432] = 25'b11010000_10110110_10000110_1;
      patterns[53433] = 25'b11010000_10110111_10000111_1;
      patterns[53434] = 25'b11010000_10111000_10001000_1;
      patterns[53435] = 25'b11010000_10111001_10001001_1;
      patterns[53436] = 25'b11010000_10111010_10001010_1;
      patterns[53437] = 25'b11010000_10111011_10001011_1;
      patterns[53438] = 25'b11010000_10111100_10001100_1;
      patterns[53439] = 25'b11010000_10111101_10001101_1;
      patterns[53440] = 25'b11010000_10111110_10001110_1;
      patterns[53441] = 25'b11010000_10111111_10001111_1;
      patterns[53442] = 25'b11010000_11000000_10010000_1;
      patterns[53443] = 25'b11010000_11000001_10010001_1;
      patterns[53444] = 25'b11010000_11000010_10010010_1;
      patterns[53445] = 25'b11010000_11000011_10010011_1;
      patterns[53446] = 25'b11010000_11000100_10010100_1;
      patterns[53447] = 25'b11010000_11000101_10010101_1;
      patterns[53448] = 25'b11010000_11000110_10010110_1;
      patterns[53449] = 25'b11010000_11000111_10010111_1;
      patterns[53450] = 25'b11010000_11001000_10011000_1;
      patterns[53451] = 25'b11010000_11001001_10011001_1;
      patterns[53452] = 25'b11010000_11001010_10011010_1;
      patterns[53453] = 25'b11010000_11001011_10011011_1;
      patterns[53454] = 25'b11010000_11001100_10011100_1;
      patterns[53455] = 25'b11010000_11001101_10011101_1;
      patterns[53456] = 25'b11010000_11001110_10011110_1;
      patterns[53457] = 25'b11010000_11001111_10011111_1;
      patterns[53458] = 25'b11010000_11010000_10100000_1;
      patterns[53459] = 25'b11010000_11010001_10100001_1;
      patterns[53460] = 25'b11010000_11010010_10100010_1;
      patterns[53461] = 25'b11010000_11010011_10100011_1;
      patterns[53462] = 25'b11010000_11010100_10100100_1;
      patterns[53463] = 25'b11010000_11010101_10100101_1;
      patterns[53464] = 25'b11010000_11010110_10100110_1;
      patterns[53465] = 25'b11010000_11010111_10100111_1;
      patterns[53466] = 25'b11010000_11011000_10101000_1;
      patterns[53467] = 25'b11010000_11011001_10101001_1;
      patterns[53468] = 25'b11010000_11011010_10101010_1;
      patterns[53469] = 25'b11010000_11011011_10101011_1;
      patterns[53470] = 25'b11010000_11011100_10101100_1;
      patterns[53471] = 25'b11010000_11011101_10101101_1;
      patterns[53472] = 25'b11010000_11011110_10101110_1;
      patterns[53473] = 25'b11010000_11011111_10101111_1;
      patterns[53474] = 25'b11010000_11100000_10110000_1;
      patterns[53475] = 25'b11010000_11100001_10110001_1;
      patterns[53476] = 25'b11010000_11100010_10110010_1;
      patterns[53477] = 25'b11010000_11100011_10110011_1;
      patterns[53478] = 25'b11010000_11100100_10110100_1;
      patterns[53479] = 25'b11010000_11100101_10110101_1;
      patterns[53480] = 25'b11010000_11100110_10110110_1;
      patterns[53481] = 25'b11010000_11100111_10110111_1;
      patterns[53482] = 25'b11010000_11101000_10111000_1;
      patterns[53483] = 25'b11010000_11101001_10111001_1;
      patterns[53484] = 25'b11010000_11101010_10111010_1;
      patterns[53485] = 25'b11010000_11101011_10111011_1;
      patterns[53486] = 25'b11010000_11101100_10111100_1;
      patterns[53487] = 25'b11010000_11101101_10111101_1;
      patterns[53488] = 25'b11010000_11101110_10111110_1;
      patterns[53489] = 25'b11010000_11101111_10111111_1;
      patterns[53490] = 25'b11010000_11110000_11000000_1;
      patterns[53491] = 25'b11010000_11110001_11000001_1;
      patterns[53492] = 25'b11010000_11110010_11000010_1;
      patterns[53493] = 25'b11010000_11110011_11000011_1;
      patterns[53494] = 25'b11010000_11110100_11000100_1;
      patterns[53495] = 25'b11010000_11110101_11000101_1;
      patterns[53496] = 25'b11010000_11110110_11000110_1;
      patterns[53497] = 25'b11010000_11110111_11000111_1;
      patterns[53498] = 25'b11010000_11111000_11001000_1;
      patterns[53499] = 25'b11010000_11111001_11001001_1;
      patterns[53500] = 25'b11010000_11111010_11001010_1;
      patterns[53501] = 25'b11010000_11111011_11001011_1;
      patterns[53502] = 25'b11010000_11111100_11001100_1;
      patterns[53503] = 25'b11010000_11111101_11001101_1;
      patterns[53504] = 25'b11010000_11111110_11001110_1;
      patterns[53505] = 25'b11010000_11111111_11001111_1;
      patterns[53506] = 25'b11010001_00000000_11010001_0;
      patterns[53507] = 25'b11010001_00000001_11010010_0;
      patterns[53508] = 25'b11010001_00000010_11010011_0;
      patterns[53509] = 25'b11010001_00000011_11010100_0;
      patterns[53510] = 25'b11010001_00000100_11010101_0;
      patterns[53511] = 25'b11010001_00000101_11010110_0;
      patterns[53512] = 25'b11010001_00000110_11010111_0;
      patterns[53513] = 25'b11010001_00000111_11011000_0;
      patterns[53514] = 25'b11010001_00001000_11011001_0;
      patterns[53515] = 25'b11010001_00001001_11011010_0;
      patterns[53516] = 25'b11010001_00001010_11011011_0;
      patterns[53517] = 25'b11010001_00001011_11011100_0;
      patterns[53518] = 25'b11010001_00001100_11011101_0;
      patterns[53519] = 25'b11010001_00001101_11011110_0;
      patterns[53520] = 25'b11010001_00001110_11011111_0;
      patterns[53521] = 25'b11010001_00001111_11100000_0;
      patterns[53522] = 25'b11010001_00010000_11100001_0;
      patterns[53523] = 25'b11010001_00010001_11100010_0;
      patterns[53524] = 25'b11010001_00010010_11100011_0;
      patterns[53525] = 25'b11010001_00010011_11100100_0;
      patterns[53526] = 25'b11010001_00010100_11100101_0;
      patterns[53527] = 25'b11010001_00010101_11100110_0;
      patterns[53528] = 25'b11010001_00010110_11100111_0;
      patterns[53529] = 25'b11010001_00010111_11101000_0;
      patterns[53530] = 25'b11010001_00011000_11101001_0;
      patterns[53531] = 25'b11010001_00011001_11101010_0;
      patterns[53532] = 25'b11010001_00011010_11101011_0;
      patterns[53533] = 25'b11010001_00011011_11101100_0;
      patterns[53534] = 25'b11010001_00011100_11101101_0;
      patterns[53535] = 25'b11010001_00011101_11101110_0;
      patterns[53536] = 25'b11010001_00011110_11101111_0;
      patterns[53537] = 25'b11010001_00011111_11110000_0;
      patterns[53538] = 25'b11010001_00100000_11110001_0;
      patterns[53539] = 25'b11010001_00100001_11110010_0;
      patterns[53540] = 25'b11010001_00100010_11110011_0;
      patterns[53541] = 25'b11010001_00100011_11110100_0;
      patterns[53542] = 25'b11010001_00100100_11110101_0;
      patterns[53543] = 25'b11010001_00100101_11110110_0;
      patterns[53544] = 25'b11010001_00100110_11110111_0;
      patterns[53545] = 25'b11010001_00100111_11111000_0;
      patterns[53546] = 25'b11010001_00101000_11111001_0;
      patterns[53547] = 25'b11010001_00101001_11111010_0;
      patterns[53548] = 25'b11010001_00101010_11111011_0;
      patterns[53549] = 25'b11010001_00101011_11111100_0;
      patterns[53550] = 25'b11010001_00101100_11111101_0;
      patterns[53551] = 25'b11010001_00101101_11111110_0;
      patterns[53552] = 25'b11010001_00101110_11111111_0;
      patterns[53553] = 25'b11010001_00101111_00000000_1;
      patterns[53554] = 25'b11010001_00110000_00000001_1;
      patterns[53555] = 25'b11010001_00110001_00000010_1;
      patterns[53556] = 25'b11010001_00110010_00000011_1;
      patterns[53557] = 25'b11010001_00110011_00000100_1;
      patterns[53558] = 25'b11010001_00110100_00000101_1;
      patterns[53559] = 25'b11010001_00110101_00000110_1;
      patterns[53560] = 25'b11010001_00110110_00000111_1;
      patterns[53561] = 25'b11010001_00110111_00001000_1;
      patterns[53562] = 25'b11010001_00111000_00001001_1;
      patterns[53563] = 25'b11010001_00111001_00001010_1;
      patterns[53564] = 25'b11010001_00111010_00001011_1;
      patterns[53565] = 25'b11010001_00111011_00001100_1;
      patterns[53566] = 25'b11010001_00111100_00001101_1;
      patterns[53567] = 25'b11010001_00111101_00001110_1;
      patterns[53568] = 25'b11010001_00111110_00001111_1;
      patterns[53569] = 25'b11010001_00111111_00010000_1;
      patterns[53570] = 25'b11010001_01000000_00010001_1;
      patterns[53571] = 25'b11010001_01000001_00010010_1;
      patterns[53572] = 25'b11010001_01000010_00010011_1;
      patterns[53573] = 25'b11010001_01000011_00010100_1;
      patterns[53574] = 25'b11010001_01000100_00010101_1;
      patterns[53575] = 25'b11010001_01000101_00010110_1;
      patterns[53576] = 25'b11010001_01000110_00010111_1;
      patterns[53577] = 25'b11010001_01000111_00011000_1;
      patterns[53578] = 25'b11010001_01001000_00011001_1;
      patterns[53579] = 25'b11010001_01001001_00011010_1;
      patterns[53580] = 25'b11010001_01001010_00011011_1;
      patterns[53581] = 25'b11010001_01001011_00011100_1;
      patterns[53582] = 25'b11010001_01001100_00011101_1;
      patterns[53583] = 25'b11010001_01001101_00011110_1;
      patterns[53584] = 25'b11010001_01001110_00011111_1;
      patterns[53585] = 25'b11010001_01001111_00100000_1;
      patterns[53586] = 25'b11010001_01010000_00100001_1;
      patterns[53587] = 25'b11010001_01010001_00100010_1;
      patterns[53588] = 25'b11010001_01010010_00100011_1;
      patterns[53589] = 25'b11010001_01010011_00100100_1;
      patterns[53590] = 25'b11010001_01010100_00100101_1;
      patterns[53591] = 25'b11010001_01010101_00100110_1;
      patterns[53592] = 25'b11010001_01010110_00100111_1;
      patterns[53593] = 25'b11010001_01010111_00101000_1;
      patterns[53594] = 25'b11010001_01011000_00101001_1;
      patterns[53595] = 25'b11010001_01011001_00101010_1;
      patterns[53596] = 25'b11010001_01011010_00101011_1;
      patterns[53597] = 25'b11010001_01011011_00101100_1;
      patterns[53598] = 25'b11010001_01011100_00101101_1;
      patterns[53599] = 25'b11010001_01011101_00101110_1;
      patterns[53600] = 25'b11010001_01011110_00101111_1;
      patterns[53601] = 25'b11010001_01011111_00110000_1;
      patterns[53602] = 25'b11010001_01100000_00110001_1;
      patterns[53603] = 25'b11010001_01100001_00110010_1;
      patterns[53604] = 25'b11010001_01100010_00110011_1;
      patterns[53605] = 25'b11010001_01100011_00110100_1;
      patterns[53606] = 25'b11010001_01100100_00110101_1;
      patterns[53607] = 25'b11010001_01100101_00110110_1;
      patterns[53608] = 25'b11010001_01100110_00110111_1;
      patterns[53609] = 25'b11010001_01100111_00111000_1;
      patterns[53610] = 25'b11010001_01101000_00111001_1;
      patterns[53611] = 25'b11010001_01101001_00111010_1;
      patterns[53612] = 25'b11010001_01101010_00111011_1;
      patterns[53613] = 25'b11010001_01101011_00111100_1;
      patterns[53614] = 25'b11010001_01101100_00111101_1;
      patterns[53615] = 25'b11010001_01101101_00111110_1;
      patterns[53616] = 25'b11010001_01101110_00111111_1;
      patterns[53617] = 25'b11010001_01101111_01000000_1;
      patterns[53618] = 25'b11010001_01110000_01000001_1;
      patterns[53619] = 25'b11010001_01110001_01000010_1;
      patterns[53620] = 25'b11010001_01110010_01000011_1;
      patterns[53621] = 25'b11010001_01110011_01000100_1;
      patterns[53622] = 25'b11010001_01110100_01000101_1;
      patterns[53623] = 25'b11010001_01110101_01000110_1;
      patterns[53624] = 25'b11010001_01110110_01000111_1;
      patterns[53625] = 25'b11010001_01110111_01001000_1;
      patterns[53626] = 25'b11010001_01111000_01001001_1;
      patterns[53627] = 25'b11010001_01111001_01001010_1;
      patterns[53628] = 25'b11010001_01111010_01001011_1;
      patterns[53629] = 25'b11010001_01111011_01001100_1;
      patterns[53630] = 25'b11010001_01111100_01001101_1;
      patterns[53631] = 25'b11010001_01111101_01001110_1;
      patterns[53632] = 25'b11010001_01111110_01001111_1;
      patterns[53633] = 25'b11010001_01111111_01010000_1;
      patterns[53634] = 25'b11010001_10000000_01010001_1;
      patterns[53635] = 25'b11010001_10000001_01010010_1;
      patterns[53636] = 25'b11010001_10000010_01010011_1;
      patterns[53637] = 25'b11010001_10000011_01010100_1;
      patterns[53638] = 25'b11010001_10000100_01010101_1;
      patterns[53639] = 25'b11010001_10000101_01010110_1;
      patterns[53640] = 25'b11010001_10000110_01010111_1;
      patterns[53641] = 25'b11010001_10000111_01011000_1;
      patterns[53642] = 25'b11010001_10001000_01011001_1;
      patterns[53643] = 25'b11010001_10001001_01011010_1;
      patterns[53644] = 25'b11010001_10001010_01011011_1;
      patterns[53645] = 25'b11010001_10001011_01011100_1;
      patterns[53646] = 25'b11010001_10001100_01011101_1;
      patterns[53647] = 25'b11010001_10001101_01011110_1;
      patterns[53648] = 25'b11010001_10001110_01011111_1;
      patterns[53649] = 25'b11010001_10001111_01100000_1;
      patterns[53650] = 25'b11010001_10010000_01100001_1;
      patterns[53651] = 25'b11010001_10010001_01100010_1;
      patterns[53652] = 25'b11010001_10010010_01100011_1;
      patterns[53653] = 25'b11010001_10010011_01100100_1;
      patterns[53654] = 25'b11010001_10010100_01100101_1;
      patterns[53655] = 25'b11010001_10010101_01100110_1;
      patterns[53656] = 25'b11010001_10010110_01100111_1;
      patterns[53657] = 25'b11010001_10010111_01101000_1;
      patterns[53658] = 25'b11010001_10011000_01101001_1;
      patterns[53659] = 25'b11010001_10011001_01101010_1;
      patterns[53660] = 25'b11010001_10011010_01101011_1;
      patterns[53661] = 25'b11010001_10011011_01101100_1;
      patterns[53662] = 25'b11010001_10011100_01101101_1;
      patterns[53663] = 25'b11010001_10011101_01101110_1;
      patterns[53664] = 25'b11010001_10011110_01101111_1;
      patterns[53665] = 25'b11010001_10011111_01110000_1;
      patterns[53666] = 25'b11010001_10100000_01110001_1;
      patterns[53667] = 25'b11010001_10100001_01110010_1;
      patterns[53668] = 25'b11010001_10100010_01110011_1;
      patterns[53669] = 25'b11010001_10100011_01110100_1;
      patterns[53670] = 25'b11010001_10100100_01110101_1;
      patterns[53671] = 25'b11010001_10100101_01110110_1;
      patterns[53672] = 25'b11010001_10100110_01110111_1;
      patterns[53673] = 25'b11010001_10100111_01111000_1;
      patterns[53674] = 25'b11010001_10101000_01111001_1;
      patterns[53675] = 25'b11010001_10101001_01111010_1;
      patterns[53676] = 25'b11010001_10101010_01111011_1;
      patterns[53677] = 25'b11010001_10101011_01111100_1;
      patterns[53678] = 25'b11010001_10101100_01111101_1;
      patterns[53679] = 25'b11010001_10101101_01111110_1;
      patterns[53680] = 25'b11010001_10101110_01111111_1;
      patterns[53681] = 25'b11010001_10101111_10000000_1;
      patterns[53682] = 25'b11010001_10110000_10000001_1;
      patterns[53683] = 25'b11010001_10110001_10000010_1;
      patterns[53684] = 25'b11010001_10110010_10000011_1;
      patterns[53685] = 25'b11010001_10110011_10000100_1;
      patterns[53686] = 25'b11010001_10110100_10000101_1;
      patterns[53687] = 25'b11010001_10110101_10000110_1;
      patterns[53688] = 25'b11010001_10110110_10000111_1;
      patterns[53689] = 25'b11010001_10110111_10001000_1;
      patterns[53690] = 25'b11010001_10111000_10001001_1;
      patterns[53691] = 25'b11010001_10111001_10001010_1;
      patterns[53692] = 25'b11010001_10111010_10001011_1;
      patterns[53693] = 25'b11010001_10111011_10001100_1;
      patterns[53694] = 25'b11010001_10111100_10001101_1;
      patterns[53695] = 25'b11010001_10111101_10001110_1;
      patterns[53696] = 25'b11010001_10111110_10001111_1;
      patterns[53697] = 25'b11010001_10111111_10010000_1;
      patterns[53698] = 25'b11010001_11000000_10010001_1;
      patterns[53699] = 25'b11010001_11000001_10010010_1;
      patterns[53700] = 25'b11010001_11000010_10010011_1;
      patterns[53701] = 25'b11010001_11000011_10010100_1;
      patterns[53702] = 25'b11010001_11000100_10010101_1;
      patterns[53703] = 25'b11010001_11000101_10010110_1;
      patterns[53704] = 25'b11010001_11000110_10010111_1;
      patterns[53705] = 25'b11010001_11000111_10011000_1;
      patterns[53706] = 25'b11010001_11001000_10011001_1;
      patterns[53707] = 25'b11010001_11001001_10011010_1;
      patterns[53708] = 25'b11010001_11001010_10011011_1;
      patterns[53709] = 25'b11010001_11001011_10011100_1;
      patterns[53710] = 25'b11010001_11001100_10011101_1;
      patterns[53711] = 25'b11010001_11001101_10011110_1;
      patterns[53712] = 25'b11010001_11001110_10011111_1;
      patterns[53713] = 25'b11010001_11001111_10100000_1;
      patterns[53714] = 25'b11010001_11010000_10100001_1;
      patterns[53715] = 25'b11010001_11010001_10100010_1;
      patterns[53716] = 25'b11010001_11010010_10100011_1;
      patterns[53717] = 25'b11010001_11010011_10100100_1;
      patterns[53718] = 25'b11010001_11010100_10100101_1;
      patterns[53719] = 25'b11010001_11010101_10100110_1;
      patterns[53720] = 25'b11010001_11010110_10100111_1;
      patterns[53721] = 25'b11010001_11010111_10101000_1;
      patterns[53722] = 25'b11010001_11011000_10101001_1;
      patterns[53723] = 25'b11010001_11011001_10101010_1;
      patterns[53724] = 25'b11010001_11011010_10101011_1;
      patterns[53725] = 25'b11010001_11011011_10101100_1;
      patterns[53726] = 25'b11010001_11011100_10101101_1;
      patterns[53727] = 25'b11010001_11011101_10101110_1;
      patterns[53728] = 25'b11010001_11011110_10101111_1;
      patterns[53729] = 25'b11010001_11011111_10110000_1;
      patterns[53730] = 25'b11010001_11100000_10110001_1;
      patterns[53731] = 25'b11010001_11100001_10110010_1;
      patterns[53732] = 25'b11010001_11100010_10110011_1;
      patterns[53733] = 25'b11010001_11100011_10110100_1;
      patterns[53734] = 25'b11010001_11100100_10110101_1;
      patterns[53735] = 25'b11010001_11100101_10110110_1;
      patterns[53736] = 25'b11010001_11100110_10110111_1;
      patterns[53737] = 25'b11010001_11100111_10111000_1;
      patterns[53738] = 25'b11010001_11101000_10111001_1;
      patterns[53739] = 25'b11010001_11101001_10111010_1;
      patterns[53740] = 25'b11010001_11101010_10111011_1;
      patterns[53741] = 25'b11010001_11101011_10111100_1;
      patterns[53742] = 25'b11010001_11101100_10111101_1;
      patterns[53743] = 25'b11010001_11101101_10111110_1;
      patterns[53744] = 25'b11010001_11101110_10111111_1;
      patterns[53745] = 25'b11010001_11101111_11000000_1;
      patterns[53746] = 25'b11010001_11110000_11000001_1;
      patterns[53747] = 25'b11010001_11110001_11000010_1;
      patterns[53748] = 25'b11010001_11110010_11000011_1;
      patterns[53749] = 25'b11010001_11110011_11000100_1;
      patterns[53750] = 25'b11010001_11110100_11000101_1;
      patterns[53751] = 25'b11010001_11110101_11000110_1;
      patterns[53752] = 25'b11010001_11110110_11000111_1;
      patterns[53753] = 25'b11010001_11110111_11001000_1;
      patterns[53754] = 25'b11010001_11111000_11001001_1;
      patterns[53755] = 25'b11010001_11111001_11001010_1;
      patterns[53756] = 25'b11010001_11111010_11001011_1;
      patterns[53757] = 25'b11010001_11111011_11001100_1;
      patterns[53758] = 25'b11010001_11111100_11001101_1;
      patterns[53759] = 25'b11010001_11111101_11001110_1;
      patterns[53760] = 25'b11010001_11111110_11001111_1;
      patterns[53761] = 25'b11010001_11111111_11010000_1;
      patterns[53762] = 25'b11010010_00000000_11010010_0;
      patterns[53763] = 25'b11010010_00000001_11010011_0;
      patterns[53764] = 25'b11010010_00000010_11010100_0;
      patterns[53765] = 25'b11010010_00000011_11010101_0;
      patterns[53766] = 25'b11010010_00000100_11010110_0;
      patterns[53767] = 25'b11010010_00000101_11010111_0;
      patterns[53768] = 25'b11010010_00000110_11011000_0;
      patterns[53769] = 25'b11010010_00000111_11011001_0;
      patterns[53770] = 25'b11010010_00001000_11011010_0;
      patterns[53771] = 25'b11010010_00001001_11011011_0;
      patterns[53772] = 25'b11010010_00001010_11011100_0;
      patterns[53773] = 25'b11010010_00001011_11011101_0;
      patterns[53774] = 25'b11010010_00001100_11011110_0;
      patterns[53775] = 25'b11010010_00001101_11011111_0;
      patterns[53776] = 25'b11010010_00001110_11100000_0;
      patterns[53777] = 25'b11010010_00001111_11100001_0;
      patterns[53778] = 25'b11010010_00010000_11100010_0;
      patterns[53779] = 25'b11010010_00010001_11100011_0;
      patterns[53780] = 25'b11010010_00010010_11100100_0;
      patterns[53781] = 25'b11010010_00010011_11100101_0;
      patterns[53782] = 25'b11010010_00010100_11100110_0;
      patterns[53783] = 25'b11010010_00010101_11100111_0;
      patterns[53784] = 25'b11010010_00010110_11101000_0;
      patterns[53785] = 25'b11010010_00010111_11101001_0;
      patterns[53786] = 25'b11010010_00011000_11101010_0;
      patterns[53787] = 25'b11010010_00011001_11101011_0;
      patterns[53788] = 25'b11010010_00011010_11101100_0;
      patterns[53789] = 25'b11010010_00011011_11101101_0;
      patterns[53790] = 25'b11010010_00011100_11101110_0;
      patterns[53791] = 25'b11010010_00011101_11101111_0;
      patterns[53792] = 25'b11010010_00011110_11110000_0;
      patterns[53793] = 25'b11010010_00011111_11110001_0;
      patterns[53794] = 25'b11010010_00100000_11110010_0;
      patterns[53795] = 25'b11010010_00100001_11110011_0;
      patterns[53796] = 25'b11010010_00100010_11110100_0;
      patterns[53797] = 25'b11010010_00100011_11110101_0;
      patterns[53798] = 25'b11010010_00100100_11110110_0;
      patterns[53799] = 25'b11010010_00100101_11110111_0;
      patterns[53800] = 25'b11010010_00100110_11111000_0;
      patterns[53801] = 25'b11010010_00100111_11111001_0;
      patterns[53802] = 25'b11010010_00101000_11111010_0;
      patterns[53803] = 25'b11010010_00101001_11111011_0;
      patterns[53804] = 25'b11010010_00101010_11111100_0;
      patterns[53805] = 25'b11010010_00101011_11111101_0;
      patterns[53806] = 25'b11010010_00101100_11111110_0;
      patterns[53807] = 25'b11010010_00101101_11111111_0;
      patterns[53808] = 25'b11010010_00101110_00000000_1;
      patterns[53809] = 25'b11010010_00101111_00000001_1;
      patterns[53810] = 25'b11010010_00110000_00000010_1;
      patterns[53811] = 25'b11010010_00110001_00000011_1;
      patterns[53812] = 25'b11010010_00110010_00000100_1;
      patterns[53813] = 25'b11010010_00110011_00000101_1;
      patterns[53814] = 25'b11010010_00110100_00000110_1;
      patterns[53815] = 25'b11010010_00110101_00000111_1;
      patterns[53816] = 25'b11010010_00110110_00001000_1;
      patterns[53817] = 25'b11010010_00110111_00001001_1;
      patterns[53818] = 25'b11010010_00111000_00001010_1;
      patterns[53819] = 25'b11010010_00111001_00001011_1;
      patterns[53820] = 25'b11010010_00111010_00001100_1;
      patterns[53821] = 25'b11010010_00111011_00001101_1;
      patterns[53822] = 25'b11010010_00111100_00001110_1;
      patterns[53823] = 25'b11010010_00111101_00001111_1;
      patterns[53824] = 25'b11010010_00111110_00010000_1;
      patterns[53825] = 25'b11010010_00111111_00010001_1;
      patterns[53826] = 25'b11010010_01000000_00010010_1;
      patterns[53827] = 25'b11010010_01000001_00010011_1;
      patterns[53828] = 25'b11010010_01000010_00010100_1;
      patterns[53829] = 25'b11010010_01000011_00010101_1;
      patterns[53830] = 25'b11010010_01000100_00010110_1;
      patterns[53831] = 25'b11010010_01000101_00010111_1;
      patterns[53832] = 25'b11010010_01000110_00011000_1;
      patterns[53833] = 25'b11010010_01000111_00011001_1;
      patterns[53834] = 25'b11010010_01001000_00011010_1;
      patterns[53835] = 25'b11010010_01001001_00011011_1;
      patterns[53836] = 25'b11010010_01001010_00011100_1;
      patterns[53837] = 25'b11010010_01001011_00011101_1;
      patterns[53838] = 25'b11010010_01001100_00011110_1;
      patterns[53839] = 25'b11010010_01001101_00011111_1;
      patterns[53840] = 25'b11010010_01001110_00100000_1;
      patterns[53841] = 25'b11010010_01001111_00100001_1;
      patterns[53842] = 25'b11010010_01010000_00100010_1;
      patterns[53843] = 25'b11010010_01010001_00100011_1;
      patterns[53844] = 25'b11010010_01010010_00100100_1;
      patterns[53845] = 25'b11010010_01010011_00100101_1;
      patterns[53846] = 25'b11010010_01010100_00100110_1;
      patterns[53847] = 25'b11010010_01010101_00100111_1;
      patterns[53848] = 25'b11010010_01010110_00101000_1;
      patterns[53849] = 25'b11010010_01010111_00101001_1;
      patterns[53850] = 25'b11010010_01011000_00101010_1;
      patterns[53851] = 25'b11010010_01011001_00101011_1;
      patterns[53852] = 25'b11010010_01011010_00101100_1;
      patterns[53853] = 25'b11010010_01011011_00101101_1;
      patterns[53854] = 25'b11010010_01011100_00101110_1;
      patterns[53855] = 25'b11010010_01011101_00101111_1;
      patterns[53856] = 25'b11010010_01011110_00110000_1;
      patterns[53857] = 25'b11010010_01011111_00110001_1;
      patterns[53858] = 25'b11010010_01100000_00110010_1;
      patterns[53859] = 25'b11010010_01100001_00110011_1;
      patterns[53860] = 25'b11010010_01100010_00110100_1;
      patterns[53861] = 25'b11010010_01100011_00110101_1;
      patterns[53862] = 25'b11010010_01100100_00110110_1;
      patterns[53863] = 25'b11010010_01100101_00110111_1;
      patterns[53864] = 25'b11010010_01100110_00111000_1;
      patterns[53865] = 25'b11010010_01100111_00111001_1;
      patterns[53866] = 25'b11010010_01101000_00111010_1;
      patterns[53867] = 25'b11010010_01101001_00111011_1;
      patterns[53868] = 25'b11010010_01101010_00111100_1;
      patterns[53869] = 25'b11010010_01101011_00111101_1;
      patterns[53870] = 25'b11010010_01101100_00111110_1;
      patterns[53871] = 25'b11010010_01101101_00111111_1;
      patterns[53872] = 25'b11010010_01101110_01000000_1;
      patterns[53873] = 25'b11010010_01101111_01000001_1;
      patterns[53874] = 25'b11010010_01110000_01000010_1;
      patterns[53875] = 25'b11010010_01110001_01000011_1;
      patterns[53876] = 25'b11010010_01110010_01000100_1;
      patterns[53877] = 25'b11010010_01110011_01000101_1;
      patterns[53878] = 25'b11010010_01110100_01000110_1;
      patterns[53879] = 25'b11010010_01110101_01000111_1;
      patterns[53880] = 25'b11010010_01110110_01001000_1;
      patterns[53881] = 25'b11010010_01110111_01001001_1;
      patterns[53882] = 25'b11010010_01111000_01001010_1;
      patterns[53883] = 25'b11010010_01111001_01001011_1;
      patterns[53884] = 25'b11010010_01111010_01001100_1;
      patterns[53885] = 25'b11010010_01111011_01001101_1;
      patterns[53886] = 25'b11010010_01111100_01001110_1;
      patterns[53887] = 25'b11010010_01111101_01001111_1;
      patterns[53888] = 25'b11010010_01111110_01010000_1;
      patterns[53889] = 25'b11010010_01111111_01010001_1;
      patterns[53890] = 25'b11010010_10000000_01010010_1;
      patterns[53891] = 25'b11010010_10000001_01010011_1;
      patterns[53892] = 25'b11010010_10000010_01010100_1;
      patterns[53893] = 25'b11010010_10000011_01010101_1;
      patterns[53894] = 25'b11010010_10000100_01010110_1;
      patterns[53895] = 25'b11010010_10000101_01010111_1;
      patterns[53896] = 25'b11010010_10000110_01011000_1;
      patterns[53897] = 25'b11010010_10000111_01011001_1;
      patterns[53898] = 25'b11010010_10001000_01011010_1;
      patterns[53899] = 25'b11010010_10001001_01011011_1;
      patterns[53900] = 25'b11010010_10001010_01011100_1;
      patterns[53901] = 25'b11010010_10001011_01011101_1;
      patterns[53902] = 25'b11010010_10001100_01011110_1;
      patterns[53903] = 25'b11010010_10001101_01011111_1;
      patterns[53904] = 25'b11010010_10001110_01100000_1;
      patterns[53905] = 25'b11010010_10001111_01100001_1;
      patterns[53906] = 25'b11010010_10010000_01100010_1;
      patterns[53907] = 25'b11010010_10010001_01100011_1;
      patterns[53908] = 25'b11010010_10010010_01100100_1;
      patterns[53909] = 25'b11010010_10010011_01100101_1;
      patterns[53910] = 25'b11010010_10010100_01100110_1;
      patterns[53911] = 25'b11010010_10010101_01100111_1;
      patterns[53912] = 25'b11010010_10010110_01101000_1;
      patterns[53913] = 25'b11010010_10010111_01101001_1;
      patterns[53914] = 25'b11010010_10011000_01101010_1;
      patterns[53915] = 25'b11010010_10011001_01101011_1;
      patterns[53916] = 25'b11010010_10011010_01101100_1;
      patterns[53917] = 25'b11010010_10011011_01101101_1;
      patterns[53918] = 25'b11010010_10011100_01101110_1;
      patterns[53919] = 25'b11010010_10011101_01101111_1;
      patterns[53920] = 25'b11010010_10011110_01110000_1;
      patterns[53921] = 25'b11010010_10011111_01110001_1;
      patterns[53922] = 25'b11010010_10100000_01110010_1;
      patterns[53923] = 25'b11010010_10100001_01110011_1;
      patterns[53924] = 25'b11010010_10100010_01110100_1;
      patterns[53925] = 25'b11010010_10100011_01110101_1;
      patterns[53926] = 25'b11010010_10100100_01110110_1;
      patterns[53927] = 25'b11010010_10100101_01110111_1;
      patterns[53928] = 25'b11010010_10100110_01111000_1;
      patterns[53929] = 25'b11010010_10100111_01111001_1;
      patterns[53930] = 25'b11010010_10101000_01111010_1;
      patterns[53931] = 25'b11010010_10101001_01111011_1;
      patterns[53932] = 25'b11010010_10101010_01111100_1;
      patterns[53933] = 25'b11010010_10101011_01111101_1;
      patterns[53934] = 25'b11010010_10101100_01111110_1;
      patterns[53935] = 25'b11010010_10101101_01111111_1;
      patterns[53936] = 25'b11010010_10101110_10000000_1;
      patterns[53937] = 25'b11010010_10101111_10000001_1;
      patterns[53938] = 25'b11010010_10110000_10000010_1;
      patterns[53939] = 25'b11010010_10110001_10000011_1;
      patterns[53940] = 25'b11010010_10110010_10000100_1;
      patterns[53941] = 25'b11010010_10110011_10000101_1;
      patterns[53942] = 25'b11010010_10110100_10000110_1;
      patterns[53943] = 25'b11010010_10110101_10000111_1;
      patterns[53944] = 25'b11010010_10110110_10001000_1;
      patterns[53945] = 25'b11010010_10110111_10001001_1;
      patterns[53946] = 25'b11010010_10111000_10001010_1;
      patterns[53947] = 25'b11010010_10111001_10001011_1;
      patterns[53948] = 25'b11010010_10111010_10001100_1;
      patterns[53949] = 25'b11010010_10111011_10001101_1;
      patterns[53950] = 25'b11010010_10111100_10001110_1;
      patterns[53951] = 25'b11010010_10111101_10001111_1;
      patterns[53952] = 25'b11010010_10111110_10010000_1;
      patterns[53953] = 25'b11010010_10111111_10010001_1;
      patterns[53954] = 25'b11010010_11000000_10010010_1;
      patterns[53955] = 25'b11010010_11000001_10010011_1;
      patterns[53956] = 25'b11010010_11000010_10010100_1;
      patterns[53957] = 25'b11010010_11000011_10010101_1;
      patterns[53958] = 25'b11010010_11000100_10010110_1;
      patterns[53959] = 25'b11010010_11000101_10010111_1;
      patterns[53960] = 25'b11010010_11000110_10011000_1;
      patterns[53961] = 25'b11010010_11000111_10011001_1;
      patterns[53962] = 25'b11010010_11001000_10011010_1;
      patterns[53963] = 25'b11010010_11001001_10011011_1;
      patterns[53964] = 25'b11010010_11001010_10011100_1;
      patterns[53965] = 25'b11010010_11001011_10011101_1;
      patterns[53966] = 25'b11010010_11001100_10011110_1;
      patterns[53967] = 25'b11010010_11001101_10011111_1;
      patterns[53968] = 25'b11010010_11001110_10100000_1;
      patterns[53969] = 25'b11010010_11001111_10100001_1;
      patterns[53970] = 25'b11010010_11010000_10100010_1;
      patterns[53971] = 25'b11010010_11010001_10100011_1;
      patterns[53972] = 25'b11010010_11010010_10100100_1;
      patterns[53973] = 25'b11010010_11010011_10100101_1;
      patterns[53974] = 25'b11010010_11010100_10100110_1;
      patterns[53975] = 25'b11010010_11010101_10100111_1;
      patterns[53976] = 25'b11010010_11010110_10101000_1;
      patterns[53977] = 25'b11010010_11010111_10101001_1;
      patterns[53978] = 25'b11010010_11011000_10101010_1;
      patterns[53979] = 25'b11010010_11011001_10101011_1;
      patterns[53980] = 25'b11010010_11011010_10101100_1;
      patterns[53981] = 25'b11010010_11011011_10101101_1;
      patterns[53982] = 25'b11010010_11011100_10101110_1;
      patterns[53983] = 25'b11010010_11011101_10101111_1;
      patterns[53984] = 25'b11010010_11011110_10110000_1;
      patterns[53985] = 25'b11010010_11011111_10110001_1;
      patterns[53986] = 25'b11010010_11100000_10110010_1;
      patterns[53987] = 25'b11010010_11100001_10110011_1;
      patterns[53988] = 25'b11010010_11100010_10110100_1;
      patterns[53989] = 25'b11010010_11100011_10110101_1;
      patterns[53990] = 25'b11010010_11100100_10110110_1;
      patterns[53991] = 25'b11010010_11100101_10110111_1;
      patterns[53992] = 25'b11010010_11100110_10111000_1;
      patterns[53993] = 25'b11010010_11100111_10111001_1;
      patterns[53994] = 25'b11010010_11101000_10111010_1;
      patterns[53995] = 25'b11010010_11101001_10111011_1;
      patterns[53996] = 25'b11010010_11101010_10111100_1;
      patterns[53997] = 25'b11010010_11101011_10111101_1;
      patterns[53998] = 25'b11010010_11101100_10111110_1;
      patterns[53999] = 25'b11010010_11101101_10111111_1;
      patterns[54000] = 25'b11010010_11101110_11000000_1;
      patterns[54001] = 25'b11010010_11101111_11000001_1;
      patterns[54002] = 25'b11010010_11110000_11000010_1;
      patterns[54003] = 25'b11010010_11110001_11000011_1;
      patterns[54004] = 25'b11010010_11110010_11000100_1;
      patterns[54005] = 25'b11010010_11110011_11000101_1;
      patterns[54006] = 25'b11010010_11110100_11000110_1;
      patterns[54007] = 25'b11010010_11110101_11000111_1;
      patterns[54008] = 25'b11010010_11110110_11001000_1;
      patterns[54009] = 25'b11010010_11110111_11001001_1;
      patterns[54010] = 25'b11010010_11111000_11001010_1;
      patterns[54011] = 25'b11010010_11111001_11001011_1;
      patterns[54012] = 25'b11010010_11111010_11001100_1;
      patterns[54013] = 25'b11010010_11111011_11001101_1;
      patterns[54014] = 25'b11010010_11111100_11001110_1;
      patterns[54015] = 25'b11010010_11111101_11001111_1;
      patterns[54016] = 25'b11010010_11111110_11010000_1;
      patterns[54017] = 25'b11010010_11111111_11010001_1;
      patterns[54018] = 25'b11010011_00000000_11010011_0;
      patterns[54019] = 25'b11010011_00000001_11010100_0;
      patterns[54020] = 25'b11010011_00000010_11010101_0;
      patterns[54021] = 25'b11010011_00000011_11010110_0;
      patterns[54022] = 25'b11010011_00000100_11010111_0;
      patterns[54023] = 25'b11010011_00000101_11011000_0;
      patterns[54024] = 25'b11010011_00000110_11011001_0;
      patterns[54025] = 25'b11010011_00000111_11011010_0;
      patterns[54026] = 25'b11010011_00001000_11011011_0;
      patterns[54027] = 25'b11010011_00001001_11011100_0;
      patterns[54028] = 25'b11010011_00001010_11011101_0;
      patterns[54029] = 25'b11010011_00001011_11011110_0;
      patterns[54030] = 25'b11010011_00001100_11011111_0;
      patterns[54031] = 25'b11010011_00001101_11100000_0;
      patterns[54032] = 25'b11010011_00001110_11100001_0;
      patterns[54033] = 25'b11010011_00001111_11100010_0;
      patterns[54034] = 25'b11010011_00010000_11100011_0;
      patterns[54035] = 25'b11010011_00010001_11100100_0;
      patterns[54036] = 25'b11010011_00010010_11100101_0;
      patterns[54037] = 25'b11010011_00010011_11100110_0;
      patterns[54038] = 25'b11010011_00010100_11100111_0;
      patterns[54039] = 25'b11010011_00010101_11101000_0;
      patterns[54040] = 25'b11010011_00010110_11101001_0;
      patterns[54041] = 25'b11010011_00010111_11101010_0;
      patterns[54042] = 25'b11010011_00011000_11101011_0;
      patterns[54043] = 25'b11010011_00011001_11101100_0;
      patterns[54044] = 25'b11010011_00011010_11101101_0;
      patterns[54045] = 25'b11010011_00011011_11101110_0;
      patterns[54046] = 25'b11010011_00011100_11101111_0;
      patterns[54047] = 25'b11010011_00011101_11110000_0;
      patterns[54048] = 25'b11010011_00011110_11110001_0;
      patterns[54049] = 25'b11010011_00011111_11110010_0;
      patterns[54050] = 25'b11010011_00100000_11110011_0;
      patterns[54051] = 25'b11010011_00100001_11110100_0;
      patterns[54052] = 25'b11010011_00100010_11110101_0;
      patterns[54053] = 25'b11010011_00100011_11110110_0;
      patterns[54054] = 25'b11010011_00100100_11110111_0;
      patterns[54055] = 25'b11010011_00100101_11111000_0;
      patterns[54056] = 25'b11010011_00100110_11111001_0;
      patterns[54057] = 25'b11010011_00100111_11111010_0;
      patterns[54058] = 25'b11010011_00101000_11111011_0;
      patterns[54059] = 25'b11010011_00101001_11111100_0;
      patterns[54060] = 25'b11010011_00101010_11111101_0;
      patterns[54061] = 25'b11010011_00101011_11111110_0;
      patterns[54062] = 25'b11010011_00101100_11111111_0;
      patterns[54063] = 25'b11010011_00101101_00000000_1;
      patterns[54064] = 25'b11010011_00101110_00000001_1;
      patterns[54065] = 25'b11010011_00101111_00000010_1;
      patterns[54066] = 25'b11010011_00110000_00000011_1;
      patterns[54067] = 25'b11010011_00110001_00000100_1;
      patterns[54068] = 25'b11010011_00110010_00000101_1;
      patterns[54069] = 25'b11010011_00110011_00000110_1;
      patterns[54070] = 25'b11010011_00110100_00000111_1;
      patterns[54071] = 25'b11010011_00110101_00001000_1;
      patterns[54072] = 25'b11010011_00110110_00001001_1;
      patterns[54073] = 25'b11010011_00110111_00001010_1;
      patterns[54074] = 25'b11010011_00111000_00001011_1;
      patterns[54075] = 25'b11010011_00111001_00001100_1;
      patterns[54076] = 25'b11010011_00111010_00001101_1;
      patterns[54077] = 25'b11010011_00111011_00001110_1;
      patterns[54078] = 25'b11010011_00111100_00001111_1;
      patterns[54079] = 25'b11010011_00111101_00010000_1;
      patterns[54080] = 25'b11010011_00111110_00010001_1;
      patterns[54081] = 25'b11010011_00111111_00010010_1;
      patterns[54082] = 25'b11010011_01000000_00010011_1;
      patterns[54083] = 25'b11010011_01000001_00010100_1;
      patterns[54084] = 25'b11010011_01000010_00010101_1;
      patterns[54085] = 25'b11010011_01000011_00010110_1;
      patterns[54086] = 25'b11010011_01000100_00010111_1;
      patterns[54087] = 25'b11010011_01000101_00011000_1;
      patterns[54088] = 25'b11010011_01000110_00011001_1;
      patterns[54089] = 25'b11010011_01000111_00011010_1;
      patterns[54090] = 25'b11010011_01001000_00011011_1;
      patterns[54091] = 25'b11010011_01001001_00011100_1;
      patterns[54092] = 25'b11010011_01001010_00011101_1;
      patterns[54093] = 25'b11010011_01001011_00011110_1;
      patterns[54094] = 25'b11010011_01001100_00011111_1;
      patterns[54095] = 25'b11010011_01001101_00100000_1;
      patterns[54096] = 25'b11010011_01001110_00100001_1;
      patterns[54097] = 25'b11010011_01001111_00100010_1;
      patterns[54098] = 25'b11010011_01010000_00100011_1;
      patterns[54099] = 25'b11010011_01010001_00100100_1;
      patterns[54100] = 25'b11010011_01010010_00100101_1;
      patterns[54101] = 25'b11010011_01010011_00100110_1;
      patterns[54102] = 25'b11010011_01010100_00100111_1;
      patterns[54103] = 25'b11010011_01010101_00101000_1;
      patterns[54104] = 25'b11010011_01010110_00101001_1;
      patterns[54105] = 25'b11010011_01010111_00101010_1;
      patterns[54106] = 25'b11010011_01011000_00101011_1;
      patterns[54107] = 25'b11010011_01011001_00101100_1;
      patterns[54108] = 25'b11010011_01011010_00101101_1;
      patterns[54109] = 25'b11010011_01011011_00101110_1;
      patterns[54110] = 25'b11010011_01011100_00101111_1;
      patterns[54111] = 25'b11010011_01011101_00110000_1;
      patterns[54112] = 25'b11010011_01011110_00110001_1;
      patterns[54113] = 25'b11010011_01011111_00110010_1;
      patterns[54114] = 25'b11010011_01100000_00110011_1;
      patterns[54115] = 25'b11010011_01100001_00110100_1;
      patterns[54116] = 25'b11010011_01100010_00110101_1;
      patterns[54117] = 25'b11010011_01100011_00110110_1;
      patterns[54118] = 25'b11010011_01100100_00110111_1;
      patterns[54119] = 25'b11010011_01100101_00111000_1;
      patterns[54120] = 25'b11010011_01100110_00111001_1;
      patterns[54121] = 25'b11010011_01100111_00111010_1;
      patterns[54122] = 25'b11010011_01101000_00111011_1;
      patterns[54123] = 25'b11010011_01101001_00111100_1;
      patterns[54124] = 25'b11010011_01101010_00111101_1;
      patterns[54125] = 25'b11010011_01101011_00111110_1;
      patterns[54126] = 25'b11010011_01101100_00111111_1;
      patterns[54127] = 25'b11010011_01101101_01000000_1;
      patterns[54128] = 25'b11010011_01101110_01000001_1;
      patterns[54129] = 25'b11010011_01101111_01000010_1;
      patterns[54130] = 25'b11010011_01110000_01000011_1;
      patterns[54131] = 25'b11010011_01110001_01000100_1;
      patterns[54132] = 25'b11010011_01110010_01000101_1;
      patterns[54133] = 25'b11010011_01110011_01000110_1;
      patterns[54134] = 25'b11010011_01110100_01000111_1;
      patterns[54135] = 25'b11010011_01110101_01001000_1;
      patterns[54136] = 25'b11010011_01110110_01001001_1;
      patterns[54137] = 25'b11010011_01110111_01001010_1;
      patterns[54138] = 25'b11010011_01111000_01001011_1;
      patterns[54139] = 25'b11010011_01111001_01001100_1;
      patterns[54140] = 25'b11010011_01111010_01001101_1;
      patterns[54141] = 25'b11010011_01111011_01001110_1;
      patterns[54142] = 25'b11010011_01111100_01001111_1;
      patterns[54143] = 25'b11010011_01111101_01010000_1;
      patterns[54144] = 25'b11010011_01111110_01010001_1;
      patterns[54145] = 25'b11010011_01111111_01010010_1;
      patterns[54146] = 25'b11010011_10000000_01010011_1;
      patterns[54147] = 25'b11010011_10000001_01010100_1;
      patterns[54148] = 25'b11010011_10000010_01010101_1;
      patterns[54149] = 25'b11010011_10000011_01010110_1;
      patterns[54150] = 25'b11010011_10000100_01010111_1;
      patterns[54151] = 25'b11010011_10000101_01011000_1;
      patterns[54152] = 25'b11010011_10000110_01011001_1;
      patterns[54153] = 25'b11010011_10000111_01011010_1;
      patterns[54154] = 25'b11010011_10001000_01011011_1;
      patterns[54155] = 25'b11010011_10001001_01011100_1;
      patterns[54156] = 25'b11010011_10001010_01011101_1;
      patterns[54157] = 25'b11010011_10001011_01011110_1;
      patterns[54158] = 25'b11010011_10001100_01011111_1;
      patterns[54159] = 25'b11010011_10001101_01100000_1;
      patterns[54160] = 25'b11010011_10001110_01100001_1;
      patterns[54161] = 25'b11010011_10001111_01100010_1;
      patterns[54162] = 25'b11010011_10010000_01100011_1;
      patterns[54163] = 25'b11010011_10010001_01100100_1;
      patterns[54164] = 25'b11010011_10010010_01100101_1;
      patterns[54165] = 25'b11010011_10010011_01100110_1;
      patterns[54166] = 25'b11010011_10010100_01100111_1;
      patterns[54167] = 25'b11010011_10010101_01101000_1;
      patterns[54168] = 25'b11010011_10010110_01101001_1;
      patterns[54169] = 25'b11010011_10010111_01101010_1;
      patterns[54170] = 25'b11010011_10011000_01101011_1;
      patterns[54171] = 25'b11010011_10011001_01101100_1;
      patterns[54172] = 25'b11010011_10011010_01101101_1;
      patterns[54173] = 25'b11010011_10011011_01101110_1;
      patterns[54174] = 25'b11010011_10011100_01101111_1;
      patterns[54175] = 25'b11010011_10011101_01110000_1;
      patterns[54176] = 25'b11010011_10011110_01110001_1;
      patterns[54177] = 25'b11010011_10011111_01110010_1;
      patterns[54178] = 25'b11010011_10100000_01110011_1;
      patterns[54179] = 25'b11010011_10100001_01110100_1;
      patterns[54180] = 25'b11010011_10100010_01110101_1;
      patterns[54181] = 25'b11010011_10100011_01110110_1;
      patterns[54182] = 25'b11010011_10100100_01110111_1;
      patterns[54183] = 25'b11010011_10100101_01111000_1;
      patterns[54184] = 25'b11010011_10100110_01111001_1;
      patterns[54185] = 25'b11010011_10100111_01111010_1;
      patterns[54186] = 25'b11010011_10101000_01111011_1;
      patterns[54187] = 25'b11010011_10101001_01111100_1;
      patterns[54188] = 25'b11010011_10101010_01111101_1;
      patterns[54189] = 25'b11010011_10101011_01111110_1;
      patterns[54190] = 25'b11010011_10101100_01111111_1;
      patterns[54191] = 25'b11010011_10101101_10000000_1;
      patterns[54192] = 25'b11010011_10101110_10000001_1;
      patterns[54193] = 25'b11010011_10101111_10000010_1;
      patterns[54194] = 25'b11010011_10110000_10000011_1;
      patterns[54195] = 25'b11010011_10110001_10000100_1;
      patterns[54196] = 25'b11010011_10110010_10000101_1;
      patterns[54197] = 25'b11010011_10110011_10000110_1;
      patterns[54198] = 25'b11010011_10110100_10000111_1;
      patterns[54199] = 25'b11010011_10110101_10001000_1;
      patterns[54200] = 25'b11010011_10110110_10001001_1;
      patterns[54201] = 25'b11010011_10110111_10001010_1;
      patterns[54202] = 25'b11010011_10111000_10001011_1;
      patterns[54203] = 25'b11010011_10111001_10001100_1;
      patterns[54204] = 25'b11010011_10111010_10001101_1;
      patterns[54205] = 25'b11010011_10111011_10001110_1;
      patterns[54206] = 25'b11010011_10111100_10001111_1;
      patterns[54207] = 25'b11010011_10111101_10010000_1;
      patterns[54208] = 25'b11010011_10111110_10010001_1;
      patterns[54209] = 25'b11010011_10111111_10010010_1;
      patterns[54210] = 25'b11010011_11000000_10010011_1;
      patterns[54211] = 25'b11010011_11000001_10010100_1;
      patterns[54212] = 25'b11010011_11000010_10010101_1;
      patterns[54213] = 25'b11010011_11000011_10010110_1;
      patterns[54214] = 25'b11010011_11000100_10010111_1;
      patterns[54215] = 25'b11010011_11000101_10011000_1;
      patterns[54216] = 25'b11010011_11000110_10011001_1;
      patterns[54217] = 25'b11010011_11000111_10011010_1;
      patterns[54218] = 25'b11010011_11001000_10011011_1;
      patterns[54219] = 25'b11010011_11001001_10011100_1;
      patterns[54220] = 25'b11010011_11001010_10011101_1;
      patterns[54221] = 25'b11010011_11001011_10011110_1;
      patterns[54222] = 25'b11010011_11001100_10011111_1;
      patterns[54223] = 25'b11010011_11001101_10100000_1;
      patterns[54224] = 25'b11010011_11001110_10100001_1;
      patterns[54225] = 25'b11010011_11001111_10100010_1;
      patterns[54226] = 25'b11010011_11010000_10100011_1;
      patterns[54227] = 25'b11010011_11010001_10100100_1;
      patterns[54228] = 25'b11010011_11010010_10100101_1;
      patterns[54229] = 25'b11010011_11010011_10100110_1;
      patterns[54230] = 25'b11010011_11010100_10100111_1;
      patterns[54231] = 25'b11010011_11010101_10101000_1;
      patterns[54232] = 25'b11010011_11010110_10101001_1;
      patterns[54233] = 25'b11010011_11010111_10101010_1;
      patterns[54234] = 25'b11010011_11011000_10101011_1;
      patterns[54235] = 25'b11010011_11011001_10101100_1;
      patterns[54236] = 25'b11010011_11011010_10101101_1;
      patterns[54237] = 25'b11010011_11011011_10101110_1;
      patterns[54238] = 25'b11010011_11011100_10101111_1;
      patterns[54239] = 25'b11010011_11011101_10110000_1;
      patterns[54240] = 25'b11010011_11011110_10110001_1;
      patterns[54241] = 25'b11010011_11011111_10110010_1;
      patterns[54242] = 25'b11010011_11100000_10110011_1;
      patterns[54243] = 25'b11010011_11100001_10110100_1;
      patterns[54244] = 25'b11010011_11100010_10110101_1;
      patterns[54245] = 25'b11010011_11100011_10110110_1;
      patterns[54246] = 25'b11010011_11100100_10110111_1;
      patterns[54247] = 25'b11010011_11100101_10111000_1;
      patterns[54248] = 25'b11010011_11100110_10111001_1;
      patterns[54249] = 25'b11010011_11100111_10111010_1;
      patterns[54250] = 25'b11010011_11101000_10111011_1;
      patterns[54251] = 25'b11010011_11101001_10111100_1;
      patterns[54252] = 25'b11010011_11101010_10111101_1;
      patterns[54253] = 25'b11010011_11101011_10111110_1;
      patterns[54254] = 25'b11010011_11101100_10111111_1;
      patterns[54255] = 25'b11010011_11101101_11000000_1;
      patterns[54256] = 25'b11010011_11101110_11000001_1;
      patterns[54257] = 25'b11010011_11101111_11000010_1;
      patterns[54258] = 25'b11010011_11110000_11000011_1;
      patterns[54259] = 25'b11010011_11110001_11000100_1;
      patterns[54260] = 25'b11010011_11110010_11000101_1;
      patterns[54261] = 25'b11010011_11110011_11000110_1;
      patterns[54262] = 25'b11010011_11110100_11000111_1;
      patterns[54263] = 25'b11010011_11110101_11001000_1;
      patterns[54264] = 25'b11010011_11110110_11001001_1;
      patterns[54265] = 25'b11010011_11110111_11001010_1;
      patterns[54266] = 25'b11010011_11111000_11001011_1;
      patterns[54267] = 25'b11010011_11111001_11001100_1;
      patterns[54268] = 25'b11010011_11111010_11001101_1;
      patterns[54269] = 25'b11010011_11111011_11001110_1;
      patterns[54270] = 25'b11010011_11111100_11001111_1;
      patterns[54271] = 25'b11010011_11111101_11010000_1;
      patterns[54272] = 25'b11010011_11111110_11010001_1;
      patterns[54273] = 25'b11010011_11111111_11010010_1;
      patterns[54274] = 25'b11010100_00000000_11010100_0;
      patterns[54275] = 25'b11010100_00000001_11010101_0;
      patterns[54276] = 25'b11010100_00000010_11010110_0;
      patterns[54277] = 25'b11010100_00000011_11010111_0;
      patterns[54278] = 25'b11010100_00000100_11011000_0;
      patterns[54279] = 25'b11010100_00000101_11011001_0;
      patterns[54280] = 25'b11010100_00000110_11011010_0;
      patterns[54281] = 25'b11010100_00000111_11011011_0;
      patterns[54282] = 25'b11010100_00001000_11011100_0;
      patterns[54283] = 25'b11010100_00001001_11011101_0;
      patterns[54284] = 25'b11010100_00001010_11011110_0;
      patterns[54285] = 25'b11010100_00001011_11011111_0;
      patterns[54286] = 25'b11010100_00001100_11100000_0;
      patterns[54287] = 25'b11010100_00001101_11100001_0;
      patterns[54288] = 25'b11010100_00001110_11100010_0;
      patterns[54289] = 25'b11010100_00001111_11100011_0;
      patterns[54290] = 25'b11010100_00010000_11100100_0;
      patterns[54291] = 25'b11010100_00010001_11100101_0;
      patterns[54292] = 25'b11010100_00010010_11100110_0;
      patterns[54293] = 25'b11010100_00010011_11100111_0;
      patterns[54294] = 25'b11010100_00010100_11101000_0;
      patterns[54295] = 25'b11010100_00010101_11101001_0;
      patterns[54296] = 25'b11010100_00010110_11101010_0;
      patterns[54297] = 25'b11010100_00010111_11101011_0;
      patterns[54298] = 25'b11010100_00011000_11101100_0;
      patterns[54299] = 25'b11010100_00011001_11101101_0;
      patterns[54300] = 25'b11010100_00011010_11101110_0;
      patterns[54301] = 25'b11010100_00011011_11101111_0;
      patterns[54302] = 25'b11010100_00011100_11110000_0;
      patterns[54303] = 25'b11010100_00011101_11110001_0;
      patterns[54304] = 25'b11010100_00011110_11110010_0;
      patterns[54305] = 25'b11010100_00011111_11110011_0;
      patterns[54306] = 25'b11010100_00100000_11110100_0;
      patterns[54307] = 25'b11010100_00100001_11110101_0;
      patterns[54308] = 25'b11010100_00100010_11110110_0;
      patterns[54309] = 25'b11010100_00100011_11110111_0;
      patterns[54310] = 25'b11010100_00100100_11111000_0;
      patterns[54311] = 25'b11010100_00100101_11111001_0;
      patterns[54312] = 25'b11010100_00100110_11111010_0;
      patterns[54313] = 25'b11010100_00100111_11111011_0;
      patterns[54314] = 25'b11010100_00101000_11111100_0;
      patterns[54315] = 25'b11010100_00101001_11111101_0;
      patterns[54316] = 25'b11010100_00101010_11111110_0;
      patterns[54317] = 25'b11010100_00101011_11111111_0;
      patterns[54318] = 25'b11010100_00101100_00000000_1;
      patterns[54319] = 25'b11010100_00101101_00000001_1;
      patterns[54320] = 25'b11010100_00101110_00000010_1;
      patterns[54321] = 25'b11010100_00101111_00000011_1;
      patterns[54322] = 25'b11010100_00110000_00000100_1;
      patterns[54323] = 25'b11010100_00110001_00000101_1;
      patterns[54324] = 25'b11010100_00110010_00000110_1;
      patterns[54325] = 25'b11010100_00110011_00000111_1;
      patterns[54326] = 25'b11010100_00110100_00001000_1;
      patterns[54327] = 25'b11010100_00110101_00001001_1;
      patterns[54328] = 25'b11010100_00110110_00001010_1;
      patterns[54329] = 25'b11010100_00110111_00001011_1;
      patterns[54330] = 25'b11010100_00111000_00001100_1;
      patterns[54331] = 25'b11010100_00111001_00001101_1;
      patterns[54332] = 25'b11010100_00111010_00001110_1;
      patterns[54333] = 25'b11010100_00111011_00001111_1;
      patterns[54334] = 25'b11010100_00111100_00010000_1;
      patterns[54335] = 25'b11010100_00111101_00010001_1;
      patterns[54336] = 25'b11010100_00111110_00010010_1;
      patterns[54337] = 25'b11010100_00111111_00010011_1;
      patterns[54338] = 25'b11010100_01000000_00010100_1;
      patterns[54339] = 25'b11010100_01000001_00010101_1;
      patterns[54340] = 25'b11010100_01000010_00010110_1;
      patterns[54341] = 25'b11010100_01000011_00010111_1;
      patterns[54342] = 25'b11010100_01000100_00011000_1;
      patterns[54343] = 25'b11010100_01000101_00011001_1;
      patterns[54344] = 25'b11010100_01000110_00011010_1;
      patterns[54345] = 25'b11010100_01000111_00011011_1;
      patterns[54346] = 25'b11010100_01001000_00011100_1;
      patterns[54347] = 25'b11010100_01001001_00011101_1;
      patterns[54348] = 25'b11010100_01001010_00011110_1;
      patterns[54349] = 25'b11010100_01001011_00011111_1;
      patterns[54350] = 25'b11010100_01001100_00100000_1;
      patterns[54351] = 25'b11010100_01001101_00100001_1;
      patterns[54352] = 25'b11010100_01001110_00100010_1;
      patterns[54353] = 25'b11010100_01001111_00100011_1;
      patterns[54354] = 25'b11010100_01010000_00100100_1;
      patterns[54355] = 25'b11010100_01010001_00100101_1;
      patterns[54356] = 25'b11010100_01010010_00100110_1;
      patterns[54357] = 25'b11010100_01010011_00100111_1;
      patterns[54358] = 25'b11010100_01010100_00101000_1;
      patterns[54359] = 25'b11010100_01010101_00101001_1;
      patterns[54360] = 25'b11010100_01010110_00101010_1;
      patterns[54361] = 25'b11010100_01010111_00101011_1;
      patterns[54362] = 25'b11010100_01011000_00101100_1;
      patterns[54363] = 25'b11010100_01011001_00101101_1;
      patterns[54364] = 25'b11010100_01011010_00101110_1;
      patterns[54365] = 25'b11010100_01011011_00101111_1;
      patterns[54366] = 25'b11010100_01011100_00110000_1;
      patterns[54367] = 25'b11010100_01011101_00110001_1;
      patterns[54368] = 25'b11010100_01011110_00110010_1;
      patterns[54369] = 25'b11010100_01011111_00110011_1;
      patterns[54370] = 25'b11010100_01100000_00110100_1;
      patterns[54371] = 25'b11010100_01100001_00110101_1;
      patterns[54372] = 25'b11010100_01100010_00110110_1;
      patterns[54373] = 25'b11010100_01100011_00110111_1;
      patterns[54374] = 25'b11010100_01100100_00111000_1;
      patterns[54375] = 25'b11010100_01100101_00111001_1;
      patterns[54376] = 25'b11010100_01100110_00111010_1;
      patterns[54377] = 25'b11010100_01100111_00111011_1;
      patterns[54378] = 25'b11010100_01101000_00111100_1;
      patterns[54379] = 25'b11010100_01101001_00111101_1;
      patterns[54380] = 25'b11010100_01101010_00111110_1;
      patterns[54381] = 25'b11010100_01101011_00111111_1;
      patterns[54382] = 25'b11010100_01101100_01000000_1;
      patterns[54383] = 25'b11010100_01101101_01000001_1;
      patterns[54384] = 25'b11010100_01101110_01000010_1;
      patterns[54385] = 25'b11010100_01101111_01000011_1;
      patterns[54386] = 25'b11010100_01110000_01000100_1;
      patterns[54387] = 25'b11010100_01110001_01000101_1;
      patterns[54388] = 25'b11010100_01110010_01000110_1;
      patterns[54389] = 25'b11010100_01110011_01000111_1;
      patterns[54390] = 25'b11010100_01110100_01001000_1;
      patterns[54391] = 25'b11010100_01110101_01001001_1;
      patterns[54392] = 25'b11010100_01110110_01001010_1;
      patterns[54393] = 25'b11010100_01110111_01001011_1;
      patterns[54394] = 25'b11010100_01111000_01001100_1;
      patterns[54395] = 25'b11010100_01111001_01001101_1;
      patterns[54396] = 25'b11010100_01111010_01001110_1;
      patterns[54397] = 25'b11010100_01111011_01001111_1;
      patterns[54398] = 25'b11010100_01111100_01010000_1;
      patterns[54399] = 25'b11010100_01111101_01010001_1;
      patterns[54400] = 25'b11010100_01111110_01010010_1;
      patterns[54401] = 25'b11010100_01111111_01010011_1;
      patterns[54402] = 25'b11010100_10000000_01010100_1;
      patterns[54403] = 25'b11010100_10000001_01010101_1;
      patterns[54404] = 25'b11010100_10000010_01010110_1;
      patterns[54405] = 25'b11010100_10000011_01010111_1;
      patterns[54406] = 25'b11010100_10000100_01011000_1;
      patterns[54407] = 25'b11010100_10000101_01011001_1;
      patterns[54408] = 25'b11010100_10000110_01011010_1;
      patterns[54409] = 25'b11010100_10000111_01011011_1;
      patterns[54410] = 25'b11010100_10001000_01011100_1;
      patterns[54411] = 25'b11010100_10001001_01011101_1;
      patterns[54412] = 25'b11010100_10001010_01011110_1;
      patterns[54413] = 25'b11010100_10001011_01011111_1;
      patterns[54414] = 25'b11010100_10001100_01100000_1;
      patterns[54415] = 25'b11010100_10001101_01100001_1;
      patterns[54416] = 25'b11010100_10001110_01100010_1;
      patterns[54417] = 25'b11010100_10001111_01100011_1;
      patterns[54418] = 25'b11010100_10010000_01100100_1;
      patterns[54419] = 25'b11010100_10010001_01100101_1;
      patterns[54420] = 25'b11010100_10010010_01100110_1;
      patterns[54421] = 25'b11010100_10010011_01100111_1;
      patterns[54422] = 25'b11010100_10010100_01101000_1;
      patterns[54423] = 25'b11010100_10010101_01101001_1;
      patterns[54424] = 25'b11010100_10010110_01101010_1;
      patterns[54425] = 25'b11010100_10010111_01101011_1;
      patterns[54426] = 25'b11010100_10011000_01101100_1;
      patterns[54427] = 25'b11010100_10011001_01101101_1;
      patterns[54428] = 25'b11010100_10011010_01101110_1;
      patterns[54429] = 25'b11010100_10011011_01101111_1;
      patterns[54430] = 25'b11010100_10011100_01110000_1;
      patterns[54431] = 25'b11010100_10011101_01110001_1;
      patterns[54432] = 25'b11010100_10011110_01110010_1;
      patterns[54433] = 25'b11010100_10011111_01110011_1;
      patterns[54434] = 25'b11010100_10100000_01110100_1;
      patterns[54435] = 25'b11010100_10100001_01110101_1;
      patterns[54436] = 25'b11010100_10100010_01110110_1;
      patterns[54437] = 25'b11010100_10100011_01110111_1;
      patterns[54438] = 25'b11010100_10100100_01111000_1;
      patterns[54439] = 25'b11010100_10100101_01111001_1;
      patterns[54440] = 25'b11010100_10100110_01111010_1;
      patterns[54441] = 25'b11010100_10100111_01111011_1;
      patterns[54442] = 25'b11010100_10101000_01111100_1;
      patterns[54443] = 25'b11010100_10101001_01111101_1;
      patterns[54444] = 25'b11010100_10101010_01111110_1;
      patterns[54445] = 25'b11010100_10101011_01111111_1;
      patterns[54446] = 25'b11010100_10101100_10000000_1;
      patterns[54447] = 25'b11010100_10101101_10000001_1;
      patterns[54448] = 25'b11010100_10101110_10000010_1;
      patterns[54449] = 25'b11010100_10101111_10000011_1;
      patterns[54450] = 25'b11010100_10110000_10000100_1;
      patterns[54451] = 25'b11010100_10110001_10000101_1;
      patterns[54452] = 25'b11010100_10110010_10000110_1;
      patterns[54453] = 25'b11010100_10110011_10000111_1;
      patterns[54454] = 25'b11010100_10110100_10001000_1;
      patterns[54455] = 25'b11010100_10110101_10001001_1;
      patterns[54456] = 25'b11010100_10110110_10001010_1;
      patterns[54457] = 25'b11010100_10110111_10001011_1;
      patterns[54458] = 25'b11010100_10111000_10001100_1;
      patterns[54459] = 25'b11010100_10111001_10001101_1;
      patterns[54460] = 25'b11010100_10111010_10001110_1;
      patterns[54461] = 25'b11010100_10111011_10001111_1;
      patterns[54462] = 25'b11010100_10111100_10010000_1;
      patterns[54463] = 25'b11010100_10111101_10010001_1;
      patterns[54464] = 25'b11010100_10111110_10010010_1;
      patterns[54465] = 25'b11010100_10111111_10010011_1;
      patterns[54466] = 25'b11010100_11000000_10010100_1;
      patterns[54467] = 25'b11010100_11000001_10010101_1;
      patterns[54468] = 25'b11010100_11000010_10010110_1;
      patterns[54469] = 25'b11010100_11000011_10010111_1;
      patterns[54470] = 25'b11010100_11000100_10011000_1;
      patterns[54471] = 25'b11010100_11000101_10011001_1;
      patterns[54472] = 25'b11010100_11000110_10011010_1;
      patterns[54473] = 25'b11010100_11000111_10011011_1;
      patterns[54474] = 25'b11010100_11001000_10011100_1;
      patterns[54475] = 25'b11010100_11001001_10011101_1;
      patterns[54476] = 25'b11010100_11001010_10011110_1;
      patterns[54477] = 25'b11010100_11001011_10011111_1;
      patterns[54478] = 25'b11010100_11001100_10100000_1;
      patterns[54479] = 25'b11010100_11001101_10100001_1;
      patterns[54480] = 25'b11010100_11001110_10100010_1;
      patterns[54481] = 25'b11010100_11001111_10100011_1;
      patterns[54482] = 25'b11010100_11010000_10100100_1;
      patterns[54483] = 25'b11010100_11010001_10100101_1;
      patterns[54484] = 25'b11010100_11010010_10100110_1;
      patterns[54485] = 25'b11010100_11010011_10100111_1;
      patterns[54486] = 25'b11010100_11010100_10101000_1;
      patterns[54487] = 25'b11010100_11010101_10101001_1;
      patterns[54488] = 25'b11010100_11010110_10101010_1;
      patterns[54489] = 25'b11010100_11010111_10101011_1;
      patterns[54490] = 25'b11010100_11011000_10101100_1;
      patterns[54491] = 25'b11010100_11011001_10101101_1;
      patterns[54492] = 25'b11010100_11011010_10101110_1;
      patterns[54493] = 25'b11010100_11011011_10101111_1;
      patterns[54494] = 25'b11010100_11011100_10110000_1;
      patterns[54495] = 25'b11010100_11011101_10110001_1;
      patterns[54496] = 25'b11010100_11011110_10110010_1;
      patterns[54497] = 25'b11010100_11011111_10110011_1;
      patterns[54498] = 25'b11010100_11100000_10110100_1;
      patterns[54499] = 25'b11010100_11100001_10110101_1;
      patterns[54500] = 25'b11010100_11100010_10110110_1;
      patterns[54501] = 25'b11010100_11100011_10110111_1;
      patterns[54502] = 25'b11010100_11100100_10111000_1;
      patterns[54503] = 25'b11010100_11100101_10111001_1;
      patterns[54504] = 25'b11010100_11100110_10111010_1;
      patterns[54505] = 25'b11010100_11100111_10111011_1;
      patterns[54506] = 25'b11010100_11101000_10111100_1;
      patterns[54507] = 25'b11010100_11101001_10111101_1;
      patterns[54508] = 25'b11010100_11101010_10111110_1;
      patterns[54509] = 25'b11010100_11101011_10111111_1;
      patterns[54510] = 25'b11010100_11101100_11000000_1;
      patterns[54511] = 25'b11010100_11101101_11000001_1;
      patterns[54512] = 25'b11010100_11101110_11000010_1;
      patterns[54513] = 25'b11010100_11101111_11000011_1;
      patterns[54514] = 25'b11010100_11110000_11000100_1;
      patterns[54515] = 25'b11010100_11110001_11000101_1;
      patterns[54516] = 25'b11010100_11110010_11000110_1;
      patterns[54517] = 25'b11010100_11110011_11000111_1;
      patterns[54518] = 25'b11010100_11110100_11001000_1;
      patterns[54519] = 25'b11010100_11110101_11001001_1;
      patterns[54520] = 25'b11010100_11110110_11001010_1;
      patterns[54521] = 25'b11010100_11110111_11001011_1;
      patterns[54522] = 25'b11010100_11111000_11001100_1;
      patterns[54523] = 25'b11010100_11111001_11001101_1;
      patterns[54524] = 25'b11010100_11111010_11001110_1;
      patterns[54525] = 25'b11010100_11111011_11001111_1;
      patterns[54526] = 25'b11010100_11111100_11010000_1;
      patterns[54527] = 25'b11010100_11111101_11010001_1;
      patterns[54528] = 25'b11010100_11111110_11010010_1;
      patterns[54529] = 25'b11010100_11111111_11010011_1;
      patterns[54530] = 25'b11010101_00000000_11010101_0;
      patterns[54531] = 25'b11010101_00000001_11010110_0;
      patterns[54532] = 25'b11010101_00000010_11010111_0;
      patterns[54533] = 25'b11010101_00000011_11011000_0;
      patterns[54534] = 25'b11010101_00000100_11011001_0;
      patterns[54535] = 25'b11010101_00000101_11011010_0;
      patterns[54536] = 25'b11010101_00000110_11011011_0;
      patterns[54537] = 25'b11010101_00000111_11011100_0;
      patterns[54538] = 25'b11010101_00001000_11011101_0;
      patterns[54539] = 25'b11010101_00001001_11011110_0;
      patterns[54540] = 25'b11010101_00001010_11011111_0;
      patterns[54541] = 25'b11010101_00001011_11100000_0;
      patterns[54542] = 25'b11010101_00001100_11100001_0;
      patterns[54543] = 25'b11010101_00001101_11100010_0;
      patterns[54544] = 25'b11010101_00001110_11100011_0;
      patterns[54545] = 25'b11010101_00001111_11100100_0;
      patterns[54546] = 25'b11010101_00010000_11100101_0;
      patterns[54547] = 25'b11010101_00010001_11100110_0;
      patterns[54548] = 25'b11010101_00010010_11100111_0;
      patterns[54549] = 25'b11010101_00010011_11101000_0;
      patterns[54550] = 25'b11010101_00010100_11101001_0;
      patterns[54551] = 25'b11010101_00010101_11101010_0;
      patterns[54552] = 25'b11010101_00010110_11101011_0;
      patterns[54553] = 25'b11010101_00010111_11101100_0;
      patterns[54554] = 25'b11010101_00011000_11101101_0;
      patterns[54555] = 25'b11010101_00011001_11101110_0;
      patterns[54556] = 25'b11010101_00011010_11101111_0;
      patterns[54557] = 25'b11010101_00011011_11110000_0;
      patterns[54558] = 25'b11010101_00011100_11110001_0;
      patterns[54559] = 25'b11010101_00011101_11110010_0;
      patterns[54560] = 25'b11010101_00011110_11110011_0;
      patterns[54561] = 25'b11010101_00011111_11110100_0;
      patterns[54562] = 25'b11010101_00100000_11110101_0;
      patterns[54563] = 25'b11010101_00100001_11110110_0;
      patterns[54564] = 25'b11010101_00100010_11110111_0;
      patterns[54565] = 25'b11010101_00100011_11111000_0;
      patterns[54566] = 25'b11010101_00100100_11111001_0;
      patterns[54567] = 25'b11010101_00100101_11111010_0;
      patterns[54568] = 25'b11010101_00100110_11111011_0;
      patterns[54569] = 25'b11010101_00100111_11111100_0;
      patterns[54570] = 25'b11010101_00101000_11111101_0;
      patterns[54571] = 25'b11010101_00101001_11111110_0;
      patterns[54572] = 25'b11010101_00101010_11111111_0;
      patterns[54573] = 25'b11010101_00101011_00000000_1;
      patterns[54574] = 25'b11010101_00101100_00000001_1;
      patterns[54575] = 25'b11010101_00101101_00000010_1;
      patterns[54576] = 25'b11010101_00101110_00000011_1;
      patterns[54577] = 25'b11010101_00101111_00000100_1;
      patterns[54578] = 25'b11010101_00110000_00000101_1;
      patterns[54579] = 25'b11010101_00110001_00000110_1;
      patterns[54580] = 25'b11010101_00110010_00000111_1;
      patterns[54581] = 25'b11010101_00110011_00001000_1;
      patterns[54582] = 25'b11010101_00110100_00001001_1;
      patterns[54583] = 25'b11010101_00110101_00001010_1;
      patterns[54584] = 25'b11010101_00110110_00001011_1;
      patterns[54585] = 25'b11010101_00110111_00001100_1;
      patterns[54586] = 25'b11010101_00111000_00001101_1;
      patterns[54587] = 25'b11010101_00111001_00001110_1;
      patterns[54588] = 25'b11010101_00111010_00001111_1;
      patterns[54589] = 25'b11010101_00111011_00010000_1;
      patterns[54590] = 25'b11010101_00111100_00010001_1;
      patterns[54591] = 25'b11010101_00111101_00010010_1;
      patterns[54592] = 25'b11010101_00111110_00010011_1;
      patterns[54593] = 25'b11010101_00111111_00010100_1;
      patterns[54594] = 25'b11010101_01000000_00010101_1;
      patterns[54595] = 25'b11010101_01000001_00010110_1;
      patterns[54596] = 25'b11010101_01000010_00010111_1;
      patterns[54597] = 25'b11010101_01000011_00011000_1;
      patterns[54598] = 25'b11010101_01000100_00011001_1;
      patterns[54599] = 25'b11010101_01000101_00011010_1;
      patterns[54600] = 25'b11010101_01000110_00011011_1;
      patterns[54601] = 25'b11010101_01000111_00011100_1;
      patterns[54602] = 25'b11010101_01001000_00011101_1;
      patterns[54603] = 25'b11010101_01001001_00011110_1;
      patterns[54604] = 25'b11010101_01001010_00011111_1;
      patterns[54605] = 25'b11010101_01001011_00100000_1;
      patterns[54606] = 25'b11010101_01001100_00100001_1;
      patterns[54607] = 25'b11010101_01001101_00100010_1;
      patterns[54608] = 25'b11010101_01001110_00100011_1;
      patterns[54609] = 25'b11010101_01001111_00100100_1;
      patterns[54610] = 25'b11010101_01010000_00100101_1;
      patterns[54611] = 25'b11010101_01010001_00100110_1;
      patterns[54612] = 25'b11010101_01010010_00100111_1;
      patterns[54613] = 25'b11010101_01010011_00101000_1;
      patterns[54614] = 25'b11010101_01010100_00101001_1;
      patterns[54615] = 25'b11010101_01010101_00101010_1;
      patterns[54616] = 25'b11010101_01010110_00101011_1;
      patterns[54617] = 25'b11010101_01010111_00101100_1;
      patterns[54618] = 25'b11010101_01011000_00101101_1;
      patterns[54619] = 25'b11010101_01011001_00101110_1;
      patterns[54620] = 25'b11010101_01011010_00101111_1;
      patterns[54621] = 25'b11010101_01011011_00110000_1;
      patterns[54622] = 25'b11010101_01011100_00110001_1;
      patterns[54623] = 25'b11010101_01011101_00110010_1;
      patterns[54624] = 25'b11010101_01011110_00110011_1;
      patterns[54625] = 25'b11010101_01011111_00110100_1;
      patterns[54626] = 25'b11010101_01100000_00110101_1;
      patterns[54627] = 25'b11010101_01100001_00110110_1;
      patterns[54628] = 25'b11010101_01100010_00110111_1;
      patterns[54629] = 25'b11010101_01100011_00111000_1;
      patterns[54630] = 25'b11010101_01100100_00111001_1;
      patterns[54631] = 25'b11010101_01100101_00111010_1;
      patterns[54632] = 25'b11010101_01100110_00111011_1;
      patterns[54633] = 25'b11010101_01100111_00111100_1;
      patterns[54634] = 25'b11010101_01101000_00111101_1;
      patterns[54635] = 25'b11010101_01101001_00111110_1;
      patterns[54636] = 25'b11010101_01101010_00111111_1;
      patterns[54637] = 25'b11010101_01101011_01000000_1;
      patterns[54638] = 25'b11010101_01101100_01000001_1;
      patterns[54639] = 25'b11010101_01101101_01000010_1;
      patterns[54640] = 25'b11010101_01101110_01000011_1;
      patterns[54641] = 25'b11010101_01101111_01000100_1;
      patterns[54642] = 25'b11010101_01110000_01000101_1;
      patterns[54643] = 25'b11010101_01110001_01000110_1;
      patterns[54644] = 25'b11010101_01110010_01000111_1;
      patterns[54645] = 25'b11010101_01110011_01001000_1;
      patterns[54646] = 25'b11010101_01110100_01001001_1;
      patterns[54647] = 25'b11010101_01110101_01001010_1;
      patterns[54648] = 25'b11010101_01110110_01001011_1;
      patterns[54649] = 25'b11010101_01110111_01001100_1;
      patterns[54650] = 25'b11010101_01111000_01001101_1;
      patterns[54651] = 25'b11010101_01111001_01001110_1;
      patterns[54652] = 25'b11010101_01111010_01001111_1;
      patterns[54653] = 25'b11010101_01111011_01010000_1;
      patterns[54654] = 25'b11010101_01111100_01010001_1;
      patterns[54655] = 25'b11010101_01111101_01010010_1;
      patterns[54656] = 25'b11010101_01111110_01010011_1;
      patterns[54657] = 25'b11010101_01111111_01010100_1;
      patterns[54658] = 25'b11010101_10000000_01010101_1;
      patterns[54659] = 25'b11010101_10000001_01010110_1;
      patterns[54660] = 25'b11010101_10000010_01010111_1;
      patterns[54661] = 25'b11010101_10000011_01011000_1;
      patterns[54662] = 25'b11010101_10000100_01011001_1;
      patterns[54663] = 25'b11010101_10000101_01011010_1;
      patterns[54664] = 25'b11010101_10000110_01011011_1;
      patterns[54665] = 25'b11010101_10000111_01011100_1;
      patterns[54666] = 25'b11010101_10001000_01011101_1;
      patterns[54667] = 25'b11010101_10001001_01011110_1;
      patterns[54668] = 25'b11010101_10001010_01011111_1;
      patterns[54669] = 25'b11010101_10001011_01100000_1;
      patterns[54670] = 25'b11010101_10001100_01100001_1;
      patterns[54671] = 25'b11010101_10001101_01100010_1;
      patterns[54672] = 25'b11010101_10001110_01100011_1;
      patterns[54673] = 25'b11010101_10001111_01100100_1;
      patterns[54674] = 25'b11010101_10010000_01100101_1;
      patterns[54675] = 25'b11010101_10010001_01100110_1;
      patterns[54676] = 25'b11010101_10010010_01100111_1;
      patterns[54677] = 25'b11010101_10010011_01101000_1;
      patterns[54678] = 25'b11010101_10010100_01101001_1;
      patterns[54679] = 25'b11010101_10010101_01101010_1;
      patterns[54680] = 25'b11010101_10010110_01101011_1;
      patterns[54681] = 25'b11010101_10010111_01101100_1;
      patterns[54682] = 25'b11010101_10011000_01101101_1;
      patterns[54683] = 25'b11010101_10011001_01101110_1;
      patterns[54684] = 25'b11010101_10011010_01101111_1;
      patterns[54685] = 25'b11010101_10011011_01110000_1;
      patterns[54686] = 25'b11010101_10011100_01110001_1;
      patterns[54687] = 25'b11010101_10011101_01110010_1;
      patterns[54688] = 25'b11010101_10011110_01110011_1;
      patterns[54689] = 25'b11010101_10011111_01110100_1;
      patterns[54690] = 25'b11010101_10100000_01110101_1;
      patterns[54691] = 25'b11010101_10100001_01110110_1;
      patterns[54692] = 25'b11010101_10100010_01110111_1;
      patterns[54693] = 25'b11010101_10100011_01111000_1;
      patterns[54694] = 25'b11010101_10100100_01111001_1;
      patterns[54695] = 25'b11010101_10100101_01111010_1;
      patterns[54696] = 25'b11010101_10100110_01111011_1;
      patterns[54697] = 25'b11010101_10100111_01111100_1;
      patterns[54698] = 25'b11010101_10101000_01111101_1;
      patterns[54699] = 25'b11010101_10101001_01111110_1;
      patterns[54700] = 25'b11010101_10101010_01111111_1;
      patterns[54701] = 25'b11010101_10101011_10000000_1;
      patterns[54702] = 25'b11010101_10101100_10000001_1;
      patterns[54703] = 25'b11010101_10101101_10000010_1;
      patterns[54704] = 25'b11010101_10101110_10000011_1;
      patterns[54705] = 25'b11010101_10101111_10000100_1;
      patterns[54706] = 25'b11010101_10110000_10000101_1;
      patterns[54707] = 25'b11010101_10110001_10000110_1;
      patterns[54708] = 25'b11010101_10110010_10000111_1;
      patterns[54709] = 25'b11010101_10110011_10001000_1;
      patterns[54710] = 25'b11010101_10110100_10001001_1;
      patterns[54711] = 25'b11010101_10110101_10001010_1;
      patterns[54712] = 25'b11010101_10110110_10001011_1;
      patterns[54713] = 25'b11010101_10110111_10001100_1;
      patterns[54714] = 25'b11010101_10111000_10001101_1;
      patterns[54715] = 25'b11010101_10111001_10001110_1;
      patterns[54716] = 25'b11010101_10111010_10001111_1;
      patterns[54717] = 25'b11010101_10111011_10010000_1;
      patterns[54718] = 25'b11010101_10111100_10010001_1;
      patterns[54719] = 25'b11010101_10111101_10010010_1;
      patterns[54720] = 25'b11010101_10111110_10010011_1;
      patterns[54721] = 25'b11010101_10111111_10010100_1;
      patterns[54722] = 25'b11010101_11000000_10010101_1;
      patterns[54723] = 25'b11010101_11000001_10010110_1;
      patterns[54724] = 25'b11010101_11000010_10010111_1;
      patterns[54725] = 25'b11010101_11000011_10011000_1;
      patterns[54726] = 25'b11010101_11000100_10011001_1;
      patterns[54727] = 25'b11010101_11000101_10011010_1;
      patterns[54728] = 25'b11010101_11000110_10011011_1;
      patterns[54729] = 25'b11010101_11000111_10011100_1;
      patterns[54730] = 25'b11010101_11001000_10011101_1;
      patterns[54731] = 25'b11010101_11001001_10011110_1;
      patterns[54732] = 25'b11010101_11001010_10011111_1;
      patterns[54733] = 25'b11010101_11001011_10100000_1;
      patterns[54734] = 25'b11010101_11001100_10100001_1;
      patterns[54735] = 25'b11010101_11001101_10100010_1;
      patterns[54736] = 25'b11010101_11001110_10100011_1;
      patterns[54737] = 25'b11010101_11001111_10100100_1;
      patterns[54738] = 25'b11010101_11010000_10100101_1;
      patterns[54739] = 25'b11010101_11010001_10100110_1;
      patterns[54740] = 25'b11010101_11010010_10100111_1;
      patterns[54741] = 25'b11010101_11010011_10101000_1;
      patterns[54742] = 25'b11010101_11010100_10101001_1;
      patterns[54743] = 25'b11010101_11010101_10101010_1;
      patterns[54744] = 25'b11010101_11010110_10101011_1;
      patterns[54745] = 25'b11010101_11010111_10101100_1;
      patterns[54746] = 25'b11010101_11011000_10101101_1;
      patterns[54747] = 25'b11010101_11011001_10101110_1;
      patterns[54748] = 25'b11010101_11011010_10101111_1;
      patterns[54749] = 25'b11010101_11011011_10110000_1;
      patterns[54750] = 25'b11010101_11011100_10110001_1;
      patterns[54751] = 25'b11010101_11011101_10110010_1;
      patterns[54752] = 25'b11010101_11011110_10110011_1;
      patterns[54753] = 25'b11010101_11011111_10110100_1;
      patterns[54754] = 25'b11010101_11100000_10110101_1;
      patterns[54755] = 25'b11010101_11100001_10110110_1;
      patterns[54756] = 25'b11010101_11100010_10110111_1;
      patterns[54757] = 25'b11010101_11100011_10111000_1;
      patterns[54758] = 25'b11010101_11100100_10111001_1;
      patterns[54759] = 25'b11010101_11100101_10111010_1;
      patterns[54760] = 25'b11010101_11100110_10111011_1;
      patterns[54761] = 25'b11010101_11100111_10111100_1;
      patterns[54762] = 25'b11010101_11101000_10111101_1;
      patterns[54763] = 25'b11010101_11101001_10111110_1;
      patterns[54764] = 25'b11010101_11101010_10111111_1;
      patterns[54765] = 25'b11010101_11101011_11000000_1;
      patterns[54766] = 25'b11010101_11101100_11000001_1;
      patterns[54767] = 25'b11010101_11101101_11000010_1;
      patterns[54768] = 25'b11010101_11101110_11000011_1;
      patterns[54769] = 25'b11010101_11101111_11000100_1;
      patterns[54770] = 25'b11010101_11110000_11000101_1;
      patterns[54771] = 25'b11010101_11110001_11000110_1;
      patterns[54772] = 25'b11010101_11110010_11000111_1;
      patterns[54773] = 25'b11010101_11110011_11001000_1;
      patterns[54774] = 25'b11010101_11110100_11001001_1;
      patterns[54775] = 25'b11010101_11110101_11001010_1;
      patterns[54776] = 25'b11010101_11110110_11001011_1;
      patterns[54777] = 25'b11010101_11110111_11001100_1;
      patterns[54778] = 25'b11010101_11111000_11001101_1;
      patterns[54779] = 25'b11010101_11111001_11001110_1;
      patterns[54780] = 25'b11010101_11111010_11001111_1;
      patterns[54781] = 25'b11010101_11111011_11010000_1;
      patterns[54782] = 25'b11010101_11111100_11010001_1;
      patterns[54783] = 25'b11010101_11111101_11010010_1;
      patterns[54784] = 25'b11010101_11111110_11010011_1;
      patterns[54785] = 25'b11010101_11111111_11010100_1;
      patterns[54786] = 25'b11010110_00000000_11010110_0;
      patterns[54787] = 25'b11010110_00000001_11010111_0;
      patterns[54788] = 25'b11010110_00000010_11011000_0;
      patterns[54789] = 25'b11010110_00000011_11011001_0;
      patterns[54790] = 25'b11010110_00000100_11011010_0;
      patterns[54791] = 25'b11010110_00000101_11011011_0;
      patterns[54792] = 25'b11010110_00000110_11011100_0;
      patterns[54793] = 25'b11010110_00000111_11011101_0;
      patterns[54794] = 25'b11010110_00001000_11011110_0;
      patterns[54795] = 25'b11010110_00001001_11011111_0;
      patterns[54796] = 25'b11010110_00001010_11100000_0;
      patterns[54797] = 25'b11010110_00001011_11100001_0;
      patterns[54798] = 25'b11010110_00001100_11100010_0;
      patterns[54799] = 25'b11010110_00001101_11100011_0;
      patterns[54800] = 25'b11010110_00001110_11100100_0;
      patterns[54801] = 25'b11010110_00001111_11100101_0;
      patterns[54802] = 25'b11010110_00010000_11100110_0;
      patterns[54803] = 25'b11010110_00010001_11100111_0;
      patterns[54804] = 25'b11010110_00010010_11101000_0;
      patterns[54805] = 25'b11010110_00010011_11101001_0;
      patterns[54806] = 25'b11010110_00010100_11101010_0;
      patterns[54807] = 25'b11010110_00010101_11101011_0;
      patterns[54808] = 25'b11010110_00010110_11101100_0;
      patterns[54809] = 25'b11010110_00010111_11101101_0;
      patterns[54810] = 25'b11010110_00011000_11101110_0;
      patterns[54811] = 25'b11010110_00011001_11101111_0;
      patterns[54812] = 25'b11010110_00011010_11110000_0;
      patterns[54813] = 25'b11010110_00011011_11110001_0;
      patterns[54814] = 25'b11010110_00011100_11110010_0;
      patterns[54815] = 25'b11010110_00011101_11110011_0;
      patterns[54816] = 25'b11010110_00011110_11110100_0;
      patterns[54817] = 25'b11010110_00011111_11110101_0;
      patterns[54818] = 25'b11010110_00100000_11110110_0;
      patterns[54819] = 25'b11010110_00100001_11110111_0;
      patterns[54820] = 25'b11010110_00100010_11111000_0;
      patterns[54821] = 25'b11010110_00100011_11111001_0;
      patterns[54822] = 25'b11010110_00100100_11111010_0;
      patterns[54823] = 25'b11010110_00100101_11111011_0;
      patterns[54824] = 25'b11010110_00100110_11111100_0;
      patterns[54825] = 25'b11010110_00100111_11111101_0;
      patterns[54826] = 25'b11010110_00101000_11111110_0;
      patterns[54827] = 25'b11010110_00101001_11111111_0;
      patterns[54828] = 25'b11010110_00101010_00000000_1;
      patterns[54829] = 25'b11010110_00101011_00000001_1;
      patterns[54830] = 25'b11010110_00101100_00000010_1;
      patterns[54831] = 25'b11010110_00101101_00000011_1;
      patterns[54832] = 25'b11010110_00101110_00000100_1;
      patterns[54833] = 25'b11010110_00101111_00000101_1;
      patterns[54834] = 25'b11010110_00110000_00000110_1;
      patterns[54835] = 25'b11010110_00110001_00000111_1;
      patterns[54836] = 25'b11010110_00110010_00001000_1;
      patterns[54837] = 25'b11010110_00110011_00001001_1;
      patterns[54838] = 25'b11010110_00110100_00001010_1;
      patterns[54839] = 25'b11010110_00110101_00001011_1;
      patterns[54840] = 25'b11010110_00110110_00001100_1;
      patterns[54841] = 25'b11010110_00110111_00001101_1;
      patterns[54842] = 25'b11010110_00111000_00001110_1;
      patterns[54843] = 25'b11010110_00111001_00001111_1;
      patterns[54844] = 25'b11010110_00111010_00010000_1;
      patterns[54845] = 25'b11010110_00111011_00010001_1;
      patterns[54846] = 25'b11010110_00111100_00010010_1;
      patterns[54847] = 25'b11010110_00111101_00010011_1;
      patterns[54848] = 25'b11010110_00111110_00010100_1;
      patterns[54849] = 25'b11010110_00111111_00010101_1;
      patterns[54850] = 25'b11010110_01000000_00010110_1;
      patterns[54851] = 25'b11010110_01000001_00010111_1;
      patterns[54852] = 25'b11010110_01000010_00011000_1;
      patterns[54853] = 25'b11010110_01000011_00011001_1;
      patterns[54854] = 25'b11010110_01000100_00011010_1;
      patterns[54855] = 25'b11010110_01000101_00011011_1;
      patterns[54856] = 25'b11010110_01000110_00011100_1;
      patterns[54857] = 25'b11010110_01000111_00011101_1;
      patterns[54858] = 25'b11010110_01001000_00011110_1;
      patterns[54859] = 25'b11010110_01001001_00011111_1;
      patterns[54860] = 25'b11010110_01001010_00100000_1;
      patterns[54861] = 25'b11010110_01001011_00100001_1;
      patterns[54862] = 25'b11010110_01001100_00100010_1;
      patterns[54863] = 25'b11010110_01001101_00100011_1;
      patterns[54864] = 25'b11010110_01001110_00100100_1;
      patterns[54865] = 25'b11010110_01001111_00100101_1;
      patterns[54866] = 25'b11010110_01010000_00100110_1;
      patterns[54867] = 25'b11010110_01010001_00100111_1;
      patterns[54868] = 25'b11010110_01010010_00101000_1;
      patterns[54869] = 25'b11010110_01010011_00101001_1;
      patterns[54870] = 25'b11010110_01010100_00101010_1;
      patterns[54871] = 25'b11010110_01010101_00101011_1;
      patterns[54872] = 25'b11010110_01010110_00101100_1;
      patterns[54873] = 25'b11010110_01010111_00101101_1;
      patterns[54874] = 25'b11010110_01011000_00101110_1;
      patterns[54875] = 25'b11010110_01011001_00101111_1;
      patterns[54876] = 25'b11010110_01011010_00110000_1;
      patterns[54877] = 25'b11010110_01011011_00110001_1;
      patterns[54878] = 25'b11010110_01011100_00110010_1;
      patterns[54879] = 25'b11010110_01011101_00110011_1;
      patterns[54880] = 25'b11010110_01011110_00110100_1;
      patterns[54881] = 25'b11010110_01011111_00110101_1;
      patterns[54882] = 25'b11010110_01100000_00110110_1;
      patterns[54883] = 25'b11010110_01100001_00110111_1;
      patterns[54884] = 25'b11010110_01100010_00111000_1;
      patterns[54885] = 25'b11010110_01100011_00111001_1;
      patterns[54886] = 25'b11010110_01100100_00111010_1;
      patterns[54887] = 25'b11010110_01100101_00111011_1;
      patterns[54888] = 25'b11010110_01100110_00111100_1;
      patterns[54889] = 25'b11010110_01100111_00111101_1;
      patterns[54890] = 25'b11010110_01101000_00111110_1;
      patterns[54891] = 25'b11010110_01101001_00111111_1;
      patterns[54892] = 25'b11010110_01101010_01000000_1;
      patterns[54893] = 25'b11010110_01101011_01000001_1;
      patterns[54894] = 25'b11010110_01101100_01000010_1;
      patterns[54895] = 25'b11010110_01101101_01000011_1;
      patterns[54896] = 25'b11010110_01101110_01000100_1;
      patterns[54897] = 25'b11010110_01101111_01000101_1;
      patterns[54898] = 25'b11010110_01110000_01000110_1;
      patterns[54899] = 25'b11010110_01110001_01000111_1;
      patterns[54900] = 25'b11010110_01110010_01001000_1;
      patterns[54901] = 25'b11010110_01110011_01001001_1;
      patterns[54902] = 25'b11010110_01110100_01001010_1;
      patterns[54903] = 25'b11010110_01110101_01001011_1;
      patterns[54904] = 25'b11010110_01110110_01001100_1;
      patterns[54905] = 25'b11010110_01110111_01001101_1;
      patterns[54906] = 25'b11010110_01111000_01001110_1;
      patterns[54907] = 25'b11010110_01111001_01001111_1;
      patterns[54908] = 25'b11010110_01111010_01010000_1;
      patterns[54909] = 25'b11010110_01111011_01010001_1;
      patterns[54910] = 25'b11010110_01111100_01010010_1;
      patterns[54911] = 25'b11010110_01111101_01010011_1;
      patterns[54912] = 25'b11010110_01111110_01010100_1;
      patterns[54913] = 25'b11010110_01111111_01010101_1;
      patterns[54914] = 25'b11010110_10000000_01010110_1;
      patterns[54915] = 25'b11010110_10000001_01010111_1;
      patterns[54916] = 25'b11010110_10000010_01011000_1;
      patterns[54917] = 25'b11010110_10000011_01011001_1;
      patterns[54918] = 25'b11010110_10000100_01011010_1;
      patterns[54919] = 25'b11010110_10000101_01011011_1;
      patterns[54920] = 25'b11010110_10000110_01011100_1;
      patterns[54921] = 25'b11010110_10000111_01011101_1;
      patterns[54922] = 25'b11010110_10001000_01011110_1;
      patterns[54923] = 25'b11010110_10001001_01011111_1;
      patterns[54924] = 25'b11010110_10001010_01100000_1;
      patterns[54925] = 25'b11010110_10001011_01100001_1;
      patterns[54926] = 25'b11010110_10001100_01100010_1;
      patterns[54927] = 25'b11010110_10001101_01100011_1;
      patterns[54928] = 25'b11010110_10001110_01100100_1;
      patterns[54929] = 25'b11010110_10001111_01100101_1;
      patterns[54930] = 25'b11010110_10010000_01100110_1;
      patterns[54931] = 25'b11010110_10010001_01100111_1;
      patterns[54932] = 25'b11010110_10010010_01101000_1;
      patterns[54933] = 25'b11010110_10010011_01101001_1;
      patterns[54934] = 25'b11010110_10010100_01101010_1;
      patterns[54935] = 25'b11010110_10010101_01101011_1;
      patterns[54936] = 25'b11010110_10010110_01101100_1;
      patterns[54937] = 25'b11010110_10010111_01101101_1;
      patterns[54938] = 25'b11010110_10011000_01101110_1;
      patterns[54939] = 25'b11010110_10011001_01101111_1;
      patterns[54940] = 25'b11010110_10011010_01110000_1;
      patterns[54941] = 25'b11010110_10011011_01110001_1;
      patterns[54942] = 25'b11010110_10011100_01110010_1;
      patterns[54943] = 25'b11010110_10011101_01110011_1;
      patterns[54944] = 25'b11010110_10011110_01110100_1;
      patterns[54945] = 25'b11010110_10011111_01110101_1;
      patterns[54946] = 25'b11010110_10100000_01110110_1;
      patterns[54947] = 25'b11010110_10100001_01110111_1;
      patterns[54948] = 25'b11010110_10100010_01111000_1;
      patterns[54949] = 25'b11010110_10100011_01111001_1;
      patterns[54950] = 25'b11010110_10100100_01111010_1;
      patterns[54951] = 25'b11010110_10100101_01111011_1;
      patterns[54952] = 25'b11010110_10100110_01111100_1;
      patterns[54953] = 25'b11010110_10100111_01111101_1;
      patterns[54954] = 25'b11010110_10101000_01111110_1;
      patterns[54955] = 25'b11010110_10101001_01111111_1;
      patterns[54956] = 25'b11010110_10101010_10000000_1;
      patterns[54957] = 25'b11010110_10101011_10000001_1;
      patterns[54958] = 25'b11010110_10101100_10000010_1;
      patterns[54959] = 25'b11010110_10101101_10000011_1;
      patterns[54960] = 25'b11010110_10101110_10000100_1;
      patterns[54961] = 25'b11010110_10101111_10000101_1;
      patterns[54962] = 25'b11010110_10110000_10000110_1;
      patterns[54963] = 25'b11010110_10110001_10000111_1;
      patterns[54964] = 25'b11010110_10110010_10001000_1;
      patterns[54965] = 25'b11010110_10110011_10001001_1;
      patterns[54966] = 25'b11010110_10110100_10001010_1;
      patterns[54967] = 25'b11010110_10110101_10001011_1;
      patterns[54968] = 25'b11010110_10110110_10001100_1;
      patterns[54969] = 25'b11010110_10110111_10001101_1;
      patterns[54970] = 25'b11010110_10111000_10001110_1;
      patterns[54971] = 25'b11010110_10111001_10001111_1;
      patterns[54972] = 25'b11010110_10111010_10010000_1;
      patterns[54973] = 25'b11010110_10111011_10010001_1;
      patterns[54974] = 25'b11010110_10111100_10010010_1;
      patterns[54975] = 25'b11010110_10111101_10010011_1;
      patterns[54976] = 25'b11010110_10111110_10010100_1;
      patterns[54977] = 25'b11010110_10111111_10010101_1;
      patterns[54978] = 25'b11010110_11000000_10010110_1;
      patterns[54979] = 25'b11010110_11000001_10010111_1;
      patterns[54980] = 25'b11010110_11000010_10011000_1;
      patterns[54981] = 25'b11010110_11000011_10011001_1;
      patterns[54982] = 25'b11010110_11000100_10011010_1;
      patterns[54983] = 25'b11010110_11000101_10011011_1;
      patterns[54984] = 25'b11010110_11000110_10011100_1;
      patterns[54985] = 25'b11010110_11000111_10011101_1;
      patterns[54986] = 25'b11010110_11001000_10011110_1;
      patterns[54987] = 25'b11010110_11001001_10011111_1;
      patterns[54988] = 25'b11010110_11001010_10100000_1;
      patterns[54989] = 25'b11010110_11001011_10100001_1;
      patterns[54990] = 25'b11010110_11001100_10100010_1;
      patterns[54991] = 25'b11010110_11001101_10100011_1;
      patterns[54992] = 25'b11010110_11001110_10100100_1;
      patterns[54993] = 25'b11010110_11001111_10100101_1;
      patterns[54994] = 25'b11010110_11010000_10100110_1;
      patterns[54995] = 25'b11010110_11010001_10100111_1;
      patterns[54996] = 25'b11010110_11010010_10101000_1;
      patterns[54997] = 25'b11010110_11010011_10101001_1;
      patterns[54998] = 25'b11010110_11010100_10101010_1;
      patterns[54999] = 25'b11010110_11010101_10101011_1;
      patterns[55000] = 25'b11010110_11010110_10101100_1;
      patterns[55001] = 25'b11010110_11010111_10101101_1;
      patterns[55002] = 25'b11010110_11011000_10101110_1;
      patterns[55003] = 25'b11010110_11011001_10101111_1;
      patterns[55004] = 25'b11010110_11011010_10110000_1;
      patterns[55005] = 25'b11010110_11011011_10110001_1;
      patterns[55006] = 25'b11010110_11011100_10110010_1;
      patterns[55007] = 25'b11010110_11011101_10110011_1;
      patterns[55008] = 25'b11010110_11011110_10110100_1;
      patterns[55009] = 25'b11010110_11011111_10110101_1;
      patterns[55010] = 25'b11010110_11100000_10110110_1;
      patterns[55011] = 25'b11010110_11100001_10110111_1;
      patterns[55012] = 25'b11010110_11100010_10111000_1;
      patterns[55013] = 25'b11010110_11100011_10111001_1;
      patterns[55014] = 25'b11010110_11100100_10111010_1;
      patterns[55015] = 25'b11010110_11100101_10111011_1;
      patterns[55016] = 25'b11010110_11100110_10111100_1;
      patterns[55017] = 25'b11010110_11100111_10111101_1;
      patterns[55018] = 25'b11010110_11101000_10111110_1;
      patterns[55019] = 25'b11010110_11101001_10111111_1;
      patterns[55020] = 25'b11010110_11101010_11000000_1;
      patterns[55021] = 25'b11010110_11101011_11000001_1;
      patterns[55022] = 25'b11010110_11101100_11000010_1;
      patterns[55023] = 25'b11010110_11101101_11000011_1;
      patterns[55024] = 25'b11010110_11101110_11000100_1;
      patterns[55025] = 25'b11010110_11101111_11000101_1;
      patterns[55026] = 25'b11010110_11110000_11000110_1;
      patterns[55027] = 25'b11010110_11110001_11000111_1;
      patterns[55028] = 25'b11010110_11110010_11001000_1;
      patterns[55029] = 25'b11010110_11110011_11001001_1;
      patterns[55030] = 25'b11010110_11110100_11001010_1;
      patterns[55031] = 25'b11010110_11110101_11001011_1;
      patterns[55032] = 25'b11010110_11110110_11001100_1;
      patterns[55033] = 25'b11010110_11110111_11001101_1;
      patterns[55034] = 25'b11010110_11111000_11001110_1;
      patterns[55035] = 25'b11010110_11111001_11001111_1;
      patterns[55036] = 25'b11010110_11111010_11010000_1;
      patterns[55037] = 25'b11010110_11111011_11010001_1;
      patterns[55038] = 25'b11010110_11111100_11010010_1;
      patterns[55039] = 25'b11010110_11111101_11010011_1;
      patterns[55040] = 25'b11010110_11111110_11010100_1;
      patterns[55041] = 25'b11010110_11111111_11010101_1;
      patterns[55042] = 25'b11010111_00000000_11010111_0;
      patterns[55043] = 25'b11010111_00000001_11011000_0;
      patterns[55044] = 25'b11010111_00000010_11011001_0;
      patterns[55045] = 25'b11010111_00000011_11011010_0;
      patterns[55046] = 25'b11010111_00000100_11011011_0;
      patterns[55047] = 25'b11010111_00000101_11011100_0;
      patterns[55048] = 25'b11010111_00000110_11011101_0;
      patterns[55049] = 25'b11010111_00000111_11011110_0;
      patterns[55050] = 25'b11010111_00001000_11011111_0;
      patterns[55051] = 25'b11010111_00001001_11100000_0;
      patterns[55052] = 25'b11010111_00001010_11100001_0;
      patterns[55053] = 25'b11010111_00001011_11100010_0;
      patterns[55054] = 25'b11010111_00001100_11100011_0;
      patterns[55055] = 25'b11010111_00001101_11100100_0;
      patterns[55056] = 25'b11010111_00001110_11100101_0;
      patterns[55057] = 25'b11010111_00001111_11100110_0;
      patterns[55058] = 25'b11010111_00010000_11100111_0;
      patterns[55059] = 25'b11010111_00010001_11101000_0;
      patterns[55060] = 25'b11010111_00010010_11101001_0;
      patterns[55061] = 25'b11010111_00010011_11101010_0;
      patterns[55062] = 25'b11010111_00010100_11101011_0;
      patterns[55063] = 25'b11010111_00010101_11101100_0;
      patterns[55064] = 25'b11010111_00010110_11101101_0;
      patterns[55065] = 25'b11010111_00010111_11101110_0;
      patterns[55066] = 25'b11010111_00011000_11101111_0;
      patterns[55067] = 25'b11010111_00011001_11110000_0;
      patterns[55068] = 25'b11010111_00011010_11110001_0;
      patterns[55069] = 25'b11010111_00011011_11110010_0;
      patterns[55070] = 25'b11010111_00011100_11110011_0;
      patterns[55071] = 25'b11010111_00011101_11110100_0;
      patterns[55072] = 25'b11010111_00011110_11110101_0;
      patterns[55073] = 25'b11010111_00011111_11110110_0;
      patterns[55074] = 25'b11010111_00100000_11110111_0;
      patterns[55075] = 25'b11010111_00100001_11111000_0;
      patterns[55076] = 25'b11010111_00100010_11111001_0;
      patterns[55077] = 25'b11010111_00100011_11111010_0;
      patterns[55078] = 25'b11010111_00100100_11111011_0;
      patterns[55079] = 25'b11010111_00100101_11111100_0;
      patterns[55080] = 25'b11010111_00100110_11111101_0;
      patterns[55081] = 25'b11010111_00100111_11111110_0;
      patterns[55082] = 25'b11010111_00101000_11111111_0;
      patterns[55083] = 25'b11010111_00101001_00000000_1;
      patterns[55084] = 25'b11010111_00101010_00000001_1;
      patterns[55085] = 25'b11010111_00101011_00000010_1;
      patterns[55086] = 25'b11010111_00101100_00000011_1;
      patterns[55087] = 25'b11010111_00101101_00000100_1;
      patterns[55088] = 25'b11010111_00101110_00000101_1;
      patterns[55089] = 25'b11010111_00101111_00000110_1;
      patterns[55090] = 25'b11010111_00110000_00000111_1;
      patterns[55091] = 25'b11010111_00110001_00001000_1;
      patterns[55092] = 25'b11010111_00110010_00001001_1;
      patterns[55093] = 25'b11010111_00110011_00001010_1;
      patterns[55094] = 25'b11010111_00110100_00001011_1;
      patterns[55095] = 25'b11010111_00110101_00001100_1;
      patterns[55096] = 25'b11010111_00110110_00001101_1;
      patterns[55097] = 25'b11010111_00110111_00001110_1;
      patterns[55098] = 25'b11010111_00111000_00001111_1;
      patterns[55099] = 25'b11010111_00111001_00010000_1;
      patterns[55100] = 25'b11010111_00111010_00010001_1;
      patterns[55101] = 25'b11010111_00111011_00010010_1;
      patterns[55102] = 25'b11010111_00111100_00010011_1;
      patterns[55103] = 25'b11010111_00111101_00010100_1;
      patterns[55104] = 25'b11010111_00111110_00010101_1;
      patterns[55105] = 25'b11010111_00111111_00010110_1;
      patterns[55106] = 25'b11010111_01000000_00010111_1;
      patterns[55107] = 25'b11010111_01000001_00011000_1;
      patterns[55108] = 25'b11010111_01000010_00011001_1;
      patterns[55109] = 25'b11010111_01000011_00011010_1;
      patterns[55110] = 25'b11010111_01000100_00011011_1;
      patterns[55111] = 25'b11010111_01000101_00011100_1;
      patterns[55112] = 25'b11010111_01000110_00011101_1;
      patterns[55113] = 25'b11010111_01000111_00011110_1;
      patterns[55114] = 25'b11010111_01001000_00011111_1;
      patterns[55115] = 25'b11010111_01001001_00100000_1;
      patterns[55116] = 25'b11010111_01001010_00100001_1;
      patterns[55117] = 25'b11010111_01001011_00100010_1;
      patterns[55118] = 25'b11010111_01001100_00100011_1;
      patterns[55119] = 25'b11010111_01001101_00100100_1;
      patterns[55120] = 25'b11010111_01001110_00100101_1;
      patterns[55121] = 25'b11010111_01001111_00100110_1;
      patterns[55122] = 25'b11010111_01010000_00100111_1;
      patterns[55123] = 25'b11010111_01010001_00101000_1;
      patterns[55124] = 25'b11010111_01010010_00101001_1;
      patterns[55125] = 25'b11010111_01010011_00101010_1;
      patterns[55126] = 25'b11010111_01010100_00101011_1;
      patterns[55127] = 25'b11010111_01010101_00101100_1;
      patterns[55128] = 25'b11010111_01010110_00101101_1;
      patterns[55129] = 25'b11010111_01010111_00101110_1;
      patterns[55130] = 25'b11010111_01011000_00101111_1;
      patterns[55131] = 25'b11010111_01011001_00110000_1;
      patterns[55132] = 25'b11010111_01011010_00110001_1;
      patterns[55133] = 25'b11010111_01011011_00110010_1;
      patterns[55134] = 25'b11010111_01011100_00110011_1;
      patterns[55135] = 25'b11010111_01011101_00110100_1;
      patterns[55136] = 25'b11010111_01011110_00110101_1;
      patterns[55137] = 25'b11010111_01011111_00110110_1;
      patterns[55138] = 25'b11010111_01100000_00110111_1;
      patterns[55139] = 25'b11010111_01100001_00111000_1;
      patterns[55140] = 25'b11010111_01100010_00111001_1;
      patterns[55141] = 25'b11010111_01100011_00111010_1;
      patterns[55142] = 25'b11010111_01100100_00111011_1;
      patterns[55143] = 25'b11010111_01100101_00111100_1;
      patterns[55144] = 25'b11010111_01100110_00111101_1;
      patterns[55145] = 25'b11010111_01100111_00111110_1;
      patterns[55146] = 25'b11010111_01101000_00111111_1;
      patterns[55147] = 25'b11010111_01101001_01000000_1;
      patterns[55148] = 25'b11010111_01101010_01000001_1;
      patterns[55149] = 25'b11010111_01101011_01000010_1;
      patterns[55150] = 25'b11010111_01101100_01000011_1;
      patterns[55151] = 25'b11010111_01101101_01000100_1;
      patterns[55152] = 25'b11010111_01101110_01000101_1;
      patterns[55153] = 25'b11010111_01101111_01000110_1;
      patterns[55154] = 25'b11010111_01110000_01000111_1;
      patterns[55155] = 25'b11010111_01110001_01001000_1;
      patterns[55156] = 25'b11010111_01110010_01001001_1;
      patterns[55157] = 25'b11010111_01110011_01001010_1;
      patterns[55158] = 25'b11010111_01110100_01001011_1;
      patterns[55159] = 25'b11010111_01110101_01001100_1;
      patterns[55160] = 25'b11010111_01110110_01001101_1;
      patterns[55161] = 25'b11010111_01110111_01001110_1;
      patterns[55162] = 25'b11010111_01111000_01001111_1;
      patterns[55163] = 25'b11010111_01111001_01010000_1;
      patterns[55164] = 25'b11010111_01111010_01010001_1;
      patterns[55165] = 25'b11010111_01111011_01010010_1;
      patterns[55166] = 25'b11010111_01111100_01010011_1;
      patterns[55167] = 25'b11010111_01111101_01010100_1;
      patterns[55168] = 25'b11010111_01111110_01010101_1;
      patterns[55169] = 25'b11010111_01111111_01010110_1;
      patterns[55170] = 25'b11010111_10000000_01010111_1;
      patterns[55171] = 25'b11010111_10000001_01011000_1;
      patterns[55172] = 25'b11010111_10000010_01011001_1;
      patterns[55173] = 25'b11010111_10000011_01011010_1;
      patterns[55174] = 25'b11010111_10000100_01011011_1;
      patterns[55175] = 25'b11010111_10000101_01011100_1;
      patterns[55176] = 25'b11010111_10000110_01011101_1;
      patterns[55177] = 25'b11010111_10000111_01011110_1;
      patterns[55178] = 25'b11010111_10001000_01011111_1;
      patterns[55179] = 25'b11010111_10001001_01100000_1;
      patterns[55180] = 25'b11010111_10001010_01100001_1;
      patterns[55181] = 25'b11010111_10001011_01100010_1;
      patterns[55182] = 25'b11010111_10001100_01100011_1;
      patterns[55183] = 25'b11010111_10001101_01100100_1;
      patterns[55184] = 25'b11010111_10001110_01100101_1;
      patterns[55185] = 25'b11010111_10001111_01100110_1;
      patterns[55186] = 25'b11010111_10010000_01100111_1;
      patterns[55187] = 25'b11010111_10010001_01101000_1;
      patterns[55188] = 25'b11010111_10010010_01101001_1;
      patterns[55189] = 25'b11010111_10010011_01101010_1;
      patterns[55190] = 25'b11010111_10010100_01101011_1;
      patterns[55191] = 25'b11010111_10010101_01101100_1;
      patterns[55192] = 25'b11010111_10010110_01101101_1;
      patterns[55193] = 25'b11010111_10010111_01101110_1;
      patterns[55194] = 25'b11010111_10011000_01101111_1;
      patterns[55195] = 25'b11010111_10011001_01110000_1;
      patterns[55196] = 25'b11010111_10011010_01110001_1;
      patterns[55197] = 25'b11010111_10011011_01110010_1;
      patterns[55198] = 25'b11010111_10011100_01110011_1;
      patterns[55199] = 25'b11010111_10011101_01110100_1;
      patterns[55200] = 25'b11010111_10011110_01110101_1;
      patterns[55201] = 25'b11010111_10011111_01110110_1;
      patterns[55202] = 25'b11010111_10100000_01110111_1;
      patterns[55203] = 25'b11010111_10100001_01111000_1;
      patterns[55204] = 25'b11010111_10100010_01111001_1;
      patterns[55205] = 25'b11010111_10100011_01111010_1;
      patterns[55206] = 25'b11010111_10100100_01111011_1;
      patterns[55207] = 25'b11010111_10100101_01111100_1;
      patterns[55208] = 25'b11010111_10100110_01111101_1;
      patterns[55209] = 25'b11010111_10100111_01111110_1;
      patterns[55210] = 25'b11010111_10101000_01111111_1;
      patterns[55211] = 25'b11010111_10101001_10000000_1;
      patterns[55212] = 25'b11010111_10101010_10000001_1;
      patterns[55213] = 25'b11010111_10101011_10000010_1;
      patterns[55214] = 25'b11010111_10101100_10000011_1;
      patterns[55215] = 25'b11010111_10101101_10000100_1;
      patterns[55216] = 25'b11010111_10101110_10000101_1;
      patterns[55217] = 25'b11010111_10101111_10000110_1;
      patterns[55218] = 25'b11010111_10110000_10000111_1;
      patterns[55219] = 25'b11010111_10110001_10001000_1;
      patterns[55220] = 25'b11010111_10110010_10001001_1;
      patterns[55221] = 25'b11010111_10110011_10001010_1;
      patterns[55222] = 25'b11010111_10110100_10001011_1;
      patterns[55223] = 25'b11010111_10110101_10001100_1;
      patterns[55224] = 25'b11010111_10110110_10001101_1;
      patterns[55225] = 25'b11010111_10110111_10001110_1;
      patterns[55226] = 25'b11010111_10111000_10001111_1;
      patterns[55227] = 25'b11010111_10111001_10010000_1;
      patterns[55228] = 25'b11010111_10111010_10010001_1;
      patterns[55229] = 25'b11010111_10111011_10010010_1;
      patterns[55230] = 25'b11010111_10111100_10010011_1;
      patterns[55231] = 25'b11010111_10111101_10010100_1;
      patterns[55232] = 25'b11010111_10111110_10010101_1;
      patterns[55233] = 25'b11010111_10111111_10010110_1;
      patterns[55234] = 25'b11010111_11000000_10010111_1;
      patterns[55235] = 25'b11010111_11000001_10011000_1;
      patterns[55236] = 25'b11010111_11000010_10011001_1;
      patterns[55237] = 25'b11010111_11000011_10011010_1;
      patterns[55238] = 25'b11010111_11000100_10011011_1;
      patterns[55239] = 25'b11010111_11000101_10011100_1;
      patterns[55240] = 25'b11010111_11000110_10011101_1;
      patterns[55241] = 25'b11010111_11000111_10011110_1;
      patterns[55242] = 25'b11010111_11001000_10011111_1;
      patterns[55243] = 25'b11010111_11001001_10100000_1;
      patterns[55244] = 25'b11010111_11001010_10100001_1;
      patterns[55245] = 25'b11010111_11001011_10100010_1;
      patterns[55246] = 25'b11010111_11001100_10100011_1;
      patterns[55247] = 25'b11010111_11001101_10100100_1;
      patterns[55248] = 25'b11010111_11001110_10100101_1;
      patterns[55249] = 25'b11010111_11001111_10100110_1;
      patterns[55250] = 25'b11010111_11010000_10100111_1;
      patterns[55251] = 25'b11010111_11010001_10101000_1;
      patterns[55252] = 25'b11010111_11010010_10101001_1;
      patterns[55253] = 25'b11010111_11010011_10101010_1;
      patterns[55254] = 25'b11010111_11010100_10101011_1;
      patterns[55255] = 25'b11010111_11010101_10101100_1;
      patterns[55256] = 25'b11010111_11010110_10101101_1;
      patterns[55257] = 25'b11010111_11010111_10101110_1;
      patterns[55258] = 25'b11010111_11011000_10101111_1;
      patterns[55259] = 25'b11010111_11011001_10110000_1;
      patterns[55260] = 25'b11010111_11011010_10110001_1;
      patterns[55261] = 25'b11010111_11011011_10110010_1;
      patterns[55262] = 25'b11010111_11011100_10110011_1;
      patterns[55263] = 25'b11010111_11011101_10110100_1;
      patterns[55264] = 25'b11010111_11011110_10110101_1;
      patterns[55265] = 25'b11010111_11011111_10110110_1;
      patterns[55266] = 25'b11010111_11100000_10110111_1;
      patterns[55267] = 25'b11010111_11100001_10111000_1;
      patterns[55268] = 25'b11010111_11100010_10111001_1;
      patterns[55269] = 25'b11010111_11100011_10111010_1;
      patterns[55270] = 25'b11010111_11100100_10111011_1;
      patterns[55271] = 25'b11010111_11100101_10111100_1;
      patterns[55272] = 25'b11010111_11100110_10111101_1;
      patterns[55273] = 25'b11010111_11100111_10111110_1;
      patterns[55274] = 25'b11010111_11101000_10111111_1;
      patterns[55275] = 25'b11010111_11101001_11000000_1;
      patterns[55276] = 25'b11010111_11101010_11000001_1;
      patterns[55277] = 25'b11010111_11101011_11000010_1;
      patterns[55278] = 25'b11010111_11101100_11000011_1;
      patterns[55279] = 25'b11010111_11101101_11000100_1;
      patterns[55280] = 25'b11010111_11101110_11000101_1;
      patterns[55281] = 25'b11010111_11101111_11000110_1;
      patterns[55282] = 25'b11010111_11110000_11000111_1;
      patterns[55283] = 25'b11010111_11110001_11001000_1;
      patterns[55284] = 25'b11010111_11110010_11001001_1;
      patterns[55285] = 25'b11010111_11110011_11001010_1;
      patterns[55286] = 25'b11010111_11110100_11001011_1;
      patterns[55287] = 25'b11010111_11110101_11001100_1;
      patterns[55288] = 25'b11010111_11110110_11001101_1;
      patterns[55289] = 25'b11010111_11110111_11001110_1;
      patterns[55290] = 25'b11010111_11111000_11001111_1;
      patterns[55291] = 25'b11010111_11111001_11010000_1;
      patterns[55292] = 25'b11010111_11111010_11010001_1;
      patterns[55293] = 25'b11010111_11111011_11010010_1;
      patterns[55294] = 25'b11010111_11111100_11010011_1;
      patterns[55295] = 25'b11010111_11111101_11010100_1;
      patterns[55296] = 25'b11010111_11111110_11010101_1;
      patterns[55297] = 25'b11010111_11111111_11010110_1;
      patterns[55298] = 25'b11011000_00000000_11011000_0;
      patterns[55299] = 25'b11011000_00000001_11011001_0;
      patterns[55300] = 25'b11011000_00000010_11011010_0;
      patterns[55301] = 25'b11011000_00000011_11011011_0;
      patterns[55302] = 25'b11011000_00000100_11011100_0;
      patterns[55303] = 25'b11011000_00000101_11011101_0;
      patterns[55304] = 25'b11011000_00000110_11011110_0;
      patterns[55305] = 25'b11011000_00000111_11011111_0;
      patterns[55306] = 25'b11011000_00001000_11100000_0;
      patterns[55307] = 25'b11011000_00001001_11100001_0;
      patterns[55308] = 25'b11011000_00001010_11100010_0;
      patterns[55309] = 25'b11011000_00001011_11100011_0;
      patterns[55310] = 25'b11011000_00001100_11100100_0;
      patterns[55311] = 25'b11011000_00001101_11100101_0;
      patterns[55312] = 25'b11011000_00001110_11100110_0;
      patterns[55313] = 25'b11011000_00001111_11100111_0;
      patterns[55314] = 25'b11011000_00010000_11101000_0;
      patterns[55315] = 25'b11011000_00010001_11101001_0;
      patterns[55316] = 25'b11011000_00010010_11101010_0;
      patterns[55317] = 25'b11011000_00010011_11101011_0;
      patterns[55318] = 25'b11011000_00010100_11101100_0;
      patterns[55319] = 25'b11011000_00010101_11101101_0;
      patterns[55320] = 25'b11011000_00010110_11101110_0;
      patterns[55321] = 25'b11011000_00010111_11101111_0;
      patterns[55322] = 25'b11011000_00011000_11110000_0;
      patterns[55323] = 25'b11011000_00011001_11110001_0;
      patterns[55324] = 25'b11011000_00011010_11110010_0;
      patterns[55325] = 25'b11011000_00011011_11110011_0;
      patterns[55326] = 25'b11011000_00011100_11110100_0;
      patterns[55327] = 25'b11011000_00011101_11110101_0;
      patterns[55328] = 25'b11011000_00011110_11110110_0;
      patterns[55329] = 25'b11011000_00011111_11110111_0;
      patterns[55330] = 25'b11011000_00100000_11111000_0;
      patterns[55331] = 25'b11011000_00100001_11111001_0;
      patterns[55332] = 25'b11011000_00100010_11111010_0;
      patterns[55333] = 25'b11011000_00100011_11111011_0;
      patterns[55334] = 25'b11011000_00100100_11111100_0;
      patterns[55335] = 25'b11011000_00100101_11111101_0;
      patterns[55336] = 25'b11011000_00100110_11111110_0;
      patterns[55337] = 25'b11011000_00100111_11111111_0;
      patterns[55338] = 25'b11011000_00101000_00000000_1;
      patterns[55339] = 25'b11011000_00101001_00000001_1;
      patterns[55340] = 25'b11011000_00101010_00000010_1;
      patterns[55341] = 25'b11011000_00101011_00000011_1;
      patterns[55342] = 25'b11011000_00101100_00000100_1;
      patterns[55343] = 25'b11011000_00101101_00000101_1;
      patterns[55344] = 25'b11011000_00101110_00000110_1;
      patterns[55345] = 25'b11011000_00101111_00000111_1;
      patterns[55346] = 25'b11011000_00110000_00001000_1;
      patterns[55347] = 25'b11011000_00110001_00001001_1;
      patterns[55348] = 25'b11011000_00110010_00001010_1;
      patterns[55349] = 25'b11011000_00110011_00001011_1;
      patterns[55350] = 25'b11011000_00110100_00001100_1;
      patterns[55351] = 25'b11011000_00110101_00001101_1;
      patterns[55352] = 25'b11011000_00110110_00001110_1;
      patterns[55353] = 25'b11011000_00110111_00001111_1;
      patterns[55354] = 25'b11011000_00111000_00010000_1;
      patterns[55355] = 25'b11011000_00111001_00010001_1;
      patterns[55356] = 25'b11011000_00111010_00010010_1;
      patterns[55357] = 25'b11011000_00111011_00010011_1;
      patterns[55358] = 25'b11011000_00111100_00010100_1;
      patterns[55359] = 25'b11011000_00111101_00010101_1;
      patterns[55360] = 25'b11011000_00111110_00010110_1;
      patterns[55361] = 25'b11011000_00111111_00010111_1;
      patterns[55362] = 25'b11011000_01000000_00011000_1;
      patterns[55363] = 25'b11011000_01000001_00011001_1;
      patterns[55364] = 25'b11011000_01000010_00011010_1;
      patterns[55365] = 25'b11011000_01000011_00011011_1;
      patterns[55366] = 25'b11011000_01000100_00011100_1;
      patterns[55367] = 25'b11011000_01000101_00011101_1;
      patterns[55368] = 25'b11011000_01000110_00011110_1;
      patterns[55369] = 25'b11011000_01000111_00011111_1;
      patterns[55370] = 25'b11011000_01001000_00100000_1;
      patterns[55371] = 25'b11011000_01001001_00100001_1;
      patterns[55372] = 25'b11011000_01001010_00100010_1;
      patterns[55373] = 25'b11011000_01001011_00100011_1;
      patterns[55374] = 25'b11011000_01001100_00100100_1;
      patterns[55375] = 25'b11011000_01001101_00100101_1;
      patterns[55376] = 25'b11011000_01001110_00100110_1;
      patterns[55377] = 25'b11011000_01001111_00100111_1;
      patterns[55378] = 25'b11011000_01010000_00101000_1;
      patterns[55379] = 25'b11011000_01010001_00101001_1;
      patterns[55380] = 25'b11011000_01010010_00101010_1;
      patterns[55381] = 25'b11011000_01010011_00101011_1;
      patterns[55382] = 25'b11011000_01010100_00101100_1;
      patterns[55383] = 25'b11011000_01010101_00101101_1;
      patterns[55384] = 25'b11011000_01010110_00101110_1;
      patterns[55385] = 25'b11011000_01010111_00101111_1;
      patterns[55386] = 25'b11011000_01011000_00110000_1;
      patterns[55387] = 25'b11011000_01011001_00110001_1;
      patterns[55388] = 25'b11011000_01011010_00110010_1;
      patterns[55389] = 25'b11011000_01011011_00110011_1;
      patterns[55390] = 25'b11011000_01011100_00110100_1;
      patterns[55391] = 25'b11011000_01011101_00110101_1;
      patterns[55392] = 25'b11011000_01011110_00110110_1;
      patterns[55393] = 25'b11011000_01011111_00110111_1;
      patterns[55394] = 25'b11011000_01100000_00111000_1;
      patterns[55395] = 25'b11011000_01100001_00111001_1;
      patterns[55396] = 25'b11011000_01100010_00111010_1;
      patterns[55397] = 25'b11011000_01100011_00111011_1;
      patterns[55398] = 25'b11011000_01100100_00111100_1;
      patterns[55399] = 25'b11011000_01100101_00111101_1;
      patterns[55400] = 25'b11011000_01100110_00111110_1;
      patterns[55401] = 25'b11011000_01100111_00111111_1;
      patterns[55402] = 25'b11011000_01101000_01000000_1;
      patterns[55403] = 25'b11011000_01101001_01000001_1;
      patterns[55404] = 25'b11011000_01101010_01000010_1;
      patterns[55405] = 25'b11011000_01101011_01000011_1;
      patterns[55406] = 25'b11011000_01101100_01000100_1;
      patterns[55407] = 25'b11011000_01101101_01000101_1;
      patterns[55408] = 25'b11011000_01101110_01000110_1;
      patterns[55409] = 25'b11011000_01101111_01000111_1;
      patterns[55410] = 25'b11011000_01110000_01001000_1;
      patterns[55411] = 25'b11011000_01110001_01001001_1;
      patterns[55412] = 25'b11011000_01110010_01001010_1;
      patterns[55413] = 25'b11011000_01110011_01001011_1;
      patterns[55414] = 25'b11011000_01110100_01001100_1;
      patterns[55415] = 25'b11011000_01110101_01001101_1;
      patterns[55416] = 25'b11011000_01110110_01001110_1;
      patterns[55417] = 25'b11011000_01110111_01001111_1;
      patterns[55418] = 25'b11011000_01111000_01010000_1;
      patterns[55419] = 25'b11011000_01111001_01010001_1;
      patterns[55420] = 25'b11011000_01111010_01010010_1;
      patterns[55421] = 25'b11011000_01111011_01010011_1;
      patterns[55422] = 25'b11011000_01111100_01010100_1;
      patterns[55423] = 25'b11011000_01111101_01010101_1;
      patterns[55424] = 25'b11011000_01111110_01010110_1;
      patterns[55425] = 25'b11011000_01111111_01010111_1;
      patterns[55426] = 25'b11011000_10000000_01011000_1;
      patterns[55427] = 25'b11011000_10000001_01011001_1;
      patterns[55428] = 25'b11011000_10000010_01011010_1;
      patterns[55429] = 25'b11011000_10000011_01011011_1;
      patterns[55430] = 25'b11011000_10000100_01011100_1;
      patterns[55431] = 25'b11011000_10000101_01011101_1;
      patterns[55432] = 25'b11011000_10000110_01011110_1;
      patterns[55433] = 25'b11011000_10000111_01011111_1;
      patterns[55434] = 25'b11011000_10001000_01100000_1;
      patterns[55435] = 25'b11011000_10001001_01100001_1;
      patterns[55436] = 25'b11011000_10001010_01100010_1;
      patterns[55437] = 25'b11011000_10001011_01100011_1;
      patterns[55438] = 25'b11011000_10001100_01100100_1;
      patterns[55439] = 25'b11011000_10001101_01100101_1;
      patterns[55440] = 25'b11011000_10001110_01100110_1;
      patterns[55441] = 25'b11011000_10001111_01100111_1;
      patterns[55442] = 25'b11011000_10010000_01101000_1;
      patterns[55443] = 25'b11011000_10010001_01101001_1;
      patterns[55444] = 25'b11011000_10010010_01101010_1;
      patterns[55445] = 25'b11011000_10010011_01101011_1;
      patterns[55446] = 25'b11011000_10010100_01101100_1;
      patterns[55447] = 25'b11011000_10010101_01101101_1;
      patterns[55448] = 25'b11011000_10010110_01101110_1;
      patterns[55449] = 25'b11011000_10010111_01101111_1;
      patterns[55450] = 25'b11011000_10011000_01110000_1;
      patterns[55451] = 25'b11011000_10011001_01110001_1;
      patterns[55452] = 25'b11011000_10011010_01110010_1;
      patterns[55453] = 25'b11011000_10011011_01110011_1;
      patterns[55454] = 25'b11011000_10011100_01110100_1;
      patterns[55455] = 25'b11011000_10011101_01110101_1;
      patterns[55456] = 25'b11011000_10011110_01110110_1;
      patterns[55457] = 25'b11011000_10011111_01110111_1;
      patterns[55458] = 25'b11011000_10100000_01111000_1;
      patterns[55459] = 25'b11011000_10100001_01111001_1;
      patterns[55460] = 25'b11011000_10100010_01111010_1;
      patterns[55461] = 25'b11011000_10100011_01111011_1;
      patterns[55462] = 25'b11011000_10100100_01111100_1;
      patterns[55463] = 25'b11011000_10100101_01111101_1;
      patterns[55464] = 25'b11011000_10100110_01111110_1;
      patterns[55465] = 25'b11011000_10100111_01111111_1;
      patterns[55466] = 25'b11011000_10101000_10000000_1;
      patterns[55467] = 25'b11011000_10101001_10000001_1;
      patterns[55468] = 25'b11011000_10101010_10000010_1;
      patterns[55469] = 25'b11011000_10101011_10000011_1;
      patterns[55470] = 25'b11011000_10101100_10000100_1;
      patterns[55471] = 25'b11011000_10101101_10000101_1;
      patterns[55472] = 25'b11011000_10101110_10000110_1;
      patterns[55473] = 25'b11011000_10101111_10000111_1;
      patterns[55474] = 25'b11011000_10110000_10001000_1;
      patterns[55475] = 25'b11011000_10110001_10001001_1;
      patterns[55476] = 25'b11011000_10110010_10001010_1;
      patterns[55477] = 25'b11011000_10110011_10001011_1;
      patterns[55478] = 25'b11011000_10110100_10001100_1;
      patterns[55479] = 25'b11011000_10110101_10001101_1;
      patterns[55480] = 25'b11011000_10110110_10001110_1;
      patterns[55481] = 25'b11011000_10110111_10001111_1;
      patterns[55482] = 25'b11011000_10111000_10010000_1;
      patterns[55483] = 25'b11011000_10111001_10010001_1;
      patterns[55484] = 25'b11011000_10111010_10010010_1;
      patterns[55485] = 25'b11011000_10111011_10010011_1;
      patterns[55486] = 25'b11011000_10111100_10010100_1;
      patterns[55487] = 25'b11011000_10111101_10010101_1;
      patterns[55488] = 25'b11011000_10111110_10010110_1;
      patterns[55489] = 25'b11011000_10111111_10010111_1;
      patterns[55490] = 25'b11011000_11000000_10011000_1;
      patterns[55491] = 25'b11011000_11000001_10011001_1;
      patterns[55492] = 25'b11011000_11000010_10011010_1;
      patterns[55493] = 25'b11011000_11000011_10011011_1;
      patterns[55494] = 25'b11011000_11000100_10011100_1;
      patterns[55495] = 25'b11011000_11000101_10011101_1;
      patterns[55496] = 25'b11011000_11000110_10011110_1;
      patterns[55497] = 25'b11011000_11000111_10011111_1;
      patterns[55498] = 25'b11011000_11001000_10100000_1;
      patterns[55499] = 25'b11011000_11001001_10100001_1;
      patterns[55500] = 25'b11011000_11001010_10100010_1;
      patterns[55501] = 25'b11011000_11001011_10100011_1;
      patterns[55502] = 25'b11011000_11001100_10100100_1;
      patterns[55503] = 25'b11011000_11001101_10100101_1;
      patterns[55504] = 25'b11011000_11001110_10100110_1;
      patterns[55505] = 25'b11011000_11001111_10100111_1;
      patterns[55506] = 25'b11011000_11010000_10101000_1;
      patterns[55507] = 25'b11011000_11010001_10101001_1;
      patterns[55508] = 25'b11011000_11010010_10101010_1;
      patterns[55509] = 25'b11011000_11010011_10101011_1;
      patterns[55510] = 25'b11011000_11010100_10101100_1;
      patterns[55511] = 25'b11011000_11010101_10101101_1;
      patterns[55512] = 25'b11011000_11010110_10101110_1;
      patterns[55513] = 25'b11011000_11010111_10101111_1;
      patterns[55514] = 25'b11011000_11011000_10110000_1;
      patterns[55515] = 25'b11011000_11011001_10110001_1;
      patterns[55516] = 25'b11011000_11011010_10110010_1;
      patterns[55517] = 25'b11011000_11011011_10110011_1;
      patterns[55518] = 25'b11011000_11011100_10110100_1;
      patterns[55519] = 25'b11011000_11011101_10110101_1;
      patterns[55520] = 25'b11011000_11011110_10110110_1;
      patterns[55521] = 25'b11011000_11011111_10110111_1;
      patterns[55522] = 25'b11011000_11100000_10111000_1;
      patterns[55523] = 25'b11011000_11100001_10111001_1;
      patterns[55524] = 25'b11011000_11100010_10111010_1;
      patterns[55525] = 25'b11011000_11100011_10111011_1;
      patterns[55526] = 25'b11011000_11100100_10111100_1;
      patterns[55527] = 25'b11011000_11100101_10111101_1;
      patterns[55528] = 25'b11011000_11100110_10111110_1;
      patterns[55529] = 25'b11011000_11100111_10111111_1;
      patterns[55530] = 25'b11011000_11101000_11000000_1;
      patterns[55531] = 25'b11011000_11101001_11000001_1;
      patterns[55532] = 25'b11011000_11101010_11000010_1;
      patterns[55533] = 25'b11011000_11101011_11000011_1;
      patterns[55534] = 25'b11011000_11101100_11000100_1;
      patterns[55535] = 25'b11011000_11101101_11000101_1;
      patterns[55536] = 25'b11011000_11101110_11000110_1;
      patterns[55537] = 25'b11011000_11101111_11000111_1;
      patterns[55538] = 25'b11011000_11110000_11001000_1;
      patterns[55539] = 25'b11011000_11110001_11001001_1;
      patterns[55540] = 25'b11011000_11110010_11001010_1;
      patterns[55541] = 25'b11011000_11110011_11001011_1;
      patterns[55542] = 25'b11011000_11110100_11001100_1;
      patterns[55543] = 25'b11011000_11110101_11001101_1;
      patterns[55544] = 25'b11011000_11110110_11001110_1;
      patterns[55545] = 25'b11011000_11110111_11001111_1;
      patterns[55546] = 25'b11011000_11111000_11010000_1;
      patterns[55547] = 25'b11011000_11111001_11010001_1;
      patterns[55548] = 25'b11011000_11111010_11010010_1;
      patterns[55549] = 25'b11011000_11111011_11010011_1;
      patterns[55550] = 25'b11011000_11111100_11010100_1;
      patterns[55551] = 25'b11011000_11111101_11010101_1;
      patterns[55552] = 25'b11011000_11111110_11010110_1;
      patterns[55553] = 25'b11011000_11111111_11010111_1;
      patterns[55554] = 25'b11011001_00000000_11011001_0;
      patterns[55555] = 25'b11011001_00000001_11011010_0;
      patterns[55556] = 25'b11011001_00000010_11011011_0;
      patterns[55557] = 25'b11011001_00000011_11011100_0;
      patterns[55558] = 25'b11011001_00000100_11011101_0;
      patterns[55559] = 25'b11011001_00000101_11011110_0;
      patterns[55560] = 25'b11011001_00000110_11011111_0;
      patterns[55561] = 25'b11011001_00000111_11100000_0;
      patterns[55562] = 25'b11011001_00001000_11100001_0;
      patterns[55563] = 25'b11011001_00001001_11100010_0;
      patterns[55564] = 25'b11011001_00001010_11100011_0;
      patterns[55565] = 25'b11011001_00001011_11100100_0;
      patterns[55566] = 25'b11011001_00001100_11100101_0;
      patterns[55567] = 25'b11011001_00001101_11100110_0;
      patterns[55568] = 25'b11011001_00001110_11100111_0;
      patterns[55569] = 25'b11011001_00001111_11101000_0;
      patterns[55570] = 25'b11011001_00010000_11101001_0;
      patterns[55571] = 25'b11011001_00010001_11101010_0;
      patterns[55572] = 25'b11011001_00010010_11101011_0;
      patterns[55573] = 25'b11011001_00010011_11101100_0;
      patterns[55574] = 25'b11011001_00010100_11101101_0;
      patterns[55575] = 25'b11011001_00010101_11101110_0;
      patterns[55576] = 25'b11011001_00010110_11101111_0;
      patterns[55577] = 25'b11011001_00010111_11110000_0;
      patterns[55578] = 25'b11011001_00011000_11110001_0;
      patterns[55579] = 25'b11011001_00011001_11110010_0;
      patterns[55580] = 25'b11011001_00011010_11110011_0;
      patterns[55581] = 25'b11011001_00011011_11110100_0;
      patterns[55582] = 25'b11011001_00011100_11110101_0;
      patterns[55583] = 25'b11011001_00011101_11110110_0;
      patterns[55584] = 25'b11011001_00011110_11110111_0;
      patterns[55585] = 25'b11011001_00011111_11111000_0;
      patterns[55586] = 25'b11011001_00100000_11111001_0;
      patterns[55587] = 25'b11011001_00100001_11111010_0;
      patterns[55588] = 25'b11011001_00100010_11111011_0;
      patterns[55589] = 25'b11011001_00100011_11111100_0;
      patterns[55590] = 25'b11011001_00100100_11111101_0;
      patterns[55591] = 25'b11011001_00100101_11111110_0;
      patterns[55592] = 25'b11011001_00100110_11111111_0;
      patterns[55593] = 25'b11011001_00100111_00000000_1;
      patterns[55594] = 25'b11011001_00101000_00000001_1;
      patterns[55595] = 25'b11011001_00101001_00000010_1;
      patterns[55596] = 25'b11011001_00101010_00000011_1;
      patterns[55597] = 25'b11011001_00101011_00000100_1;
      patterns[55598] = 25'b11011001_00101100_00000101_1;
      patterns[55599] = 25'b11011001_00101101_00000110_1;
      patterns[55600] = 25'b11011001_00101110_00000111_1;
      patterns[55601] = 25'b11011001_00101111_00001000_1;
      patterns[55602] = 25'b11011001_00110000_00001001_1;
      patterns[55603] = 25'b11011001_00110001_00001010_1;
      patterns[55604] = 25'b11011001_00110010_00001011_1;
      patterns[55605] = 25'b11011001_00110011_00001100_1;
      patterns[55606] = 25'b11011001_00110100_00001101_1;
      patterns[55607] = 25'b11011001_00110101_00001110_1;
      patterns[55608] = 25'b11011001_00110110_00001111_1;
      patterns[55609] = 25'b11011001_00110111_00010000_1;
      patterns[55610] = 25'b11011001_00111000_00010001_1;
      patterns[55611] = 25'b11011001_00111001_00010010_1;
      patterns[55612] = 25'b11011001_00111010_00010011_1;
      patterns[55613] = 25'b11011001_00111011_00010100_1;
      patterns[55614] = 25'b11011001_00111100_00010101_1;
      patterns[55615] = 25'b11011001_00111101_00010110_1;
      patterns[55616] = 25'b11011001_00111110_00010111_1;
      patterns[55617] = 25'b11011001_00111111_00011000_1;
      patterns[55618] = 25'b11011001_01000000_00011001_1;
      patterns[55619] = 25'b11011001_01000001_00011010_1;
      patterns[55620] = 25'b11011001_01000010_00011011_1;
      patterns[55621] = 25'b11011001_01000011_00011100_1;
      patterns[55622] = 25'b11011001_01000100_00011101_1;
      patterns[55623] = 25'b11011001_01000101_00011110_1;
      patterns[55624] = 25'b11011001_01000110_00011111_1;
      patterns[55625] = 25'b11011001_01000111_00100000_1;
      patterns[55626] = 25'b11011001_01001000_00100001_1;
      patterns[55627] = 25'b11011001_01001001_00100010_1;
      patterns[55628] = 25'b11011001_01001010_00100011_1;
      patterns[55629] = 25'b11011001_01001011_00100100_1;
      patterns[55630] = 25'b11011001_01001100_00100101_1;
      patterns[55631] = 25'b11011001_01001101_00100110_1;
      patterns[55632] = 25'b11011001_01001110_00100111_1;
      patterns[55633] = 25'b11011001_01001111_00101000_1;
      patterns[55634] = 25'b11011001_01010000_00101001_1;
      patterns[55635] = 25'b11011001_01010001_00101010_1;
      patterns[55636] = 25'b11011001_01010010_00101011_1;
      patterns[55637] = 25'b11011001_01010011_00101100_1;
      patterns[55638] = 25'b11011001_01010100_00101101_1;
      patterns[55639] = 25'b11011001_01010101_00101110_1;
      patterns[55640] = 25'b11011001_01010110_00101111_1;
      patterns[55641] = 25'b11011001_01010111_00110000_1;
      patterns[55642] = 25'b11011001_01011000_00110001_1;
      patterns[55643] = 25'b11011001_01011001_00110010_1;
      patterns[55644] = 25'b11011001_01011010_00110011_1;
      patterns[55645] = 25'b11011001_01011011_00110100_1;
      patterns[55646] = 25'b11011001_01011100_00110101_1;
      patterns[55647] = 25'b11011001_01011101_00110110_1;
      patterns[55648] = 25'b11011001_01011110_00110111_1;
      patterns[55649] = 25'b11011001_01011111_00111000_1;
      patterns[55650] = 25'b11011001_01100000_00111001_1;
      patterns[55651] = 25'b11011001_01100001_00111010_1;
      patterns[55652] = 25'b11011001_01100010_00111011_1;
      patterns[55653] = 25'b11011001_01100011_00111100_1;
      patterns[55654] = 25'b11011001_01100100_00111101_1;
      patterns[55655] = 25'b11011001_01100101_00111110_1;
      patterns[55656] = 25'b11011001_01100110_00111111_1;
      patterns[55657] = 25'b11011001_01100111_01000000_1;
      patterns[55658] = 25'b11011001_01101000_01000001_1;
      patterns[55659] = 25'b11011001_01101001_01000010_1;
      patterns[55660] = 25'b11011001_01101010_01000011_1;
      patterns[55661] = 25'b11011001_01101011_01000100_1;
      patterns[55662] = 25'b11011001_01101100_01000101_1;
      patterns[55663] = 25'b11011001_01101101_01000110_1;
      patterns[55664] = 25'b11011001_01101110_01000111_1;
      patterns[55665] = 25'b11011001_01101111_01001000_1;
      patterns[55666] = 25'b11011001_01110000_01001001_1;
      patterns[55667] = 25'b11011001_01110001_01001010_1;
      patterns[55668] = 25'b11011001_01110010_01001011_1;
      patterns[55669] = 25'b11011001_01110011_01001100_1;
      patterns[55670] = 25'b11011001_01110100_01001101_1;
      patterns[55671] = 25'b11011001_01110101_01001110_1;
      patterns[55672] = 25'b11011001_01110110_01001111_1;
      patterns[55673] = 25'b11011001_01110111_01010000_1;
      patterns[55674] = 25'b11011001_01111000_01010001_1;
      patterns[55675] = 25'b11011001_01111001_01010010_1;
      patterns[55676] = 25'b11011001_01111010_01010011_1;
      patterns[55677] = 25'b11011001_01111011_01010100_1;
      patterns[55678] = 25'b11011001_01111100_01010101_1;
      patterns[55679] = 25'b11011001_01111101_01010110_1;
      patterns[55680] = 25'b11011001_01111110_01010111_1;
      patterns[55681] = 25'b11011001_01111111_01011000_1;
      patterns[55682] = 25'b11011001_10000000_01011001_1;
      patterns[55683] = 25'b11011001_10000001_01011010_1;
      patterns[55684] = 25'b11011001_10000010_01011011_1;
      patterns[55685] = 25'b11011001_10000011_01011100_1;
      patterns[55686] = 25'b11011001_10000100_01011101_1;
      patterns[55687] = 25'b11011001_10000101_01011110_1;
      patterns[55688] = 25'b11011001_10000110_01011111_1;
      patterns[55689] = 25'b11011001_10000111_01100000_1;
      patterns[55690] = 25'b11011001_10001000_01100001_1;
      patterns[55691] = 25'b11011001_10001001_01100010_1;
      patterns[55692] = 25'b11011001_10001010_01100011_1;
      patterns[55693] = 25'b11011001_10001011_01100100_1;
      patterns[55694] = 25'b11011001_10001100_01100101_1;
      patterns[55695] = 25'b11011001_10001101_01100110_1;
      patterns[55696] = 25'b11011001_10001110_01100111_1;
      patterns[55697] = 25'b11011001_10001111_01101000_1;
      patterns[55698] = 25'b11011001_10010000_01101001_1;
      patterns[55699] = 25'b11011001_10010001_01101010_1;
      patterns[55700] = 25'b11011001_10010010_01101011_1;
      patterns[55701] = 25'b11011001_10010011_01101100_1;
      patterns[55702] = 25'b11011001_10010100_01101101_1;
      patterns[55703] = 25'b11011001_10010101_01101110_1;
      patterns[55704] = 25'b11011001_10010110_01101111_1;
      patterns[55705] = 25'b11011001_10010111_01110000_1;
      patterns[55706] = 25'b11011001_10011000_01110001_1;
      patterns[55707] = 25'b11011001_10011001_01110010_1;
      patterns[55708] = 25'b11011001_10011010_01110011_1;
      patterns[55709] = 25'b11011001_10011011_01110100_1;
      patterns[55710] = 25'b11011001_10011100_01110101_1;
      patterns[55711] = 25'b11011001_10011101_01110110_1;
      patterns[55712] = 25'b11011001_10011110_01110111_1;
      patterns[55713] = 25'b11011001_10011111_01111000_1;
      patterns[55714] = 25'b11011001_10100000_01111001_1;
      patterns[55715] = 25'b11011001_10100001_01111010_1;
      patterns[55716] = 25'b11011001_10100010_01111011_1;
      patterns[55717] = 25'b11011001_10100011_01111100_1;
      patterns[55718] = 25'b11011001_10100100_01111101_1;
      patterns[55719] = 25'b11011001_10100101_01111110_1;
      patterns[55720] = 25'b11011001_10100110_01111111_1;
      patterns[55721] = 25'b11011001_10100111_10000000_1;
      patterns[55722] = 25'b11011001_10101000_10000001_1;
      patterns[55723] = 25'b11011001_10101001_10000010_1;
      patterns[55724] = 25'b11011001_10101010_10000011_1;
      patterns[55725] = 25'b11011001_10101011_10000100_1;
      patterns[55726] = 25'b11011001_10101100_10000101_1;
      patterns[55727] = 25'b11011001_10101101_10000110_1;
      patterns[55728] = 25'b11011001_10101110_10000111_1;
      patterns[55729] = 25'b11011001_10101111_10001000_1;
      patterns[55730] = 25'b11011001_10110000_10001001_1;
      patterns[55731] = 25'b11011001_10110001_10001010_1;
      patterns[55732] = 25'b11011001_10110010_10001011_1;
      patterns[55733] = 25'b11011001_10110011_10001100_1;
      patterns[55734] = 25'b11011001_10110100_10001101_1;
      patterns[55735] = 25'b11011001_10110101_10001110_1;
      patterns[55736] = 25'b11011001_10110110_10001111_1;
      patterns[55737] = 25'b11011001_10110111_10010000_1;
      patterns[55738] = 25'b11011001_10111000_10010001_1;
      patterns[55739] = 25'b11011001_10111001_10010010_1;
      patterns[55740] = 25'b11011001_10111010_10010011_1;
      patterns[55741] = 25'b11011001_10111011_10010100_1;
      patterns[55742] = 25'b11011001_10111100_10010101_1;
      patterns[55743] = 25'b11011001_10111101_10010110_1;
      patterns[55744] = 25'b11011001_10111110_10010111_1;
      patterns[55745] = 25'b11011001_10111111_10011000_1;
      patterns[55746] = 25'b11011001_11000000_10011001_1;
      patterns[55747] = 25'b11011001_11000001_10011010_1;
      patterns[55748] = 25'b11011001_11000010_10011011_1;
      patterns[55749] = 25'b11011001_11000011_10011100_1;
      patterns[55750] = 25'b11011001_11000100_10011101_1;
      patterns[55751] = 25'b11011001_11000101_10011110_1;
      patterns[55752] = 25'b11011001_11000110_10011111_1;
      patterns[55753] = 25'b11011001_11000111_10100000_1;
      patterns[55754] = 25'b11011001_11001000_10100001_1;
      patterns[55755] = 25'b11011001_11001001_10100010_1;
      patterns[55756] = 25'b11011001_11001010_10100011_1;
      patterns[55757] = 25'b11011001_11001011_10100100_1;
      patterns[55758] = 25'b11011001_11001100_10100101_1;
      patterns[55759] = 25'b11011001_11001101_10100110_1;
      patterns[55760] = 25'b11011001_11001110_10100111_1;
      patterns[55761] = 25'b11011001_11001111_10101000_1;
      patterns[55762] = 25'b11011001_11010000_10101001_1;
      patterns[55763] = 25'b11011001_11010001_10101010_1;
      patterns[55764] = 25'b11011001_11010010_10101011_1;
      patterns[55765] = 25'b11011001_11010011_10101100_1;
      patterns[55766] = 25'b11011001_11010100_10101101_1;
      patterns[55767] = 25'b11011001_11010101_10101110_1;
      patterns[55768] = 25'b11011001_11010110_10101111_1;
      patterns[55769] = 25'b11011001_11010111_10110000_1;
      patterns[55770] = 25'b11011001_11011000_10110001_1;
      patterns[55771] = 25'b11011001_11011001_10110010_1;
      patterns[55772] = 25'b11011001_11011010_10110011_1;
      patterns[55773] = 25'b11011001_11011011_10110100_1;
      patterns[55774] = 25'b11011001_11011100_10110101_1;
      patterns[55775] = 25'b11011001_11011101_10110110_1;
      patterns[55776] = 25'b11011001_11011110_10110111_1;
      patterns[55777] = 25'b11011001_11011111_10111000_1;
      patterns[55778] = 25'b11011001_11100000_10111001_1;
      patterns[55779] = 25'b11011001_11100001_10111010_1;
      patterns[55780] = 25'b11011001_11100010_10111011_1;
      patterns[55781] = 25'b11011001_11100011_10111100_1;
      patterns[55782] = 25'b11011001_11100100_10111101_1;
      patterns[55783] = 25'b11011001_11100101_10111110_1;
      patterns[55784] = 25'b11011001_11100110_10111111_1;
      patterns[55785] = 25'b11011001_11100111_11000000_1;
      patterns[55786] = 25'b11011001_11101000_11000001_1;
      patterns[55787] = 25'b11011001_11101001_11000010_1;
      patterns[55788] = 25'b11011001_11101010_11000011_1;
      patterns[55789] = 25'b11011001_11101011_11000100_1;
      patterns[55790] = 25'b11011001_11101100_11000101_1;
      patterns[55791] = 25'b11011001_11101101_11000110_1;
      patterns[55792] = 25'b11011001_11101110_11000111_1;
      patterns[55793] = 25'b11011001_11101111_11001000_1;
      patterns[55794] = 25'b11011001_11110000_11001001_1;
      patterns[55795] = 25'b11011001_11110001_11001010_1;
      patterns[55796] = 25'b11011001_11110010_11001011_1;
      patterns[55797] = 25'b11011001_11110011_11001100_1;
      patterns[55798] = 25'b11011001_11110100_11001101_1;
      patterns[55799] = 25'b11011001_11110101_11001110_1;
      patterns[55800] = 25'b11011001_11110110_11001111_1;
      patterns[55801] = 25'b11011001_11110111_11010000_1;
      patterns[55802] = 25'b11011001_11111000_11010001_1;
      patterns[55803] = 25'b11011001_11111001_11010010_1;
      patterns[55804] = 25'b11011001_11111010_11010011_1;
      patterns[55805] = 25'b11011001_11111011_11010100_1;
      patterns[55806] = 25'b11011001_11111100_11010101_1;
      patterns[55807] = 25'b11011001_11111101_11010110_1;
      patterns[55808] = 25'b11011001_11111110_11010111_1;
      patterns[55809] = 25'b11011001_11111111_11011000_1;
      patterns[55810] = 25'b11011010_00000000_11011010_0;
      patterns[55811] = 25'b11011010_00000001_11011011_0;
      patterns[55812] = 25'b11011010_00000010_11011100_0;
      patterns[55813] = 25'b11011010_00000011_11011101_0;
      patterns[55814] = 25'b11011010_00000100_11011110_0;
      patterns[55815] = 25'b11011010_00000101_11011111_0;
      patterns[55816] = 25'b11011010_00000110_11100000_0;
      patterns[55817] = 25'b11011010_00000111_11100001_0;
      patterns[55818] = 25'b11011010_00001000_11100010_0;
      patterns[55819] = 25'b11011010_00001001_11100011_0;
      patterns[55820] = 25'b11011010_00001010_11100100_0;
      patterns[55821] = 25'b11011010_00001011_11100101_0;
      patterns[55822] = 25'b11011010_00001100_11100110_0;
      patterns[55823] = 25'b11011010_00001101_11100111_0;
      patterns[55824] = 25'b11011010_00001110_11101000_0;
      patterns[55825] = 25'b11011010_00001111_11101001_0;
      patterns[55826] = 25'b11011010_00010000_11101010_0;
      patterns[55827] = 25'b11011010_00010001_11101011_0;
      patterns[55828] = 25'b11011010_00010010_11101100_0;
      patterns[55829] = 25'b11011010_00010011_11101101_0;
      patterns[55830] = 25'b11011010_00010100_11101110_0;
      patterns[55831] = 25'b11011010_00010101_11101111_0;
      patterns[55832] = 25'b11011010_00010110_11110000_0;
      patterns[55833] = 25'b11011010_00010111_11110001_0;
      patterns[55834] = 25'b11011010_00011000_11110010_0;
      patterns[55835] = 25'b11011010_00011001_11110011_0;
      patterns[55836] = 25'b11011010_00011010_11110100_0;
      patterns[55837] = 25'b11011010_00011011_11110101_0;
      patterns[55838] = 25'b11011010_00011100_11110110_0;
      patterns[55839] = 25'b11011010_00011101_11110111_0;
      patterns[55840] = 25'b11011010_00011110_11111000_0;
      patterns[55841] = 25'b11011010_00011111_11111001_0;
      patterns[55842] = 25'b11011010_00100000_11111010_0;
      patterns[55843] = 25'b11011010_00100001_11111011_0;
      patterns[55844] = 25'b11011010_00100010_11111100_0;
      patterns[55845] = 25'b11011010_00100011_11111101_0;
      patterns[55846] = 25'b11011010_00100100_11111110_0;
      patterns[55847] = 25'b11011010_00100101_11111111_0;
      patterns[55848] = 25'b11011010_00100110_00000000_1;
      patterns[55849] = 25'b11011010_00100111_00000001_1;
      patterns[55850] = 25'b11011010_00101000_00000010_1;
      patterns[55851] = 25'b11011010_00101001_00000011_1;
      patterns[55852] = 25'b11011010_00101010_00000100_1;
      patterns[55853] = 25'b11011010_00101011_00000101_1;
      patterns[55854] = 25'b11011010_00101100_00000110_1;
      patterns[55855] = 25'b11011010_00101101_00000111_1;
      patterns[55856] = 25'b11011010_00101110_00001000_1;
      patterns[55857] = 25'b11011010_00101111_00001001_1;
      patterns[55858] = 25'b11011010_00110000_00001010_1;
      patterns[55859] = 25'b11011010_00110001_00001011_1;
      patterns[55860] = 25'b11011010_00110010_00001100_1;
      patterns[55861] = 25'b11011010_00110011_00001101_1;
      patterns[55862] = 25'b11011010_00110100_00001110_1;
      patterns[55863] = 25'b11011010_00110101_00001111_1;
      patterns[55864] = 25'b11011010_00110110_00010000_1;
      patterns[55865] = 25'b11011010_00110111_00010001_1;
      patterns[55866] = 25'b11011010_00111000_00010010_1;
      patterns[55867] = 25'b11011010_00111001_00010011_1;
      patterns[55868] = 25'b11011010_00111010_00010100_1;
      patterns[55869] = 25'b11011010_00111011_00010101_1;
      patterns[55870] = 25'b11011010_00111100_00010110_1;
      patterns[55871] = 25'b11011010_00111101_00010111_1;
      patterns[55872] = 25'b11011010_00111110_00011000_1;
      patterns[55873] = 25'b11011010_00111111_00011001_1;
      patterns[55874] = 25'b11011010_01000000_00011010_1;
      patterns[55875] = 25'b11011010_01000001_00011011_1;
      patterns[55876] = 25'b11011010_01000010_00011100_1;
      patterns[55877] = 25'b11011010_01000011_00011101_1;
      patterns[55878] = 25'b11011010_01000100_00011110_1;
      patterns[55879] = 25'b11011010_01000101_00011111_1;
      patterns[55880] = 25'b11011010_01000110_00100000_1;
      patterns[55881] = 25'b11011010_01000111_00100001_1;
      patterns[55882] = 25'b11011010_01001000_00100010_1;
      patterns[55883] = 25'b11011010_01001001_00100011_1;
      patterns[55884] = 25'b11011010_01001010_00100100_1;
      patterns[55885] = 25'b11011010_01001011_00100101_1;
      patterns[55886] = 25'b11011010_01001100_00100110_1;
      patterns[55887] = 25'b11011010_01001101_00100111_1;
      patterns[55888] = 25'b11011010_01001110_00101000_1;
      patterns[55889] = 25'b11011010_01001111_00101001_1;
      patterns[55890] = 25'b11011010_01010000_00101010_1;
      patterns[55891] = 25'b11011010_01010001_00101011_1;
      patterns[55892] = 25'b11011010_01010010_00101100_1;
      patterns[55893] = 25'b11011010_01010011_00101101_1;
      patterns[55894] = 25'b11011010_01010100_00101110_1;
      patterns[55895] = 25'b11011010_01010101_00101111_1;
      patterns[55896] = 25'b11011010_01010110_00110000_1;
      patterns[55897] = 25'b11011010_01010111_00110001_1;
      patterns[55898] = 25'b11011010_01011000_00110010_1;
      patterns[55899] = 25'b11011010_01011001_00110011_1;
      patterns[55900] = 25'b11011010_01011010_00110100_1;
      patterns[55901] = 25'b11011010_01011011_00110101_1;
      patterns[55902] = 25'b11011010_01011100_00110110_1;
      patterns[55903] = 25'b11011010_01011101_00110111_1;
      patterns[55904] = 25'b11011010_01011110_00111000_1;
      patterns[55905] = 25'b11011010_01011111_00111001_1;
      patterns[55906] = 25'b11011010_01100000_00111010_1;
      patterns[55907] = 25'b11011010_01100001_00111011_1;
      patterns[55908] = 25'b11011010_01100010_00111100_1;
      patterns[55909] = 25'b11011010_01100011_00111101_1;
      patterns[55910] = 25'b11011010_01100100_00111110_1;
      patterns[55911] = 25'b11011010_01100101_00111111_1;
      patterns[55912] = 25'b11011010_01100110_01000000_1;
      patterns[55913] = 25'b11011010_01100111_01000001_1;
      patterns[55914] = 25'b11011010_01101000_01000010_1;
      patterns[55915] = 25'b11011010_01101001_01000011_1;
      patterns[55916] = 25'b11011010_01101010_01000100_1;
      patterns[55917] = 25'b11011010_01101011_01000101_1;
      patterns[55918] = 25'b11011010_01101100_01000110_1;
      patterns[55919] = 25'b11011010_01101101_01000111_1;
      patterns[55920] = 25'b11011010_01101110_01001000_1;
      patterns[55921] = 25'b11011010_01101111_01001001_1;
      patterns[55922] = 25'b11011010_01110000_01001010_1;
      patterns[55923] = 25'b11011010_01110001_01001011_1;
      patterns[55924] = 25'b11011010_01110010_01001100_1;
      patterns[55925] = 25'b11011010_01110011_01001101_1;
      patterns[55926] = 25'b11011010_01110100_01001110_1;
      patterns[55927] = 25'b11011010_01110101_01001111_1;
      patterns[55928] = 25'b11011010_01110110_01010000_1;
      patterns[55929] = 25'b11011010_01110111_01010001_1;
      patterns[55930] = 25'b11011010_01111000_01010010_1;
      patterns[55931] = 25'b11011010_01111001_01010011_1;
      patterns[55932] = 25'b11011010_01111010_01010100_1;
      patterns[55933] = 25'b11011010_01111011_01010101_1;
      patterns[55934] = 25'b11011010_01111100_01010110_1;
      patterns[55935] = 25'b11011010_01111101_01010111_1;
      patterns[55936] = 25'b11011010_01111110_01011000_1;
      patterns[55937] = 25'b11011010_01111111_01011001_1;
      patterns[55938] = 25'b11011010_10000000_01011010_1;
      patterns[55939] = 25'b11011010_10000001_01011011_1;
      patterns[55940] = 25'b11011010_10000010_01011100_1;
      patterns[55941] = 25'b11011010_10000011_01011101_1;
      patterns[55942] = 25'b11011010_10000100_01011110_1;
      patterns[55943] = 25'b11011010_10000101_01011111_1;
      patterns[55944] = 25'b11011010_10000110_01100000_1;
      patterns[55945] = 25'b11011010_10000111_01100001_1;
      patterns[55946] = 25'b11011010_10001000_01100010_1;
      patterns[55947] = 25'b11011010_10001001_01100011_1;
      patterns[55948] = 25'b11011010_10001010_01100100_1;
      patterns[55949] = 25'b11011010_10001011_01100101_1;
      patterns[55950] = 25'b11011010_10001100_01100110_1;
      patterns[55951] = 25'b11011010_10001101_01100111_1;
      patterns[55952] = 25'b11011010_10001110_01101000_1;
      patterns[55953] = 25'b11011010_10001111_01101001_1;
      patterns[55954] = 25'b11011010_10010000_01101010_1;
      patterns[55955] = 25'b11011010_10010001_01101011_1;
      patterns[55956] = 25'b11011010_10010010_01101100_1;
      patterns[55957] = 25'b11011010_10010011_01101101_1;
      patterns[55958] = 25'b11011010_10010100_01101110_1;
      patterns[55959] = 25'b11011010_10010101_01101111_1;
      patterns[55960] = 25'b11011010_10010110_01110000_1;
      patterns[55961] = 25'b11011010_10010111_01110001_1;
      patterns[55962] = 25'b11011010_10011000_01110010_1;
      patterns[55963] = 25'b11011010_10011001_01110011_1;
      patterns[55964] = 25'b11011010_10011010_01110100_1;
      patterns[55965] = 25'b11011010_10011011_01110101_1;
      patterns[55966] = 25'b11011010_10011100_01110110_1;
      patterns[55967] = 25'b11011010_10011101_01110111_1;
      patterns[55968] = 25'b11011010_10011110_01111000_1;
      patterns[55969] = 25'b11011010_10011111_01111001_1;
      patterns[55970] = 25'b11011010_10100000_01111010_1;
      patterns[55971] = 25'b11011010_10100001_01111011_1;
      patterns[55972] = 25'b11011010_10100010_01111100_1;
      patterns[55973] = 25'b11011010_10100011_01111101_1;
      patterns[55974] = 25'b11011010_10100100_01111110_1;
      patterns[55975] = 25'b11011010_10100101_01111111_1;
      patterns[55976] = 25'b11011010_10100110_10000000_1;
      patterns[55977] = 25'b11011010_10100111_10000001_1;
      patterns[55978] = 25'b11011010_10101000_10000010_1;
      patterns[55979] = 25'b11011010_10101001_10000011_1;
      patterns[55980] = 25'b11011010_10101010_10000100_1;
      patterns[55981] = 25'b11011010_10101011_10000101_1;
      patterns[55982] = 25'b11011010_10101100_10000110_1;
      patterns[55983] = 25'b11011010_10101101_10000111_1;
      patterns[55984] = 25'b11011010_10101110_10001000_1;
      patterns[55985] = 25'b11011010_10101111_10001001_1;
      patterns[55986] = 25'b11011010_10110000_10001010_1;
      patterns[55987] = 25'b11011010_10110001_10001011_1;
      patterns[55988] = 25'b11011010_10110010_10001100_1;
      patterns[55989] = 25'b11011010_10110011_10001101_1;
      patterns[55990] = 25'b11011010_10110100_10001110_1;
      patterns[55991] = 25'b11011010_10110101_10001111_1;
      patterns[55992] = 25'b11011010_10110110_10010000_1;
      patterns[55993] = 25'b11011010_10110111_10010001_1;
      patterns[55994] = 25'b11011010_10111000_10010010_1;
      patterns[55995] = 25'b11011010_10111001_10010011_1;
      patterns[55996] = 25'b11011010_10111010_10010100_1;
      patterns[55997] = 25'b11011010_10111011_10010101_1;
      patterns[55998] = 25'b11011010_10111100_10010110_1;
      patterns[55999] = 25'b11011010_10111101_10010111_1;
      patterns[56000] = 25'b11011010_10111110_10011000_1;
      patterns[56001] = 25'b11011010_10111111_10011001_1;
      patterns[56002] = 25'b11011010_11000000_10011010_1;
      patterns[56003] = 25'b11011010_11000001_10011011_1;
      patterns[56004] = 25'b11011010_11000010_10011100_1;
      patterns[56005] = 25'b11011010_11000011_10011101_1;
      patterns[56006] = 25'b11011010_11000100_10011110_1;
      patterns[56007] = 25'b11011010_11000101_10011111_1;
      patterns[56008] = 25'b11011010_11000110_10100000_1;
      patterns[56009] = 25'b11011010_11000111_10100001_1;
      patterns[56010] = 25'b11011010_11001000_10100010_1;
      patterns[56011] = 25'b11011010_11001001_10100011_1;
      patterns[56012] = 25'b11011010_11001010_10100100_1;
      patterns[56013] = 25'b11011010_11001011_10100101_1;
      patterns[56014] = 25'b11011010_11001100_10100110_1;
      patterns[56015] = 25'b11011010_11001101_10100111_1;
      patterns[56016] = 25'b11011010_11001110_10101000_1;
      patterns[56017] = 25'b11011010_11001111_10101001_1;
      patterns[56018] = 25'b11011010_11010000_10101010_1;
      patterns[56019] = 25'b11011010_11010001_10101011_1;
      patterns[56020] = 25'b11011010_11010010_10101100_1;
      patterns[56021] = 25'b11011010_11010011_10101101_1;
      patterns[56022] = 25'b11011010_11010100_10101110_1;
      patterns[56023] = 25'b11011010_11010101_10101111_1;
      patterns[56024] = 25'b11011010_11010110_10110000_1;
      patterns[56025] = 25'b11011010_11010111_10110001_1;
      patterns[56026] = 25'b11011010_11011000_10110010_1;
      patterns[56027] = 25'b11011010_11011001_10110011_1;
      patterns[56028] = 25'b11011010_11011010_10110100_1;
      patterns[56029] = 25'b11011010_11011011_10110101_1;
      patterns[56030] = 25'b11011010_11011100_10110110_1;
      patterns[56031] = 25'b11011010_11011101_10110111_1;
      patterns[56032] = 25'b11011010_11011110_10111000_1;
      patterns[56033] = 25'b11011010_11011111_10111001_1;
      patterns[56034] = 25'b11011010_11100000_10111010_1;
      patterns[56035] = 25'b11011010_11100001_10111011_1;
      patterns[56036] = 25'b11011010_11100010_10111100_1;
      patterns[56037] = 25'b11011010_11100011_10111101_1;
      patterns[56038] = 25'b11011010_11100100_10111110_1;
      patterns[56039] = 25'b11011010_11100101_10111111_1;
      patterns[56040] = 25'b11011010_11100110_11000000_1;
      patterns[56041] = 25'b11011010_11100111_11000001_1;
      patterns[56042] = 25'b11011010_11101000_11000010_1;
      patterns[56043] = 25'b11011010_11101001_11000011_1;
      patterns[56044] = 25'b11011010_11101010_11000100_1;
      patterns[56045] = 25'b11011010_11101011_11000101_1;
      patterns[56046] = 25'b11011010_11101100_11000110_1;
      patterns[56047] = 25'b11011010_11101101_11000111_1;
      patterns[56048] = 25'b11011010_11101110_11001000_1;
      patterns[56049] = 25'b11011010_11101111_11001001_1;
      patterns[56050] = 25'b11011010_11110000_11001010_1;
      patterns[56051] = 25'b11011010_11110001_11001011_1;
      patterns[56052] = 25'b11011010_11110010_11001100_1;
      patterns[56053] = 25'b11011010_11110011_11001101_1;
      patterns[56054] = 25'b11011010_11110100_11001110_1;
      patterns[56055] = 25'b11011010_11110101_11001111_1;
      patterns[56056] = 25'b11011010_11110110_11010000_1;
      patterns[56057] = 25'b11011010_11110111_11010001_1;
      patterns[56058] = 25'b11011010_11111000_11010010_1;
      patterns[56059] = 25'b11011010_11111001_11010011_1;
      patterns[56060] = 25'b11011010_11111010_11010100_1;
      patterns[56061] = 25'b11011010_11111011_11010101_1;
      patterns[56062] = 25'b11011010_11111100_11010110_1;
      patterns[56063] = 25'b11011010_11111101_11010111_1;
      patterns[56064] = 25'b11011010_11111110_11011000_1;
      patterns[56065] = 25'b11011010_11111111_11011001_1;
      patterns[56066] = 25'b11011011_00000000_11011011_0;
      patterns[56067] = 25'b11011011_00000001_11011100_0;
      patterns[56068] = 25'b11011011_00000010_11011101_0;
      patterns[56069] = 25'b11011011_00000011_11011110_0;
      patterns[56070] = 25'b11011011_00000100_11011111_0;
      patterns[56071] = 25'b11011011_00000101_11100000_0;
      patterns[56072] = 25'b11011011_00000110_11100001_0;
      patterns[56073] = 25'b11011011_00000111_11100010_0;
      patterns[56074] = 25'b11011011_00001000_11100011_0;
      patterns[56075] = 25'b11011011_00001001_11100100_0;
      patterns[56076] = 25'b11011011_00001010_11100101_0;
      patterns[56077] = 25'b11011011_00001011_11100110_0;
      patterns[56078] = 25'b11011011_00001100_11100111_0;
      patterns[56079] = 25'b11011011_00001101_11101000_0;
      patterns[56080] = 25'b11011011_00001110_11101001_0;
      patterns[56081] = 25'b11011011_00001111_11101010_0;
      patterns[56082] = 25'b11011011_00010000_11101011_0;
      patterns[56083] = 25'b11011011_00010001_11101100_0;
      patterns[56084] = 25'b11011011_00010010_11101101_0;
      patterns[56085] = 25'b11011011_00010011_11101110_0;
      patterns[56086] = 25'b11011011_00010100_11101111_0;
      patterns[56087] = 25'b11011011_00010101_11110000_0;
      patterns[56088] = 25'b11011011_00010110_11110001_0;
      patterns[56089] = 25'b11011011_00010111_11110010_0;
      patterns[56090] = 25'b11011011_00011000_11110011_0;
      patterns[56091] = 25'b11011011_00011001_11110100_0;
      patterns[56092] = 25'b11011011_00011010_11110101_0;
      patterns[56093] = 25'b11011011_00011011_11110110_0;
      patterns[56094] = 25'b11011011_00011100_11110111_0;
      patterns[56095] = 25'b11011011_00011101_11111000_0;
      patterns[56096] = 25'b11011011_00011110_11111001_0;
      patterns[56097] = 25'b11011011_00011111_11111010_0;
      patterns[56098] = 25'b11011011_00100000_11111011_0;
      patterns[56099] = 25'b11011011_00100001_11111100_0;
      patterns[56100] = 25'b11011011_00100010_11111101_0;
      patterns[56101] = 25'b11011011_00100011_11111110_0;
      patterns[56102] = 25'b11011011_00100100_11111111_0;
      patterns[56103] = 25'b11011011_00100101_00000000_1;
      patterns[56104] = 25'b11011011_00100110_00000001_1;
      patterns[56105] = 25'b11011011_00100111_00000010_1;
      patterns[56106] = 25'b11011011_00101000_00000011_1;
      patterns[56107] = 25'b11011011_00101001_00000100_1;
      patterns[56108] = 25'b11011011_00101010_00000101_1;
      patterns[56109] = 25'b11011011_00101011_00000110_1;
      patterns[56110] = 25'b11011011_00101100_00000111_1;
      patterns[56111] = 25'b11011011_00101101_00001000_1;
      patterns[56112] = 25'b11011011_00101110_00001001_1;
      patterns[56113] = 25'b11011011_00101111_00001010_1;
      patterns[56114] = 25'b11011011_00110000_00001011_1;
      patterns[56115] = 25'b11011011_00110001_00001100_1;
      patterns[56116] = 25'b11011011_00110010_00001101_1;
      patterns[56117] = 25'b11011011_00110011_00001110_1;
      patterns[56118] = 25'b11011011_00110100_00001111_1;
      patterns[56119] = 25'b11011011_00110101_00010000_1;
      patterns[56120] = 25'b11011011_00110110_00010001_1;
      patterns[56121] = 25'b11011011_00110111_00010010_1;
      patterns[56122] = 25'b11011011_00111000_00010011_1;
      patterns[56123] = 25'b11011011_00111001_00010100_1;
      patterns[56124] = 25'b11011011_00111010_00010101_1;
      patterns[56125] = 25'b11011011_00111011_00010110_1;
      patterns[56126] = 25'b11011011_00111100_00010111_1;
      patterns[56127] = 25'b11011011_00111101_00011000_1;
      patterns[56128] = 25'b11011011_00111110_00011001_1;
      patterns[56129] = 25'b11011011_00111111_00011010_1;
      patterns[56130] = 25'b11011011_01000000_00011011_1;
      patterns[56131] = 25'b11011011_01000001_00011100_1;
      patterns[56132] = 25'b11011011_01000010_00011101_1;
      patterns[56133] = 25'b11011011_01000011_00011110_1;
      patterns[56134] = 25'b11011011_01000100_00011111_1;
      patterns[56135] = 25'b11011011_01000101_00100000_1;
      patterns[56136] = 25'b11011011_01000110_00100001_1;
      patterns[56137] = 25'b11011011_01000111_00100010_1;
      patterns[56138] = 25'b11011011_01001000_00100011_1;
      patterns[56139] = 25'b11011011_01001001_00100100_1;
      patterns[56140] = 25'b11011011_01001010_00100101_1;
      patterns[56141] = 25'b11011011_01001011_00100110_1;
      patterns[56142] = 25'b11011011_01001100_00100111_1;
      patterns[56143] = 25'b11011011_01001101_00101000_1;
      patterns[56144] = 25'b11011011_01001110_00101001_1;
      patterns[56145] = 25'b11011011_01001111_00101010_1;
      patterns[56146] = 25'b11011011_01010000_00101011_1;
      patterns[56147] = 25'b11011011_01010001_00101100_1;
      patterns[56148] = 25'b11011011_01010010_00101101_1;
      patterns[56149] = 25'b11011011_01010011_00101110_1;
      patterns[56150] = 25'b11011011_01010100_00101111_1;
      patterns[56151] = 25'b11011011_01010101_00110000_1;
      patterns[56152] = 25'b11011011_01010110_00110001_1;
      patterns[56153] = 25'b11011011_01010111_00110010_1;
      patterns[56154] = 25'b11011011_01011000_00110011_1;
      patterns[56155] = 25'b11011011_01011001_00110100_1;
      patterns[56156] = 25'b11011011_01011010_00110101_1;
      patterns[56157] = 25'b11011011_01011011_00110110_1;
      patterns[56158] = 25'b11011011_01011100_00110111_1;
      patterns[56159] = 25'b11011011_01011101_00111000_1;
      patterns[56160] = 25'b11011011_01011110_00111001_1;
      patterns[56161] = 25'b11011011_01011111_00111010_1;
      patterns[56162] = 25'b11011011_01100000_00111011_1;
      patterns[56163] = 25'b11011011_01100001_00111100_1;
      patterns[56164] = 25'b11011011_01100010_00111101_1;
      patterns[56165] = 25'b11011011_01100011_00111110_1;
      patterns[56166] = 25'b11011011_01100100_00111111_1;
      patterns[56167] = 25'b11011011_01100101_01000000_1;
      patterns[56168] = 25'b11011011_01100110_01000001_1;
      patterns[56169] = 25'b11011011_01100111_01000010_1;
      patterns[56170] = 25'b11011011_01101000_01000011_1;
      patterns[56171] = 25'b11011011_01101001_01000100_1;
      patterns[56172] = 25'b11011011_01101010_01000101_1;
      patterns[56173] = 25'b11011011_01101011_01000110_1;
      patterns[56174] = 25'b11011011_01101100_01000111_1;
      patterns[56175] = 25'b11011011_01101101_01001000_1;
      patterns[56176] = 25'b11011011_01101110_01001001_1;
      patterns[56177] = 25'b11011011_01101111_01001010_1;
      patterns[56178] = 25'b11011011_01110000_01001011_1;
      patterns[56179] = 25'b11011011_01110001_01001100_1;
      patterns[56180] = 25'b11011011_01110010_01001101_1;
      patterns[56181] = 25'b11011011_01110011_01001110_1;
      patterns[56182] = 25'b11011011_01110100_01001111_1;
      patterns[56183] = 25'b11011011_01110101_01010000_1;
      patterns[56184] = 25'b11011011_01110110_01010001_1;
      patterns[56185] = 25'b11011011_01110111_01010010_1;
      patterns[56186] = 25'b11011011_01111000_01010011_1;
      patterns[56187] = 25'b11011011_01111001_01010100_1;
      patterns[56188] = 25'b11011011_01111010_01010101_1;
      patterns[56189] = 25'b11011011_01111011_01010110_1;
      patterns[56190] = 25'b11011011_01111100_01010111_1;
      patterns[56191] = 25'b11011011_01111101_01011000_1;
      patterns[56192] = 25'b11011011_01111110_01011001_1;
      patterns[56193] = 25'b11011011_01111111_01011010_1;
      patterns[56194] = 25'b11011011_10000000_01011011_1;
      patterns[56195] = 25'b11011011_10000001_01011100_1;
      patterns[56196] = 25'b11011011_10000010_01011101_1;
      patterns[56197] = 25'b11011011_10000011_01011110_1;
      patterns[56198] = 25'b11011011_10000100_01011111_1;
      patterns[56199] = 25'b11011011_10000101_01100000_1;
      patterns[56200] = 25'b11011011_10000110_01100001_1;
      patterns[56201] = 25'b11011011_10000111_01100010_1;
      patterns[56202] = 25'b11011011_10001000_01100011_1;
      patterns[56203] = 25'b11011011_10001001_01100100_1;
      patterns[56204] = 25'b11011011_10001010_01100101_1;
      patterns[56205] = 25'b11011011_10001011_01100110_1;
      patterns[56206] = 25'b11011011_10001100_01100111_1;
      patterns[56207] = 25'b11011011_10001101_01101000_1;
      patterns[56208] = 25'b11011011_10001110_01101001_1;
      patterns[56209] = 25'b11011011_10001111_01101010_1;
      patterns[56210] = 25'b11011011_10010000_01101011_1;
      patterns[56211] = 25'b11011011_10010001_01101100_1;
      patterns[56212] = 25'b11011011_10010010_01101101_1;
      patterns[56213] = 25'b11011011_10010011_01101110_1;
      patterns[56214] = 25'b11011011_10010100_01101111_1;
      patterns[56215] = 25'b11011011_10010101_01110000_1;
      patterns[56216] = 25'b11011011_10010110_01110001_1;
      patterns[56217] = 25'b11011011_10010111_01110010_1;
      patterns[56218] = 25'b11011011_10011000_01110011_1;
      patterns[56219] = 25'b11011011_10011001_01110100_1;
      patterns[56220] = 25'b11011011_10011010_01110101_1;
      patterns[56221] = 25'b11011011_10011011_01110110_1;
      patterns[56222] = 25'b11011011_10011100_01110111_1;
      patterns[56223] = 25'b11011011_10011101_01111000_1;
      patterns[56224] = 25'b11011011_10011110_01111001_1;
      patterns[56225] = 25'b11011011_10011111_01111010_1;
      patterns[56226] = 25'b11011011_10100000_01111011_1;
      patterns[56227] = 25'b11011011_10100001_01111100_1;
      patterns[56228] = 25'b11011011_10100010_01111101_1;
      patterns[56229] = 25'b11011011_10100011_01111110_1;
      patterns[56230] = 25'b11011011_10100100_01111111_1;
      patterns[56231] = 25'b11011011_10100101_10000000_1;
      patterns[56232] = 25'b11011011_10100110_10000001_1;
      patterns[56233] = 25'b11011011_10100111_10000010_1;
      patterns[56234] = 25'b11011011_10101000_10000011_1;
      patterns[56235] = 25'b11011011_10101001_10000100_1;
      patterns[56236] = 25'b11011011_10101010_10000101_1;
      patterns[56237] = 25'b11011011_10101011_10000110_1;
      patterns[56238] = 25'b11011011_10101100_10000111_1;
      patterns[56239] = 25'b11011011_10101101_10001000_1;
      patterns[56240] = 25'b11011011_10101110_10001001_1;
      patterns[56241] = 25'b11011011_10101111_10001010_1;
      patterns[56242] = 25'b11011011_10110000_10001011_1;
      patterns[56243] = 25'b11011011_10110001_10001100_1;
      patterns[56244] = 25'b11011011_10110010_10001101_1;
      patterns[56245] = 25'b11011011_10110011_10001110_1;
      patterns[56246] = 25'b11011011_10110100_10001111_1;
      patterns[56247] = 25'b11011011_10110101_10010000_1;
      patterns[56248] = 25'b11011011_10110110_10010001_1;
      patterns[56249] = 25'b11011011_10110111_10010010_1;
      patterns[56250] = 25'b11011011_10111000_10010011_1;
      patterns[56251] = 25'b11011011_10111001_10010100_1;
      patterns[56252] = 25'b11011011_10111010_10010101_1;
      patterns[56253] = 25'b11011011_10111011_10010110_1;
      patterns[56254] = 25'b11011011_10111100_10010111_1;
      patterns[56255] = 25'b11011011_10111101_10011000_1;
      patterns[56256] = 25'b11011011_10111110_10011001_1;
      patterns[56257] = 25'b11011011_10111111_10011010_1;
      patterns[56258] = 25'b11011011_11000000_10011011_1;
      patterns[56259] = 25'b11011011_11000001_10011100_1;
      patterns[56260] = 25'b11011011_11000010_10011101_1;
      patterns[56261] = 25'b11011011_11000011_10011110_1;
      patterns[56262] = 25'b11011011_11000100_10011111_1;
      patterns[56263] = 25'b11011011_11000101_10100000_1;
      patterns[56264] = 25'b11011011_11000110_10100001_1;
      patterns[56265] = 25'b11011011_11000111_10100010_1;
      patterns[56266] = 25'b11011011_11001000_10100011_1;
      patterns[56267] = 25'b11011011_11001001_10100100_1;
      patterns[56268] = 25'b11011011_11001010_10100101_1;
      patterns[56269] = 25'b11011011_11001011_10100110_1;
      patterns[56270] = 25'b11011011_11001100_10100111_1;
      patterns[56271] = 25'b11011011_11001101_10101000_1;
      patterns[56272] = 25'b11011011_11001110_10101001_1;
      patterns[56273] = 25'b11011011_11001111_10101010_1;
      patterns[56274] = 25'b11011011_11010000_10101011_1;
      patterns[56275] = 25'b11011011_11010001_10101100_1;
      patterns[56276] = 25'b11011011_11010010_10101101_1;
      patterns[56277] = 25'b11011011_11010011_10101110_1;
      patterns[56278] = 25'b11011011_11010100_10101111_1;
      patterns[56279] = 25'b11011011_11010101_10110000_1;
      patterns[56280] = 25'b11011011_11010110_10110001_1;
      patterns[56281] = 25'b11011011_11010111_10110010_1;
      patterns[56282] = 25'b11011011_11011000_10110011_1;
      patterns[56283] = 25'b11011011_11011001_10110100_1;
      patterns[56284] = 25'b11011011_11011010_10110101_1;
      patterns[56285] = 25'b11011011_11011011_10110110_1;
      patterns[56286] = 25'b11011011_11011100_10110111_1;
      patterns[56287] = 25'b11011011_11011101_10111000_1;
      patterns[56288] = 25'b11011011_11011110_10111001_1;
      patterns[56289] = 25'b11011011_11011111_10111010_1;
      patterns[56290] = 25'b11011011_11100000_10111011_1;
      patterns[56291] = 25'b11011011_11100001_10111100_1;
      patterns[56292] = 25'b11011011_11100010_10111101_1;
      patterns[56293] = 25'b11011011_11100011_10111110_1;
      patterns[56294] = 25'b11011011_11100100_10111111_1;
      patterns[56295] = 25'b11011011_11100101_11000000_1;
      patterns[56296] = 25'b11011011_11100110_11000001_1;
      patterns[56297] = 25'b11011011_11100111_11000010_1;
      patterns[56298] = 25'b11011011_11101000_11000011_1;
      patterns[56299] = 25'b11011011_11101001_11000100_1;
      patterns[56300] = 25'b11011011_11101010_11000101_1;
      patterns[56301] = 25'b11011011_11101011_11000110_1;
      patterns[56302] = 25'b11011011_11101100_11000111_1;
      patterns[56303] = 25'b11011011_11101101_11001000_1;
      patterns[56304] = 25'b11011011_11101110_11001001_1;
      patterns[56305] = 25'b11011011_11101111_11001010_1;
      patterns[56306] = 25'b11011011_11110000_11001011_1;
      patterns[56307] = 25'b11011011_11110001_11001100_1;
      patterns[56308] = 25'b11011011_11110010_11001101_1;
      patterns[56309] = 25'b11011011_11110011_11001110_1;
      patterns[56310] = 25'b11011011_11110100_11001111_1;
      patterns[56311] = 25'b11011011_11110101_11010000_1;
      patterns[56312] = 25'b11011011_11110110_11010001_1;
      patterns[56313] = 25'b11011011_11110111_11010010_1;
      patterns[56314] = 25'b11011011_11111000_11010011_1;
      patterns[56315] = 25'b11011011_11111001_11010100_1;
      patterns[56316] = 25'b11011011_11111010_11010101_1;
      patterns[56317] = 25'b11011011_11111011_11010110_1;
      patterns[56318] = 25'b11011011_11111100_11010111_1;
      patterns[56319] = 25'b11011011_11111101_11011000_1;
      patterns[56320] = 25'b11011011_11111110_11011001_1;
      patterns[56321] = 25'b11011011_11111111_11011010_1;
      patterns[56322] = 25'b11011100_00000000_11011100_0;
      patterns[56323] = 25'b11011100_00000001_11011101_0;
      patterns[56324] = 25'b11011100_00000010_11011110_0;
      patterns[56325] = 25'b11011100_00000011_11011111_0;
      patterns[56326] = 25'b11011100_00000100_11100000_0;
      patterns[56327] = 25'b11011100_00000101_11100001_0;
      patterns[56328] = 25'b11011100_00000110_11100010_0;
      patterns[56329] = 25'b11011100_00000111_11100011_0;
      patterns[56330] = 25'b11011100_00001000_11100100_0;
      patterns[56331] = 25'b11011100_00001001_11100101_0;
      patterns[56332] = 25'b11011100_00001010_11100110_0;
      patterns[56333] = 25'b11011100_00001011_11100111_0;
      patterns[56334] = 25'b11011100_00001100_11101000_0;
      patterns[56335] = 25'b11011100_00001101_11101001_0;
      patterns[56336] = 25'b11011100_00001110_11101010_0;
      patterns[56337] = 25'b11011100_00001111_11101011_0;
      patterns[56338] = 25'b11011100_00010000_11101100_0;
      patterns[56339] = 25'b11011100_00010001_11101101_0;
      patterns[56340] = 25'b11011100_00010010_11101110_0;
      patterns[56341] = 25'b11011100_00010011_11101111_0;
      patterns[56342] = 25'b11011100_00010100_11110000_0;
      patterns[56343] = 25'b11011100_00010101_11110001_0;
      patterns[56344] = 25'b11011100_00010110_11110010_0;
      patterns[56345] = 25'b11011100_00010111_11110011_0;
      patterns[56346] = 25'b11011100_00011000_11110100_0;
      patterns[56347] = 25'b11011100_00011001_11110101_0;
      patterns[56348] = 25'b11011100_00011010_11110110_0;
      patterns[56349] = 25'b11011100_00011011_11110111_0;
      patterns[56350] = 25'b11011100_00011100_11111000_0;
      patterns[56351] = 25'b11011100_00011101_11111001_0;
      patterns[56352] = 25'b11011100_00011110_11111010_0;
      patterns[56353] = 25'b11011100_00011111_11111011_0;
      patterns[56354] = 25'b11011100_00100000_11111100_0;
      patterns[56355] = 25'b11011100_00100001_11111101_0;
      patterns[56356] = 25'b11011100_00100010_11111110_0;
      patterns[56357] = 25'b11011100_00100011_11111111_0;
      patterns[56358] = 25'b11011100_00100100_00000000_1;
      patterns[56359] = 25'b11011100_00100101_00000001_1;
      patterns[56360] = 25'b11011100_00100110_00000010_1;
      patterns[56361] = 25'b11011100_00100111_00000011_1;
      patterns[56362] = 25'b11011100_00101000_00000100_1;
      patterns[56363] = 25'b11011100_00101001_00000101_1;
      patterns[56364] = 25'b11011100_00101010_00000110_1;
      patterns[56365] = 25'b11011100_00101011_00000111_1;
      patterns[56366] = 25'b11011100_00101100_00001000_1;
      patterns[56367] = 25'b11011100_00101101_00001001_1;
      patterns[56368] = 25'b11011100_00101110_00001010_1;
      patterns[56369] = 25'b11011100_00101111_00001011_1;
      patterns[56370] = 25'b11011100_00110000_00001100_1;
      patterns[56371] = 25'b11011100_00110001_00001101_1;
      patterns[56372] = 25'b11011100_00110010_00001110_1;
      patterns[56373] = 25'b11011100_00110011_00001111_1;
      patterns[56374] = 25'b11011100_00110100_00010000_1;
      patterns[56375] = 25'b11011100_00110101_00010001_1;
      patterns[56376] = 25'b11011100_00110110_00010010_1;
      patterns[56377] = 25'b11011100_00110111_00010011_1;
      patterns[56378] = 25'b11011100_00111000_00010100_1;
      patterns[56379] = 25'b11011100_00111001_00010101_1;
      patterns[56380] = 25'b11011100_00111010_00010110_1;
      patterns[56381] = 25'b11011100_00111011_00010111_1;
      patterns[56382] = 25'b11011100_00111100_00011000_1;
      patterns[56383] = 25'b11011100_00111101_00011001_1;
      patterns[56384] = 25'b11011100_00111110_00011010_1;
      patterns[56385] = 25'b11011100_00111111_00011011_1;
      patterns[56386] = 25'b11011100_01000000_00011100_1;
      patterns[56387] = 25'b11011100_01000001_00011101_1;
      patterns[56388] = 25'b11011100_01000010_00011110_1;
      patterns[56389] = 25'b11011100_01000011_00011111_1;
      patterns[56390] = 25'b11011100_01000100_00100000_1;
      patterns[56391] = 25'b11011100_01000101_00100001_1;
      patterns[56392] = 25'b11011100_01000110_00100010_1;
      patterns[56393] = 25'b11011100_01000111_00100011_1;
      patterns[56394] = 25'b11011100_01001000_00100100_1;
      patterns[56395] = 25'b11011100_01001001_00100101_1;
      patterns[56396] = 25'b11011100_01001010_00100110_1;
      patterns[56397] = 25'b11011100_01001011_00100111_1;
      patterns[56398] = 25'b11011100_01001100_00101000_1;
      patterns[56399] = 25'b11011100_01001101_00101001_1;
      patterns[56400] = 25'b11011100_01001110_00101010_1;
      patterns[56401] = 25'b11011100_01001111_00101011_1;
      patterns[56402] = 25'b11011100_01010000_00101100_1;
      patterns[56403] = 25'b11011100_01010001_00101101_1;
      patterns[56404] = 25'b11011100_01010010_00101110_1;
      patterns[56405] = 25'b11011100_01010011_00101111_1;
      patterns[56406] = 25'b11011100_01010100_00110000_1;
      patterns[56407] = 25'b11011100_01010101_00110001_1;
      patterns[56408] = 25'b11011100_01010110_00110010_1;
      patterns[56409] = 25'b11011100_01010111_00110011_1;
      patterns[56410] = 25'b11011100_01011000_00110100_1;
      patterns[56411] = 25'b11011100_01011001_00110101_1;
      patterns[56412] = 25'b11011100_01011010_00110110_1;
      patterns[56413] = 25'b11011100_01011011_00110111_1;
      patterns[56414] = 25'b11011100_01011100_00111000_1;
      patterns[56415] = 25'b11011100_01011101_00111001_1;
      patterns[56416] = 25'b11011100_01011110_00111010_1;
      patterns[56417] = 25'b11011100_01011111_00111011_1;
      patterns[56418] = 25'b11011100_01100000_00111100_1;
      patterns[56419] = 25'b11011100_01100001_00111101_1;
      patterns[56420] = 25'b11011100_01100010_00111110_1;
      patterns[56421] = 25'b11011100_01100011_00111111_1;
      patterns[56422] = 25'b11011100_01100100_01000000_1;
      patterns[56423] = 25'b11011100_01100101_01000001_1;
      patterns[56424] = 25'b11011100_01100110_01000010_1;
      patterns[56425] = 25'b11011100_01100111_01000011_1;
      patterns[56426] = 25'b11011100_01101000_01000100_1;
      patterns[56427] = 25'b11011100_01101001_01000101_1;
      patterns[56428] = 25'b11011100_01101010_01000110_1;
      patterns[56429] = 25'b11011100_01101011_01000111_1;
      patterns[56430] = 25'b11011100_01101100_01001000_1;
      patterns[56431] = 25'b11011100_01101101_01001001_1;
      patterns[56432] = 25'b11011100_01101110_01001010_1;
      patterns[56433] = 25'b11011100_01101111_01001011_1;
      patterns[56434] = 25'b11011100_01110000_01001100_1;
      patterns[56435] = 25'b11011100_01110001_01001101_1;
      patterns[56436] = 25'b11011100_01110010_01001110_1;
      patterns[56437] = 25'b11011100_01110011_01001111_1;
      patterns[56438] = 25'b11011100_01110100_01010000_1;
      patterns[56439] = 25'b11011100_01110101_01010001_1;
      patterns[56440] = 25'b11011100_01110110_01010010_1;
      patterns[56441] = 25'b11011100_01110111_01010011_1;
      patterns[56442] = 25'b11011100_01111000_01010100_1;
      patterns[56443] = 25'b11011100_01111001_01010101_1;
      patterns[56444] = 25'b11011100_01111010_01010110_1;
      patterns[56445] = 25'b11011100_01111011_01010111_1;
      patterns[56446] = 25'b11011100_01111100_01011000_1;
      patterns[56447] = 25'b11011100_01111101_01011001_1;
      patterns[56448] = 25'b11011100_01111110_01011010_1;
      patterns[56449] = 25'b11011100_01111111_01011011_1;
      patterns[56450] = 25'b11011100_10000000_01011100_1;
      patterns[56451] = 25'b11011100_10000001_01011101_1;
      patterns[56452] = 25'b11011100_10000010_01011110_1;
      patterns[56453] = 25'b11011100_10000011_01011111_1;
      patterns[56454] = 25'b11011100_10000100_01100000_1;
      patterns[56455] = 25'b11011100_10000101_01100001_1;
      patterns[56456] = 25'b11011100_10000110_01100010_1;
      patterns[56457] = 25'b11011100_10000111_01100011_1;
      patterns[56458] = 25'b11011100_10001000_01100100_1;
      patterns[56459] = 25'b11011100_10001001_01100101_1;
      patterns[56460] = 25'b11011100_10001010_01100110_1;
      patterns[56461] = 25'b11011100_10001011_01100111_1;
      patterns[56462] = 25'b11011100_10001100_01101000_1;
      patterns[56463] = 25'b11011100_10001101_01101001_1;
      patterns[56464] = 25'b11011100_10001110_01101010_1;
      patterns[56465] = 25'b11011100_10001111_01101011_1;
      patterns[56466] = 25'b11011100_10010000_01101100_1;
      patterns[56467] = 25'b11011100_10010001_01101101_1;
      patterns[56468] = 25'b11011100_10010010_01101110_1;
      patterns[56469] = 25'b11011100_10010011_01101111_1;
      patterns[56470] = 25'b11011100_10010100_01110000_1;
      patterns[56471] = 25'b11011100_10010101_01110001_1;
      patterns[56472] = 25'b11011100_10010110_01110010_1;
      patterns[56473] = 25'b11011100_10010111_01110011_1;
      patterns[56474] = 25'b11011100_10011000_01110100_1;
      patterns[56475] = 25'b11011100_10011001_01110101_1;
      patterns[56476] = 25'b11011100_10011010_01110110_1;
      patterns[56477] = 25'b11011100_10011011_01110111_1;
      patterns[56478] = 25'b11011100_10011100_01111000_1;
      patterns[56479] = 25'b11011100_10011101_01111001_1;
      patterns[56480] = 25'b11011100_10011110_01111010_1;
      patterns[56481] = 25'b11011100_10011111_01111011_1;
      patterns[56482] = 25'b11011100_10100000_01111100_1;
      patterns[56483] = 25'b11011100_10100001_01111101_1;
      patterns[56484] = 25'b11011100_10100010_01111110_1;
      patterns[56485] = 25'b11011100_10100011_01111111_1;
      patterns[56486] = 25'b11011100_10100100_10000000_1;
      patterns[56487] = 25'b11011100_10100101_10000001_1;
      patterns[56488] = 25'b11011100_10100110_10000010_1;
      patterns[56489] = 25'b11011100_10100111_10000011_1;
      patterns[56490] = 25'b11011100_10101000_10000100_1;
      patterns[56491] = 25'b11011100_10101001_10000101_1;
      patterns[56492] = 25'b11011100_10101010_10000110_1;
      patterns[56493] = 25'b11011100_10101011_10000111_1;
      patterns[56494] = 25'b11011100_10101100_10001000_1;
      patterns[56495] = 25'b11011100_10101101_10001001_1;
      patterns[56496] = 25'b11011100_10101110_10001010_1;
      patterns[56497] = 25'b11011100_10101111_10001011_1;
      patterns[56498] = 25'b11011100_10110000_10001100_1;
      patterns[56499] = 25'b11011100_10110001_10001101_1;
      patterns[56500] = 25'b11011100_10110010_10001110_1;
      patterns[56501] = 25'b11011100_10110011_10001111_1;
      patterns[56502] = 25'b11011100_10110100_10010000_1;
      patterns[56503] = 25'b11011100_10110101_10010001_1;
      patterns[56504] = 25'b11011100_10110110_10010010_1;
      patterns[56505] = 25'b11011100_10110111_10010011_1;
      patterns[56506] = 25'b11011100_10111000_10010100_1;
      patterns[56507] = 25'b11011100_10111001_10010101_1;
      patterns[56508] = 25'b11011100_10111010_10010110_1;
      patterns[56509] = 25'b11011100_10111011_10010111_1;
      patterns[56510] = 25'b11011100_10111100_10011000_1;
      patterns[56511] = 25'b11011100_10111101_10011001_1;
      patterns[56512] = 25'b11011100_10111110_10011010_1;
      patterns[56513] = 25'b11011100_10111111_10011011_1;
      patterns[56514] = 25'b11011100_11000000_10011100_1;
      patterns[56515] = 25'b11011100_11000001_10011101_1;
      patterns[56516] = 25'b11011100_11000010_10011110_1;
      patterns[56517] = 25'b11011100_11000011_10011111_1;
      patterns[56518] = 25'b11011100_11000100_10100000_1;
      patterns[56519] = 25'b11011100_11000101_10100001_1;
      patterns[56520] = 25'b11011100_11000110_10100010_1;
      patterns[56521] = 25'b11011100_11000111_10100011_1;
      patterns[56522] = 25'b11011100_11001000_10100100_1;
      patterns[56523] = 25'b11011100_11001001_10100101_1;
      patterns[56524] = 25'b11011100_11001010_10100110_1;
      patterns[56525] = 25'b11011100_11001011_10100111_1;
      patterns[56526] = 25'b11011100_11001100_10101000_1;
      patterns[56527] = 25'b11011100_11001101_10101001_1;
      patterns[56528] = 25'b11011100_11001110_10101010_1;
      patterns[56529] = 25'b11011100_11001111_10101011_1;
      patterns[56530] = 25'b11011100_11010000_10101100_1;
      patterns[56531] = 25'b11011100_11010001_10101101_1;
      patterns[56532] = 25'b11011100_11010010_10101110_1;
      patterns[56533] = 25'b11011100_11010011_10101111_1;
      patterns[56534] = 25'b11011100_11010100_10110000_1;
      patterns[56535] = 25'b11011100_11010101_10110001_1;
      patterns[56536] = 25'b11011100_11010110_10110010_1;
      patterns[56537] = 25'b11011100_11010111_10110011_1;
      patterns[56538] = 25'b11011100_11011000_10110100_1;
      patterns[56539] = 25'b11011100_11011001_10110101_1;
      patterns[56540] = 25'b11011100_11011010_10110110_1;
      patterns[56541] = 25'b11011100_11011011_10110111_1;
      patterns[56542] = 25'b11011100_11011100_10111000_1;
      patterns[56543] = 25'b11011100_11011101_10111001_1;
      patterns[56544] = 25'b11011100_11011110_10111010_1;
      patterns[56545] = 25'b11011100_11011111_10111011_1;
      patterns[56546] = 25'b11011100_11100000_10111100_1;
      patterns[56547] = 25'b11011100_11100001_10111101_1;
      patterns[56548] = 25'b11011100_11100010_10111110_1;
      patterns[56549] = 25'b11011100_11100011_10111111_1;
      patterns[56550] = 25'b11011100_11100100_11000000_1;
      patterns[56551] = 25'b11011100_11100101_11000001_1;
      patterns[56552] = 25'b11011100_11100110_11000010_1;
      patterns[56553] = 25'b11011100_11100111_11000011_1;
      patterns[56554] = 25'b11011100_11101000_11000100_1;
      patterns[56555] = 25'b11011100_11101001_11000101_1;
      patterns[56556] = 25'b11011100_11101010_11000110_1;
      patterns[56557] = 25'b11011100_11101011_11000111_1;
      patterns[56558] = 25'b11011100_11101100_11001000_1;
      patterns[56559] = 25'b11011100_11101101_11001001_1;
      patterns[56560] = 25'b11011100_11101110_11001010_1;
      patterns[56561] = 25'b11011100_11101111_11001011_1;
      patterns[56562] = 25'b11011100_11110000_11001100_1;
      patterns[56563] = 25'b11011100_11110001_11001101_1;
      patterns[56564] = 25'b11011100_11110010_11001110_1;
      patterns[56565] = 25'b11011100_11110011_11001111_1;
      patterns[56566] = 25'b11011100_11110100_11010000_1;
      patterns[56567] = 25'b11011100_11110101_11010001_1;
      patterns[56568] = 25'b11011100_11110110_11010010_1;
      patterns[56569] = 25'b11011100_11110111_11010011_1;
      patterns[56570] = 25'b11011100_11111000_11010100_1;
      patterns[56571] = 25'b11011100_11111001_11010101_1;
      patterns[56572] = 25'b11011100_11111010_11010110_1;
      patterns[56573] = 25'b11011100_11111011_11010111_1;
      patterns[56574] = 25'b11011100_11111100_11011000_1;
      patterns[56575] = 25'b11011100_11111101_11011001_1;
      patterns[56576] = 25'b11011100_11111110_11011010_1;
      patterns[56577] = 25'b11011100_11111111_11011011_1;
      patterns[56578] = 25'b11011101_00000000_11011101_0;
      patterns[56579] = 25'b11011101_00000001_11011110_0;
      patterns[56580] = 25'b11011101_00000010_11011111_0;
      patterns[56581] = 25'b11011101_00000011_11100000_0;
      patterns[56582] = 25'b11011101_00000100_11100001_0;
      patterns[56583] = 25'b11011101_00000101_11100010_0;
      patterns[56584] = 25'b11011101_00000110_11100011_0;
      patterns[56585] = 25'b11011101_00000111_11100100_0;
      patterns[56586] = 25'b11011101_00001000_11100101_0;
      patterns[56587] = 25'b11011101_00001001_11100110_0;
      patterns[56588] = 25'b11011101_00001010_11100111_0;
      patterns[56589] = 25'b11011101_00001011_11101000_0;
      patterns[56590] = 25'b11011101_00001100_11101001_0;
      patterns[56591] = 25'b11011101_00001101_11101010_0;
      patterns[56592] = 25'b11011101_00001110_11101011_0;
      patterns[56593] = 25'b11011101_00001111_11101100_0;
      patterns[56594] = 25'b11011101_00010000_11101101_0;
      patterns[56595] = 25'b11011101_00010001_11101110_0;
      patterns[56596] = 25'b11011101_00010010_11101111_0;
      patterns[56597] = 25'b11011101_00010011_11110000_0;
      patterns[56598] = 25'b11011101_00010100_11110001_0;
      patterns[56599] = 25'b11011101_00010101_11110010_0;
      patterns[56600] = 25'b11011101_00010110_11110011_0;
      patterns[56601] = 25'b11011101_00010111_11110100_0;
      patterns[56602] = 25'b11011101_00011000_11110101_0;
      patterns[56603] = 25'b11011101_00011001_11110110_0;
      patterns[56604] = 25'b11011101_00011010_11110111_0;
      patterns[56605] = 25'b11011101_00011011_11111000_0;
      patterns[56606] = 25'b11011101_00011100_11111001_0;
      patterns[56607] = 25'b11011101_00011101_11111010_0;
      patterns[56608] = 25'b11011101_00011110_11111011_0;
      patterns[56609] = 25'b11011101_00011111_11111100_0;
      patterns[56610] = 25'b11011101_00100000_11111101_0;
      patterns[56611] = 25'b11011101_00100001_11111110_0;
      patterns[56612] = 25'b11011101_00100010_11111111_0;
      patterns[56613] = 25'b11011101_00100011_00000000_1;
      patterns[56614] = 25'b11011101_00100100_00000001_1;
      patterns[56615] = 25'b11011101_00100101_00000010_1;
      patterns[56616] = 25'b11011101_00100110_00000011_1;
      patterns[56617] = 25'b11011101_00100111_00000100_1;
      patterns[56618] = 25'b11011101_00101000_00000101_1;
      patterns[56619] = 25'b11011101_00101001_00000110_1;
      patterns[56620] = 25'b11011101_00101010_00000111_1;
      patterns[56621] = 25'b11011101_00101011_00001000_1;
      patterns[56622] = 25'b11011101_00101100_00001001_1;
      patterns[56623] = 25'b11011101_00101101_00001010_1;
      patterns[56624] = 25'b11011101_00101110_00001011_1;
      patterns[56625] = 25'b11011101_00101111_00001100_1;
      patterns[56626] = 25'b11011101_00110000_00001101_1;
      patterns[56627] = 25'b11011101_00110001_00001110_1;
      patterns[56628] = 25'b11011101_00110010_00001111_1;
      patterns[56629] = 25'b11011101_00110011_00010000_1;
      patterns[56630] = 25'b11011101_00110100_00010001_1;
      patterns[56631] = 25'b11011101_00110101_00010010_1;
      patterns[56632] = 25'b11011101_00110110_00010011_1;
      patterns[56633] = 25'b11011101_00110111_00010100_1;
      patterns[56634] = 25'b11011101_00111000_00010101_1;
      patterns[56635] = 25'b11011101_00111001_00010110_1;
      patterns[56636] = 25'b11011101_00111010_00010111_1;
      patterns[56637] = 25'b11011101_00111011_00011000_1;
      patterns[56638] = 25'b11011101_00111100_00011001_1;
      patterns[56639] = 25'b11011101_00111101_00011010_1;
      patterns[56640] = 25'b11011101_00111110_00011011_1;
      patterns[56641] = 25'b11011101_00111111_00011100_1;
      patterns[56642] = 25'b11011101_01000000_00011101_1;
      patterns[56643] = 25'b11011101_01000001_00011110_1;
      patterns[56644] = 25'b11011101_01000010_00011111_1;
      patterns[56645] = 25'b11011101_01000011_00100000_1;
      patterns[56646] = 25'b11011101_01000100_00100001_1;
      patterns[56647] = 25'b11011101_01000101_00100010_1;
      patterns[56648] = 25'b11011101_01000110_00100011_1;
      patterns[56649] = 25'b11011101_01000111_00100100_1;
      patterns[56650] = 25'b11011101_01001000_00100101_1;
      patterns[56651] = 25'b11011101_01001001_00100110_1;
      patterns[56652] = 25'b11011101_01001010_00100111_1;
      patterns[56653] = 25'b11011101_01001011_00101000_1;
      patterns[56654] = 25'b11011101_01001100_00101001_1;
      patterns[56655] = 25'b11011101_01001101_00101010_1;
      patterns[56656] = 25'b11011101_01001110_00101011_1;
      patterns[56657] = 25'b11011101_01001111_00101100_1;
      patterns[56658] = 25'b11011101_01010000_00101101_1;
      patterns[56659] = 25'b11011101_01010001_00101110_1;
      patterns[56660] = 25'b11011101_01010010_00101111_1;
      patterns[56661] = 25'b11011101_01010011_00110000_1;
      patterns[56662] = 25'b11011101_01010100_00110001_1;
      patterns[56663] = 25'b11011101_01010101_00110010_1;
      patterns[56664] = 25'b11011101_01010110_00110011_1;
      patterns[56665] = 25'b11011101_01010111_00110100_1;
      patterns[56666] = 25'b11011101_01011000_00110101_1;
      patterns[56667] = 25'b11011101_01011001_00110110_1;
      patterns[56668] = 25'b11011101_01011010_00110111_1;
      patterns[56669] = 25'b11011101_01011011_00111000_1;
      patterns[56670] = 25'b11011101_01011100_00111001_1;
      patterns[56671] = 25'b11011101_01011101_00111010_1;
      patterns[56672] = 25'b11011101_01011110_00111011_1;
      patterns[56673] = 25'b11011101_01011111_00111100_1;
      patterns[56674] = 25'b11011101_01100000_00111101_1;
      patterns[56675] = 25'b11011101_01100001_00111110_1;
      patterns[56676] = 25'b11011101_01100010_00111111_1;
      patterns[56677] = 25'b11011101_01100011_01000000_1;
      patterns[56678] = 25'b11011101_01100100_01000001_1;
      patterns[56679] = 25'b11011101_01100101_01000010_1;
      patterns[56680] = 25'b11011101_01100110_01000011_1;
      patterns[56681] = 25'b11011101_01100111_01000100_1;
      patterns[56682] = 25'b11011101_01101000_01000101_1;
      patterns[56683] = 25'b11011101_01101001_01000110_1;
      patterns[56684] = 25'b11011101_01101010_01000111_1;
      patterns[56685] = 25'b11011101_01101011_01001000_1;
      patterns[56686] = 25'b11011101_01101100_01001001_1;
      patterns[56687] = 25'b11011101_01101101_01001010_1;
      patterns[56688] = 25'b11011101_01101110_01001011_1;
      patterns[56689] = 25'b11011101_01101111_01001100_1;
      patterns[56690] = 25'b11011101_01110000_01001101_1;
      patterns[56691] = 25'b11011101_01110001_01001110_1;
      patterns[56692] = 25'b11011101_01110010_01001111_1;
      patterns[56693] = 25'b11011101_01110011_01010000_1;
      patterns[56694] = 25'b11011101_01110100_01010001_1;
      patterns[56695] = 25'b11011101_01110101_01010010_1;
      patterns[56696] = 25'b11011101_01110110_01010011_1;
      patterns[56697] = 25'b11011101_01110111_01010100_1;
      patterns[56698] = 25'b11011101_01111000_01010101_1;
      patterns[56699] = 25'b11011101_01111001_01010110_1;
      patterns[56700] = 25'b11011101_01111010_01010111_1;
      patterns[56701] = 25'b11011101_01111011_01011000_1;
      patterns[56702] = 25'b11011101_01111100_01011001_1;
      patterns[56703] = 25'b11011101_01111101_01011010_1;
      patterns[56704] = 25'b11011101_01111110_01011011_1;
      patterns[56705] = 25'b11011101_01111111_01011100_1;
      patterns[56706] = 25'b11011101_10000000_01011101_1;
      patterns[56707] = 25'b11011101_10000001_01011110_1;
      patterns[56708] = 25'b11011101_10000010_01011111_1;
      patterns[56709] = 25'b11011101_10000011_01100000_1;
      patterns[56710] = 25'b11011101_10000100_01100001_1;
      patterns[56711] = 25'b11011101_10000101_01100010_1;
      patterns[56712] = 25'b11011101_10000110_01100011_1;
      patterns[56713] = 25'b11011101_10000111_01100100_1;
      patterns[56714] = 25'b11011101_10001000_01100101_1;
      patterns[56715] = 25'b11011101_10001001_01100110_1;
      patterns[56716] = 25'b11011101_10001010_01100111_1;
      patterns[56717] = 25'b11011101_10001011_01101000_1;
      patterns[56718] = 25'b11011101_10001100_01101001_1;
      patterns[56719] = 25'b11011101_10001101_01101010_1;
      patterns[56720] = 25'b11011101_10001110_01101011_1;
      patterns[56721] = 25'b11011101_10001111_01101100_1;
      patterns[56722] = 25'b11011101_10010000_01101101_1;
      patterns[56723] = 25'b11011101_10010001_01101110_1;
      patterns[56724] = 25'b11011101_10010010_01101111_1;
      patterns[56725] = 25'b11011101_10010011_01110000_1;
      patterns[56726] = 25'b11011101_10010100_01110001_1;
      patterns[56727] = 25'b11011101_10010101_01110010_1;
      patterns[56728] = 25'b11011101_10010110_01110011_1;
      patterns[56729] = 25'b11011101_10010111_01110100_1;
      patterns[56730] = 25'b11011101_10011000_01110101_1;
      patterns[56731] = 25'b11011101_10011001_01110110_1;
      patterns[56732] = 25'b11011101_10011010_01110111_1;
      patterns[56733] = 25'b11011101_10011011_01111000_1;
      patterns[56734] = 25'b11011101_10011100_01111001_1;
      patterns[56735] = 25'b11011101_10011101_01111010_1;
      patterns[56736] = 25'b11011101_10011110_01111011_1;
      patterns[56737] = 25'b11011101_10011111_01111100_1;
      patterns[56738] = 25'b11011101_10100000_01111101_1;
      patterns[56739] = 25'b11011101_10100001_01111110_1;
      patterns[56740] = 25'b11011101_10100010_01111111_1;
      patterns[56741] = 25'b11011101_10100011_10000000_1;
      patterns[56742] = 25'b11011101_10100100_10000001_1;
      patterns[56743] = 25'b11011101_10100101_10000010_1;
      patterns[56744] = 25'b11011101_10100110_10000011_1;
      patterns[56745] = 25'b11011101_10100111_10000100_1;
      patterns[56746] = 25'b11011101_10101000_10000101_1;
      patterns[56747] = 25'b11011101_10101001_10000110_1;
      patterns[56748] = 25'b11011101_10101010_10000111_1;
      patterns[56749] = 25'b11011101_10101011_10001000_1;
      patterns[56750] = 25'b11011101_10101100_10001001_1;
      patterns[56751] = 25'b11011101_10101101_10001010_1;
      patterns[56752] = 25'b11011101_10101110_10001011_1;
      patterns[56753] = 25'b11011101_10101111_10001100_1;
      patterns[56754] = 25'b11011101_10110000_10001101_1;
      patterns[56755] = 25'b11011101_10110001_10001110_1;
      patterns[56756] = 25'b11011101_10110010_10001111_1;
      patterns[56757] = 25'b11011101_10110011_10010000_1;
      patterns[56758] = 25'b11011101_10110100_10010001_1;
      patterns[56759] = 25'b11011101_10110101_10010010_1;
      patterns[56760] = 25'b11011101_10110110_10010011_1;
      patterns[56761] = 25'b11011101_10110111_10010100_1;
      patterns[56762] = 25'b11011101_10111000_10010101_1;
      patterns[56763] = 25'b11011101_10111001_10010110_1;
      patterns[56764] = 25'b11011101_10111010_10010111_1;
      patterns[56765] = 25'b11011101_10111011_10011000_1;
      patterns[56766] = 25'b11011101_10111100_10011001_1;
      patterns[56767] = 25'b11011101_10111101_10011010_1;
      patterns[56768] = 25'b11011101_10111110_10011011_1;
      patterns[56769] = 25'b11011101_10111111_10011100_1;
      patterns[56770] = 25'b11011101_11000000_10011101_1;
      patterns[56771] = 25'b11011101_11000001_10011110_1;
      patterns[56772] = 25'b11011101_11000010_10011111_1;
      patterns[56773] = 25'b11011101_11000011_10100000_1;
      patterns[56774] = 25'b11011101_11000100_10100001_1;
      patterns[56775] = 25'b11011101_11000101_10100010_1;
      patterns[56776] = 25'b11011101_11000110_10100011_1;
      patterns[56777] = 25'b11011101_11000111_10100100_1;
      patterns[56778] = 25'b11011101_11001000_10100101_1;
      patterns[56779] = 25'b11011101_11001001_10100110_1;
      patterns[56780] = 25'b11011101_11001010_10100111_1;
      patterns[56781] = 25'b11011101_11001011_10101000_1;
      patterns[56782] = 25'b11011101_11001100_10101001_1;
      patterns[56783] = 25'b11011101_11001101_10101010_1;
      patterns[56784] = 25'b11011101_11001110_10101011_1;
      patterns[56785] = 25'b11011101_11001111_10101100_1;
      patterns[56786] = 25'b11011101_11010000_10101101_1;
      patterns[56787] = 25'b11011101_11010001_10101110_1;
      patterns[56788] = 25'b11011101_11010010_10101111_1;
      patterns[56789] = 25'b11011101_11010011_10110000_1;
      patterns[56790] = 25'b11011101_11010100_10110001_1;
      patterns[56791] = 25'b11011101_11010101_10110010_1;
      patterns[56792] = 25'b11011101_11010110_10110011_1;
      patterns[56793] = 25'b11011101_11010111_10110100_1;
      patterns[56794] = 25'b11011101_11011000_10110101_1;
      patterns[56795] = 25'b11011101_11011001_10110110_1;
      patterns[56796] = 25'b11011101_11011010_10110111_1;
      patterns[56797] = 25'b11011101_11011011_10111000_1;
      patterns[56798] = 25'b11011101_11011100_10111001_1;
      patterns[56799] = 25'b11011101_11011101_10111010_1;
      patterns[56800] = 25'b11011101_11011110_10111011_1;
      patterns[56801] = 25'b11011101_11011111_10111100_1;
      patterns[56802] = 25'b11011101_11100000_10111101_1;
      patterns[56803] = 25'b11011101_11100001_10111110_1;
      patterns[56804] = 25'b11011101_11100010_10111111_1;
      patterns[56805] = 25'b11011101_11100011_11000000_1;
      patterns[56806] = 25'b11011101_11100100_11000001_1;
      patterns[56807] = 25'b11011101_11100101_11000010_1;
      patterns[56808] = 25'b11011101_11100110_11000011_1;
      patterns[56809] = 25'b11011101_11100111_11000100_1;
      patterns[56810] = 25'b11011101_11101000_11000101_1;
      patterns[56811] = 25'b11011101_11101001_11000110_1;
      patterns[56812] = 25'b11011101_11101010_11000111_1;
      patterns[56813] = 25'b11011101_11101011_11001000_1;
      patterns[56814] = 25'b11011101_11101100_11001001_1;
      patterns[56815] = 25'b11011101_11101101_11001010_1;
      patterns[56816] = 25'b11011101_11101110_11001011_1;
      patterns[56817] = 25'b11011101_11101111_11001100_1;
      patterns[56818] = 25'b11011101_11110000_11001101_1;
      patterns[56819] = 25'b11011101_11110001_11001110_1;
      patterns[56820] = 25'b11011101_11110010_11001111_1;
      patterns[56821] = 25'b11011101_11110011_11010000_1;
      patterns[56822] = 25'b11011101_11110100_11010001_1;
      patterns[56823] = 25'b11011101_11110101_11010010_1;
      patterns[56824] = 25'b11011101_11110110_11010011_1;
      patterns[56825] = 25'b11011101_11110111_11010100_1;
      patterns[56826] = 25'b11011101_11111000_11010101_1;
      patterns[56827] = 25'b11011101_11111001_11010110_1;
      patterns[56828] = 25'b11011101_11111010_11010111_1;
      patterns[56829] = 25'b11011101_11111011_11011000_1;
      patterns[56830] = 25'b11011101_11111100_11011001_1;
      patterns[56831] = 25'b11011101_11111101_11011010_1;
      patterns[56832] = 25'b11011101_11111110_11011011_1;
      patterns[56833] = 25'b11011101_11111111_11011100_1;
      patterns[56834] = 25'b11011110_00000000_11011110_0;
      patterns[56835] = 25'b11011110_00000001_11011111_0;
      patterns[56836] = 25'b11011110_00000010_11100000_0;
      patterns[56837] = 25'b11011110_00000011_11100001_0;
      patterns[56838] = 25'b11011110_00000100_11100010_0;
      patterns[56839] = 25'b11011110_00000101_11100011_0;
      patterns[56840] = 25'b11011110_00000110_11100100_0;
      patterns[56841] = 25'b11011110_00000111_11100101_0;
      patterns[56842] = 25'b11011110_00001000_11100110_0;
      patterns[56843] = 25'b11011110_00001001_11100111_0;
      patterns[56844] = 25'b11011110_00001010_11101000_0;
      patterns[56845] = 25'b11011110_00001011_11101001_0;
      patterns[56846] = 25'b11011110_00001100_11101010_0;
      patterns[56847] = 25'b11011110_00001101_11101011_0;
      patterns[56848] = 25'b11011110_00001110_11101100_0;
      patterns[56849] = 25'b11011110_00001111_11101101_0;
      patterns[56850] = 25'b11011110_00010000_11101110_0;
      patterns[56851] = 25'b11011110_00010001_11101111_0;
      patterns[56852] = 25'b11011110_00010010_11110000_0;
      patterns[56853] = 25'b11011110_00010011_11110001_0;
      patterns[56854] = 25'b11011110_00010100_11110010_0;
      patterns[56855] = 25'b11011110_00010101_11110011_0;
      patterns[56856] = 25'b11011110_00010110_11110100_0;
      patterns[56857] = 25'b11011110_00010111_11110101_0;
      patterns[56858] = 25'b11011110_00011000_11110110_0;
      patterns[56859] = 25'b11011110_00011001_11110111_0;
      patterns[56860] = 25'b11011110_00011010_11111000_0;
      patterns[56861] = 25'b11011110_00011011_11111001_0;
      patterns[56862] = 25'b11011110_00011100_11111010_0;
      patterns[56863] = 25'b11011110_00011101_11111011_0;
      patterns[56864] = 25'b11011110_00011110_11111100_0;
      patterns[56865] = 25'b11011110_00011111_11111101_0;
      patterns[56866] = 25'b11011110_00100000_11111110_0;
      patterns[56867] = 25'b11011110_00100001_11111111_0;
      patterns[56868] = 25'b11011110_00100010_00000000_1;
      patterns[56869] = 25'b11011110_00100011_00000001_1;
      patterns[56870] = 25'b11011110_00100100_00000010_1;
      patterns[56871] = 25'b11011110_00100101_00000011_1;
      patterns[56872] = 25'b11011110_00100110_00000100_1;
      patterns[56873] = 25'b11011110_00100111_00000101_1;
      patterns[56874] = 25'b11011110_00101000_00000110_1;
      patterns[56875] = 25'b11011110_00101001_00000111_1;
      patterns[56876] = 25'b11011110_00101010_00001000_1;
      patterns[56877] = 25'b11011110_00101011_00001001_1;
      patterns[56878] = 25'b11011110_00101100_00001010_1;
      patterns[56879] = 25'b11011110_00101101_00001011_1;
      patterns[56880] = 25'b11011110_00101110_00001100_1;
      patterns[56881] = 25'b11011110_00101111_00001101_1;
      patterns[56882] = 25'b11011110_00110000_00001110_1;
      patterns[56883] = 25'b11011110_00110001_00001111_1;
      patterns[56884] = 25'b11011110_00110010_00010000_1;
      patterns[56885] = 25'b11011110_00110011_00010001_1;
      patterns[56886] = 25'b11011110_00110100_00010010_1;
      patterns[56887] = 25'b11011110_00110101_00010011_1;
      patterns[56888] = 25'b11011110_00110110_00010100_1;
      patterns[56889] = 25'b11011110_00110111_00010101_1;
      patterns[56890] = 25'b11011110_00111000_00010110_1;
      patterns[56891] = 25'b11011110_00111001_00010111_1;
      patterns[56892] = 25'b11011110_00111010_00011000_1;
      patterns[56893] = 25'b11011110_00111011_00011001_1;
      patterns[56894] = 25'b11011110_00111100_00011010_1;
      patterns[56895] = 25'b11011110_00111101_00011011_1;
      patterns[56896] = 25'b11011110_00111110_00011100_1;
      patterns[56897] = 25'b11011110_00111111_00011101_1;
      patterns[56898] = 25'b11011110_01000000_00011110_1;
      patterns[56899] = 25'b11011110_01000001_00011111_1;
      patterns[56900] = 25'b11011110_01000010_00100000_1;
      patterns[56901] = 25'b11011110_01000011_00100001_1;
      patterns[56902] = 25'b11011110_01000100_00100010_1;
      patterns[56903] = 25'b11011110_01000101_00100011_1;
      patterns[56904] = 25'b11011110_01000110_00100100_1;
      patterns[56905] = 25'b11011110_01000111_00100101_1;
      patterns[56906] = 25'b11011110_01001000_00100110_1;
      patterns[56907] = 25'b11011110_01001001_00100111_1;
      patterns[56908] = 25'b11011110_01001010_00101000_1;
      patterns[56909] = 25'b11011110_01001011_00101001_1;
      patterns[56910] = 25'b11011110_01001100_00101010_1;
      patterns[56911] = 25'b11011110_01001101_00101011_1;
      patterns[56912] = 25'b11011110_01001110_00101100_1;
      patterns[56913] = 25'b11011110_01001111_00101101_1;
      patterns[56914] = 25'b11011110_01010000_00101110_1;
      patterns[56915] = 25'b11011110_01010001_00101111_1;
      patterns[56916] = 25'b11011110_01010010_00110000_1;
      patterns[56917] = 25'b11011110_01010011_00110001_1;
      patterns[56918] = 25'b11011110_01010100_00110010_1;
      patterns[56919] = 25'b11011110_01010101_00110011_1;
      patterns[56920] = 25'b11011110_01010110_00110100_1;
      patterns[56921] = 25'b11011110_01010111_00110101_1;
      patterns[56922] = 25'b11011110_01011000_00110110_1;
      patterns[56923] = 25'b11011110_01011001_00110111_1;
      patterns[56924] = 25'b11011110_01011010_00111000_1;
      patterns[56925] = 25'b11011110_01011011_00111001_1;
      patterns[56926] = 25'b11011110_01011100_00111010_1;
      patterns[56927] = 25'b11011110_01011101_00111011_1;
      patterns[56928] = 25'b11011110_01011110_00111100_1;
      patterns[56929] = 25'b11011110_01011111_00111101_1;
      patterns[56930] = 25'b11011110_01100000_00111110_1;
      patterns[56931] = 25'b11011110_01100001_00111111_1;
      patterns[56932] = 25'b11011110_01100010_01000000_1;
      patterns[56933] = 25'b11011110_01100011_01000001_1;
      patterns[56934] = 25'b11011110_01100100_01000010_1;
      patterns[56935] = 25'b11011110_01100101_01000011_1;
      patterns[56936] = 25'b11011110_01100110_01000100_1;
      patterns[56937] = 25'b11011110_01100111_01000101_1;
      patterns[56938] = 25'b11011110_01101000_01000110_1;
      patterns[56939] = 25'b11011110_01101001_01000111_1;
      patterns[56940] = 25'b11011110_01101010_01001000_1;
      patterns[56941] = 25'b11011110_01101011_01001001_1;
      patterns[56942] = 25'b11011110_01101100_01001010_1;
      patterns[56943] = 25'b11011110_01101101_01001011_1;
      patterns[56944] = 25'b11011110_01101110_01001100_1;
      patterns[56945] = 25'b11011110_01101111_01001101_1;
      patterns[56946] = 25'b11011110_01110000_01001110_1;
      patterns[56947] = 25'b11011110_01110001_01001111_1;
      patterns[56948] = 25'b11011110_01110010_01010000_1;
      patterns[56949] = 25'b11011110_01110011_01010001_1;
      patterns[56950] = 25'b11011110_01110100_01010010_1;
      patterns[56951] = 25'b11011110_01110101_01010011_1;
      patterns[56952] = 25'b11011110_01110110_01010100_1;
      patterns[56953] = 25'b11011110_01110111_01010101_1;
      patterns[56954] = 25'b11011110_01111000_01010110_1;
      patterns[56955] = 25'b11011110_01111001_01010111_1;
      patterns[56956] = 25'b11011110_01111010_01011000_1;
      patterns[56957] = 25'b11011110_01111011_01011001_1;
      patterns[56958] = 25'b11011110_01111100_01011010_1;
      patterns[56959] = 25'b11011110_01111101_01011011_1;
      patterns[56960] = 25'b11011110_01111110_01011100_1;
      patterns[56961] = 25'b11011110_01111111_01011101_1;
      patterns[56962] = 25'b11011110_10000000_01011110_1;
      patterns[56963] = 25'b11011110_10000001_01011111_1;
      patterns[56964] = 25'b11011110_10000010_01100000_1;
      patterns[56965] = 25'b11011110_10000011_01100001_1;
      patterns[56966] = 25'b11011110_10000100_01100010_1;
      patterns[56967] = 25'b11011110_10000101_01100011_1;
      patterns[56968] = 25'b11011110_10000110_01100100_1;
      patterns[56969] = 25'b11011110_10000111_01100101_1;
      patterns[56970] = 25'b11011110_10001000_01100110_1;
      patterns[56971] = 25'b11011110_10001001_01100111_1;
      patterns[56972] = 25'b11011110_10001010_01101000_1;
      patterns[56973] = 25'b11011110_10001011_01101001_1;
      patterns[56974] = 25'b11011110_10001100_01101010_1;
      patterns[56975] = 25'b11011110_10001101_01101011_1;
      patterns[56976] = 25'b11011110_10001110_01101100_1;
      patterns[56977] = 25'b11011110_10001111_01101101_1;
      patterns[56978] = 25'b11011110_10010000_01101110_1;
      patterns[56979] = 25'b11011110_10010001_01101111_1;
      patterns[56980] = 25'b11011110_10010010_01110000_1;
      patterns[56981] = 25'b11011110_10010011_01110001_1;
      patterns[56982] = 25'b11011110_10010100_01110010_1;
      patterns[56983] = 25'b11011110_10010101_01110011_1;
      patterns[56984] = 25'b11011110_10010110_01110100_1;
      patterns[56985] = 25'b11011110_10010111_01110101_1;
      patterns[56986] = 25'b11011110_10011000_01110110_1;
      patterns[56987] = 25'b11011110_10011001_01110111_1;
      patterns[56988] = 25'b11011110_10011010_01111000_1;
      patterns[56989] = 25'b11011110_10011011_01111001_1;
      patterns[56990] = 25'b11011110_10011100_01111010_1;
      patterns[56991] = 25'b11011110_10011101_01111011_1;
      patterns[56992] = 25'b11011110_10011110_01111100_1;
      patterns[56993] = 25'b11011110_10011111_01111101_1;
      patterns[56994] = 25'b11011110_10100000_01111110_1;
      patterns[56995] = 25'b11011110_10100001_01111111_1;
      patterns[56996] = 25'b11011110_10100010_10000000_1;
      patterns[56997] = 25'b11011110_10100011_10000001_1;
      patterns[56998] = 25'b11011110_10100100_10000010_1;
      patterns[56999] = 25'b11011110_10100101_10000011_1;
      patterns[57000] = 25'b11011110_10100110_10000100_1;
      patterns[57001] = 25'b11011110_10100111_10000101_1;
      patterns[57002] = 25'b11011110_10101000_10000110_1;
      patterns[57003] = 25'b11011110_10101001_10000111_1;
      patterns[57004] = 25'b11011110_10101010_10001000_1;
      patterns[57005] = 25'b11011110_10101011_10001001_1;
      patterns[57006] = 25'b11011110_10101100_10001010_1;
      patterns[57007] = 25'b11011110_10101101_10001011_1;
      patterns[57008] = 25'b11011110_10101110_10001100_1;
      patterns[57009] = 25'b11011110_10101111_10001101_1;
      patterns[57010] = 25'b11011110_10110000_10001110_1;
      patterns[57011] = 25'b11011110_10110001_10001111_1;
      patterns[57012] = 25'b11011110_10110010_10010000_1;
      patterns[57013] = 25'b11011110_10110011_10010001_1;
      patterns[57014] = 25'b11011110_10110100_10010010_1;
      patterns[57015] = 25'b11011110_10110101_10010011_1;
      patterns[57016] = 25'b11011110_10110110_10010100_1;
      patterns[57017] = 25'b11011110_10110111_10010101_1;
      patterns[57018] = 25'b11011110_10111000_10010110_1;
      patterns[57019] = 25'b11011110_10111001_10010111_1;
      patterns[57020] = 25'b11011110_10111010_10011000_1;
      patterns[57021] = 25'b11011110_10111011_10011001_1;
      patterns[57022] = 25'b11011110_10111100_10011010_1;
      patterns[57023] = 25'b11011110_10111101_10011011_1;
      patterns[57024] = 25'b11011110_10111110_10011100_1;
      patterns[57025] = 25'b11011110_10111111_10011101_1;
      patterns[57026] = 25'b11011110_11000000_10011110_1;
      patterns[57027] = 25'b11011110_11000001_10011111_1;
      patterns[57028] = 25'b11011110_11000010_10100000_1;
      patterns[57029] = 25'b11011110_11000011_10100001_1;
      patterns[57030] = 25'b11011110_11000100_10100010_1;
      patterns[57031] = 25'b11011110_11000101_10100011_1;
      patterns[57032] = 25'b11011110_11000110_10100100_1;
      patterns[57033] = 25'b11011110_11000111_10100101_1;
      patterns[57034] = 25'b11011110_11001000_10100110_1;
      patterns[57035] = 25'b11011110_11001001_10100111_1;
      patterns[57036] = 25'b11011110_11001010_10101000_1;
      patterns[57037] = 25'b11011110_11001011_10101001_1;
      patterns[57038] = 25'b11011110_11001100_10101010_1;
      patterns[57039] = 25'b11011110_11001101_10101011_1;
      patterns[57040] = 25'b11011110_11001110_10101100_1;
      patterns[57041] = 25'b11011110_11001111_10101101_1;
      patterns[57042] = 25'b11011110_11010000_10101110_1;
      patterns[57043] = 25'b11011110_11010001_10101111_1;
      patterns[57044] = 25'b11011110_11010010_10110000_1;
      patterns[57045] = 25'b11011110_11010011_10110001_1;
      patterns[57046] = 25'b11011110_11010100_10110010_1;
      patterns[57047] = 25'b11011110_11010101_10110011_1;
      patterns[57048] = 25'b11011110_11010110_10110100_1;
      patterns[57049] = 25'b11011110_11010111_10110101_1;
      patterns[57050] = 25'b11011110_11011000_10110110_1;
      patterns[57051] = 25'b11011110_11011001_10110111_1;
      patterns[57052] = 25'b11011110_11011010_10111000_1;
      patterns[57053] = 25'b11011110_11011011_10111001_1;
      patterns[57054] = 25'b11011110_11011100_10111010_1;
      patterns[57055] = 25'b11011110_11011101_10111011_1;
      patterns[57056] = 25'b11011110_11011110_10111100_1;
      patterns[57057] = 25'b11011110_11011111_10111101_1;
      patterns[57058] = 25'b11011110_11100000_10111110_1;
      patterns[57059] = 25'b11011110_11100001_10111111_1;
      patterns[57060] = 25'b11011110_11100010_11000000_1;
      patterns[57061] = 25'b11011110_11100011_11000001_1;
      patterns[57062] = 25'b11011110_11100100_11000010_1;
      patterns[57063] = 25'b11011110_11100101_11000011_1;
      patterns[57064] = 25'b11011110_11100110_11000100_1;
      patterns[57065] = 25'b11011110_11100111_11000101_1;
      patterns[57066] = 25'b11011110_11101000_11000110_1;
      patterns[57067] = 25'b11011110_11101001_11000111_1;
      patterns[57068] = 25'b11011110_11101010_11001000_1;
      patterns[57069] = 25'b11011110_11101011_11001001_1;
      patterns[57070] = 25'b11011110_11101100_11001010_1;
      patterns[57071] = 25'b11011110_11101101_11001011_1;
      patterns[57072] = 25'b11011110_11101110_11001100_1;
      patterns[57073] = 25'b11011110_11101111_11001101_1;
      patterns[57074] = 25'b11011110_11110000_11001110_1;
      patterns[57075] = 25'b11011110_11110001_11001111_1;
      patterns[57076] = 25'b11011110_11110010_11010000_1;
      patterns[57077] = 25'b11011110_11110011_11010001_1;
      patterns[57078] = 25'b11011110_11110100_11010010_1;
      patterns[57079] = 25'b11011110_11110101_11010011_1;
      patterns[57080] = 25'b11011110_11110110_11010100_1;
      patterns[57081] = 25'b11011110_11110111_11010101_1;
      patterns[57082] = 25'b11011110_11111000_11010110_1;
      patterns[57083] = 25'b11011110_11111001_11010111_1;
      patterns[57084] = 25'b11011110_11111010_11011000_1;
      patterns[57085] = 25'b11011110_11111011_11011001_1;
      patterns[57086] = 25'b11011110_11111100_11011010_1;
      patterns[57087] = 25'b11011110_11111101_11011011_1;
      patterns[57088] = 25'b11011110_11111110_11011100_1;
      patterns[57089] = 25'b11011110_11111111_11011101_1;
      patterns[57090] = 25'b11011111_00000000_11011111_0;
      patterns[57091] = 25'b11011111_00000001_11100000_0;
      patterns[57092] = 25'b11011111_00000010_11100001_0;
      patterns[57093] = 25'b11011111_00000011_11100010_0;
      patterns[57094] = 25'b11011111_00000100_11100011_0;
      patterns[57095] = 25'b11011111_00000101_11100100_0;
      patterns[57096] = 25'b11011111_00000110_11100101_0;
      patterns[57097] = 25'b11011111_00000111_11100110_0;
      patterns[57098] = 25'b11011111_00001000_11100111_0;
      patterns[57099] = 25'b11011111_00001001_11101000_0;
      patterns[57100] = 25'b11011111_00001010_11101001_0;
      patterns[57101] = 25'b11011111_00001011_11101010_0;
      patterns[57102] = 25'b11011111_00001100_11101011_0;
      patterns[57103] = 25'b11011111_00001101_11101100_0;
      patterns[57104] = 25'b11011111_00001110_11101101_0;
      patterns[57105] = 25'b11011111_00001111_11101110_0;
      patterns[57106] = 25'b11011111_00010000_11101111_0;
      patterns[57107] = 25'b11011111_00010001_11110000_0;
      patterns[57108] = 25'b11011111_00010010_11110001_0;
      patterns[57109] = 25'b11011111_00010011_11110010_0;
      patterns[57110] = 25'b11011111_00010100_11110011_0;
      patterns[57111] = 25'b11011111_00010101_11110100_0;
      patterns[57112] = 25'b11011111_00010110_11110101_0;
      patterns[57113] = 25'b11011111_00010111_11110110_0;
      patterns[57114] = 25'b11011111_00011000_11110111_0;
      patterns[57115] = 25'b11011111_00011001_11111000_0;
      patterns[57116] = 25'b11011111_00011010_11111001_0;
      patterns[57117] = 25'b11011111_00011011_11111010_0;
      patterns[57118] = 25'b11011111_00011100_11111011_0;
      patterns[57119] = 25'b11011111_00011101_11111100_0;
      patterns[57120] = 25'b11011111_00011110_11111101_0;
      patterns[57121] = 25'b11011111_00011111_11111110_0;
      patterns[57122] = 25'b11011111_00100000_11111111_0;
      patterns[57123] = 25'b11011111_00100001_00000000_1;
      patterns[57124] = 25'b11011111_00100010_00000001_1;
      patterns[57125] = 25'b11011111_00100011_00000010_1;
      patterns[57126] = 25'b11011111_00100100_00000011_1;
      patterns[57127] = 25'b11011111_00100101_00000100_1;
      patterns[57128] = 25'b11011111_00100110_00000101_1;
      patterns[57129] = 25'b11011111_00100111_00000110_1;
      patterns[57130] = 25'b11011111_00101000_00000111_1;
      patterns[57131] = 25'b11011111_00101001_00001000_1;
      patterns[57132] = 25'b11011111_00101010_00001001_1;
      patterns[57133] = 25'b11011111_00101011_00001010_1;
      patterns[57134] = 25'b11011111_00101100_00001011_1;
      patterns[57135] = 25'b11011111_00101101_00001100_1;
      patterns[57136] = 25'b11011111_00101110_00001101_1;
      patterns[57137] = 25'b11011111_00101111_00001110_1;
      patterns[57138] = 25'b11011111_00110000_00001111_1;
      patterns[57139] = 25'b11011111_00110001_00010000_1;
      patterns[57140] = 25'b11011111_00110010_00010001_1;
      patterns[57141] = 25'b11011111_00110011_00010010_1;
      patterns[57142] = 25'b11011111_00110100_00010011_1;
      patterns[57143] = 25'b11011111_00110101_00010100_1;
      patterns[57144] = 25'b11011111_00110110_00010101_1;
      patterns[57145] = 25'b11011111_00110111_00010110_1;
      patterns[57146] = 25'b11011111_00111000_00010111_1;
      patterns[57147] = 25'b11011111_00111001_00011000_1;
      patterns[57148] = 25'b11011111_00111010_00011001_1;
      patterns[57149] = 25'b11011111_00111011_00011010_1;
      patterns[57150] = 25'b11011111_00111100_00011011_1;
      patterns[57151] = 25'b11011111_00111101_00011100_1;
      patterns[57152] = 25'b11011111_00111110_00011101_1;
      patterns[57153] = 25'b11011111_00111111_00011110_1;
      patterns[57154] = 25'b11011111_01000000_00011111_1;
      patterns[57155] = 25'b11011111_01000001_00100000_1;
      patterns[57156] = 25'b11011111_01000010_00100001_1;
      patterns[57157] = 25'b11011111_01000011_00100010_1;
      patterns[57158] = 25'b11011111_01000100_00100011_1;
      patterns[57159] = 25'b11011111_01000101_00100100_1;
      patterns[57160] = 25'b11011111_01000110_00100101_1;
      patterns[57161] = 25'b11011111_01000111_00100110_1;
      patterns[57162] = 25'b11011111_01001000_00100111_1;
      patterns[57163] = 25'b11011111_01001001_00101000_1;
      patterns[57164] = 25'b11011111_01001010_00101001_1;
      patterns[57165] = 25'b11011111_01001011_00101010_1;
      patterns[57166] = 25'b11011111_01001100_00101011_1;
      patterns[57167] = 25'b11011111_01001101_00101100_1;
      patterns[57168] = 25'b11011111_01001110_00101101_1;
      patterns[57169] = 25'b11011111_01001111_00101110_1;
      patterns[57170] = 25'b11011111_01010000_00101111_1;
      patterns[57171] = 25'b11011111_01010001_00110000_1;
      patterns[57172] = 25'b11011111_01010010_00110001_1;
      patterns[57173] = 25'b11011111_01010011_00110010_1;
      patterns[57174] = 25'b11011111_01010100_00110011_1;
      patterns[57175] = 25'b11011111_01010101_00110100_1;
      patterns[57176] = 25'b11011111_01010110_00110101_1;
      patterns[57177] = 25'b11011111_01010111_00110110_1;
      patterns[57178] = 25'b11011111_01011000_00110111_1;
      patterns[57179] = 25'b11011111_01011001_00111000_1;
      patterns[57180] = 25'b11011111_01011010_00111001_1;
      patterns[57181] = 25'b11011111_01011011_00111010_1;
      patterns[57182] = 25'b11011111_01011100_00111011_1;
      patterns[57183] = 25'b11011111_01011101_00111100_1;
      patterns[57184] = 25'b11011111_01011110_00111101_1;
      patterns[57185] = 25'b11011111_01011111_00111110_1;
      patterns[57186] = 25'b11011111_01100000_00111111_1;
      patterns[57187] = 25'b11011111_01100001_01000000_1;
      patterns[57188] = 25'b11011111_01100010_01000001_1;
      patterns[57189] = 25'b11011111_01100011_01000010_1;
      patterns[57190] = 25'b11011111_01100100_01000011_1;
      patterns[57191] = 25'b11011111_01100101_01000100_1;
      patterns[57192] = 25'b11011111_01100110_01000101_1;
      patterns[57193] = 25'b11011111_01100111_01000110_1;
      patterns[57194] = 25'b11011111_01101000_01000111_1;
      patterns[57195] = 25'b11011111_01101001_01001000_1;
      patterns[57196] = 25'b11011111_01101010_01001001_1;
      patterns[57197] = 25'b11011111_01101011_01001010_1;
      patterns[57198] = 25'b11011111_01101100_01001011_1;
      patterns[57199] = 25'b11011111_01101101_01001100_1;
      patterns[57200] = 25'b11011111_01101110_01001101_1;
      patterns[57201] = 25'b11011111_01101111_01001110_1;
      patterns[57202] = 25'b11011111_01110000_01001111_1;
      patterns[57203] = 25'b11011111_01110001_01010000_1;
      patterns[57204] = 25'b11011111_01110010_01010001_1;
      patterns[57205] = 25'b11011111_01110011_01010010_1;
      patterns[57206] = 25'b11011111_01110100_01010011_1;
      patterns[57207] = 25'b11011111_01110101_01010100_1;
      patterns[57208] = 25'b11011111_01110110_01010101_1;
      patterns[57209] = 25'b11011111_01110111_01010110_1;
      patterns[57210] = 25'b11011111_01111000_01010111_1;
      patterns[57211] = 25'b11011111_01111001_01011000_1;
      patterns[57212] = 25'b11011111_01111010_01011001_1;
      patterns[57213] = 25'b11011111_01111011_01011010_1;
      patterns[57214] = 25'b11011111_01111100_01011011_1;
      patterns[57215] = 25'b11011111_01111101_01011100_1;
      patterns[57216] = 25'b11011111_01111110_01011101_1;
      patterns[57217] = 25'b11011111_01111111_01011110_1;
      patterns[57218] = 25'b11011111_10000000_01011111_1;
      patterns[57219] = 25'b11011111_10000001_01100000_1;
      patterns[57220] = 25'b11011111_10000010_01100001_1;
      patterns[57221] = 25'b11011111_10000011_01100010_1;
      patterns[57222] = 25'b11011111_10000100_01100011_1;
      patterns[57223] = 25'b11011111_10000101_01100100_1;
      patterns[57224] = 25'b11011111_10000110_01100101_1;
      patterns[57225] = 25'b11011111_10000111_01100110_1;
      patterns[57226] = 25'b11011111_10001000_01100111_1;
      patterns[57227] = 25'b11011111_10001001_01101000_1;
      patterns[57228] = 25'b11011111_10001010_01101001_1;
      patterns[57229] = 25'b11011111_10001011_01101010_1;
      patterns[57230] = 25'b11011111_10001100_01101011_1;
      patterns[57231] = 25'b11011111_10001101_01101100_1;
      patterns[57232] = 25'b11011111_10001110_01101101_1;
      patterns[57233] = 25'b11011111_10001111_01101110_1;
      patterns[57234] = 25'b11011111_10010000_01101111_1;
      patterns[57235] = 25'b11011111_10010001_01110000_1;
      patterns[57236] = 25'b11011111_10010010_01110001_1;
      patterns[57237] = 25'b11011111_10010011_01110010_1;
      patterns[57238] = 25'b11011111_10010100_01110011_1;
      patterns[57239] = 25'b11011111_10010101_01110100_1;
      patterns[57240] = 25'b11011111_10010110_01110101_1;
      patterns[57241] = 25'b11011111_10010111_01110110_1;
      patterns[57242] = 25'b11011111_10011000_01110111_1;
      patterns[57243] = 25'b11011111_10011001_01111000_1;
      patterns[57244] = 25'b11011111_10011010_01111001_1;
      patterns[57245] = 25'b11011111_10011011_01111010_1;
      patterns[57246] = 25'b11011111_10011100_01111011_1;
      patterns[57247] = 25'b11011111_10011101_01111100_1;
      patterns[57248] = 25'b11011111_10011110_01111101_1;
      patterns[57249] = 25'b11011111_10011111_01111110_1;
      patterns[57250] = 25'b11011111_10100000_01111111_1;
      patterns[57251] = 25'b11011111_10100001_10000000_1;
      patterns[57252] = 25'b11011111_10100010_10000001_1;
      patterns[57253] = 25'b11011111_10100011_10000010_1;
      patterns[57254] = 25'b11011111_10100100_10000011_1;
      patterns[57255] = 25'b11011111_10100101_10000100_1;
      patterns[57256] = 25'b11011111_10100110_10000101_1;
      patterns[57257] = 25'b11011111_10100111_10000110_1;
      patterns[57258] = 25'b11011111_10101000_10000111_1;
      patterns[57259] = 25'b11011111_10101001_10001000_1;
      patterns[57260] = 25'b11011111_10101010_10001001_1;
      patterns[57261] = 25'b11011111_10101011_10001010_1;
      patterns[57262] = 25'b11011111_10101100_10001011_1;
      patterns[57263] = 25'b11011111_10101101_10001100_1;
      patterns[57264] = 25'b11011111_10101110_10001101_1;
      patterns[57265] = 25'b11011111_10101111_10001110_1;
      patterns[57266] = 25'b11011111_10110000_10001111_1;
      patterns[57267] = 25'b11011111_10110001_10010000_1;
      patterns[57268] = 25'b11011111_10110010_10010001_1;
      patterns[57269] = 25'b11011111_10110011_10010010_1;
      patterns[57270] = 25'b11011111_10110100_10010011_1;
      patterns[57271] = 25'b11011111_10110101_10010100_1;
      patterns[57272] = 25'b11011111_10110110_10010101_1;
      patterns[57273] = 25'b11011111_10110111_10010110_1;
      patterns[57274] = 25'b11011111_10111000_10010111_1;
      patterns[57275] = 25'b11011111_10111001_10011000_1;
      patterns[57276] = 25'b11011111_10111010_10011001_1;
      patterns[57277] = 25'b11011111_10111011_10011010_1;
      patterns[57278] = 25'b11011111_10111100_10011011_1;
      patterns[57279] = 25'b11011111_10111101_10011100_1;
      patterns[57280] = 25'b11011111_10111110_10011101_1;
      patterns[57281] = 25'b11011111_10111111_10011110_1;
      patterns[57282] = 25'b11011111_11000000_10011111_1;
      patterns[57283] = 25'b11011111_11000001_10100000_1;
      patterns[57284] = 25'b11011111_11000010_10100001_1;
      patterns[57285] = 25'b11011111_11000011_10100010_1;
      patterns[57286] = 25'b11011111_11000100_10100011_1;
      patterns[57287] = 25'b11011111_11000101_10100100_1;
      patterns[57288] = 25'b11011111_11000110_10100101_1;
      patterns[57289] = 25'b11011111_11000111_10100110_1;
      patterns[57290] = 25'b11011111_11001000_10100111_1;
      patterns[57291] = 25'b11011111_11001001_10101000_1;
      patterns[57292] = 25'b11011111_11001010_10101001_1;
      patterns[57293] = 25'b11011111_11001011_10101010_1;
      patterns[57294] = 25'b11011111_11001100_10101011_1;
      patterns[57295] = 25'b11011111_11001101_10101100_1;
      patterns[57296] = 25'b11011111_11001110_10101101_1;
      patterns[57297] = 25'b11011111_11001111_10101110_1;
      patterns[57298] = 25'b11011111_11010000_10101111_1;
      patterns[57299] = 25'b11011111_11010001_10110000_1;
      patterns[57300] = 25'b11011111_11010010_10110001_1;
      patterns[57301] = 25'b11011111_11010011_10110010_1;
      patterns[57302] = 25'b11011111_11010100_10110011_1;
      patterns[57303] = 25'b11011111_11010101_10110100_1;
      patterns[57304] = 25'b11011111_11010110_10110101_1;
      patterns[57305] = 25'b11011111_11010111_10110110_1;
      patterns[57306] = 25'b11011111_11011000_10110111_1;
      patterns[57307] = 25'b11011111_11011001_10111000_1;
      patterns[57308] = 25'b11011111_11011010_10111001_1;
      patterns[57309] = 25'b11011111_11011011_10111010_1;
      patterns[57310] = 25'b11011111_11011100_10111011_1;
      patterns[57311] = 25'b11011111_11011101_10111100_1;
      patterns[57312] = 25'b11011111_11011110_10111101_1;
      patterns[57313] = 25'b11011111_11011111_10111110_1;
      patterns[57314] = 25'b11011111_11100000_10111111_1;
      patterns[57315] = 25'b11011111_11100001_11000000_1;
      patterns[57316] = 25'b11011111_11100010_11000001_1;
      patterns[57317] = 25'b11011111_11100011_11000010_1;
      patterns[57318] = 25'b11011111_11100100_11000011_1;
      patterns[57319] = 25'b11011111_11100101_11000100_1;
      patterns[57320] = 25'b11011111_11100110_11000101_1;
      patterns[57321] = 25'b11011111_11100111_11000110_1;
      patterns[57322] = 25'b11011111_11101000_11000111_1;
      patterns[57323] = 25'b11011111_11101001_11001000_1;
      patterns[57324] = 25'b11011111_11101010_11001001_1;
      patterns[57325] = 25'b11011111_11101011_11001010_1;
      patterns[57326] = 25'b11011111_11101100_11001011_1;
      patterns[57327] = 25'b11011111_11101101_11001100_1;
      patterns[57328] = 25'b11011111_11101110_11001101_1;
      patterns[57329] = 25'b11011111_11101111_11001110_1;
      patterns[57330] = 25'b11011111_11110000_11001111_1;
      patterns[57331] = 25'b11011111_11110001_11010000_1;
      patterns[57332] = 25'b11011111_11110010_11010001_1;
      patterns[57333] = 25'b11011111_11110011_11010010_1;
      patterns[57334] = 25'b11011111_11110100_11010011_1;
      patterns[57335] = 25'b11011111_11110101_11010100_1;
      patterns[57336] = 25'b11011111_11110110_11010101_1;
      patterns[57337] = 25'b11011111_11110111_11010110_1;
      patterns[57338] = 25'b11011111_11111000_11010111_1;
      patterns[57339] = 25'b11011111_11111001_11011000_1;
      patterns[57340] = 25'b11011111_11111010_11011001_1;
      patterns[57341] = 25'b11011111_11111011_11011010_1;
      patterns[57342] = 25'b11011111_11111100_11011011_1;
      patterns[57343] = 25'b11011111_11111101_11011100_1;
      patterns[57344] = 25'b11011111_11111110_11011101_1;
      patterns[57345] = 25'b11011111_11111111_11011110_1;
      patterns[57346] = 25'b11100000_00000000_11100000_0;
      patterns[57347] = 25'b11100000_00000001_11100001_0;
      patterns[57348] = 25'b11100000_00000010_11100010_0;
      patterns[57349] = 25'b11100000_00000011_11100011_0;
      patterns[57350] = 25'b11100000_00000100_11100100_0;
      patterns[57351] = 25'b11100000_00000101_11100101_0;
      patterns[57352] = 25'b11100000_00000110_11100110_0;
      patterns[57353] = 25'b11100000_00000111_11100111_0;
      patterns[57354] = 25'b11100000_00001000_11101000_0;
      patterns[57355] = 25'b11100000_00001001_11101001_0;
      patterns[57356] = 25'b11100000_00001010_11101010_0;
      patterns[57357] = 25'b11100000_00001011_11101011_0;
      patterns[57358] = 25'b11100000_00001100_11101100_0;
      patterns[57359] = 25'b11100000_00001101_11101101_0;
      patterns[57360] = 25'b11100000_00001110_11101110_0;
      patterns[57361] = 25'b11100000_00001111_11101111_0;
      patterns[57362] = 25'b11100000_00010000_11110000_0;
      patterns[57363] = 25'b11100000_00010001_11110001_0;
      patterns[57364] = 25'b11100000_00010010_11110010_0;
      patterns[57365] = 25'b11100000_00010011_11110011_0;
      patterns[57366] = 25'b11100000_00010100_11110100_0;
      patterns[57367] = 25'b11100000_00010101_11110101_0;
      patterns[57368] = 25'b11100000_00010110_11110110_0;
      patterns[57369] = 25'b11100000_00010111_11110111_0;
      patterns[57370] = 25'b11100000_00011000_11111000_0;
      patterns[57371] = 25'b11100000_00011001_11111001_0;
      patterns[57372] = 25'b11100000_00011010_11111010_0;
      patterns[57373] = 25'b11100000_00011011_11111011_0;
      patterns[57374] = 25'b11100000_00011100_11111100_0;
      patterns[57375] = 25'b11100000_00011101_11111101_0;
      patterns[57376] = 25'b11100000_00011110_11111110_0;
      patterns[57377] = 25'b11100000_00011111_11111111_0;
      patterns[57378] = 25'b11100000_00100000_00000000_1;
      patterns[57379] = 25'b11100000_00100001_00000001_1;
      patterns[57380] = 25'b11100000_00100010_00000010_1;
      patterns[57381] = 25'b11100000_00100011_00000011_1;
      patterns[57382] = 25'b11100000_00100100_00000100_1;
      patterns[57383] = 25'b11100000_00100101_00000101_1;
      patterns[57384] = 25'b11100000_00100110_00000110_1;
      patterns[57385] = 25'b11100000_00100111_00000111_1;
      patterns[57386] = 25'b11100000_00101000_00001000_1;
      patterns[57387] = 25'b11100000_00101001_00001001_1;
      patterns[57388] = 25'b11100000_00101010_00001010_1;
      patterns[57389] = 25'b11100000_00101011_00001011_1;
      patterns[57390] = 25'b11100000_00101100_00001100_1;
      patterns[57391] = 25'b11100000_00101101_00001101_1;
      patterns[57392] = 25'b11100000_00101110_00001110_1;
      patterns[57393] = 25'b11100000_00101111_00001111_1;
      patterns[57394] = 25'b11100000_00110000_00010000_1;
      patterns[57395] = 25'b11100000_00110001_00010001_1;
      patterns[57396] = 25'b11100000_00110010_00010010_1;
      patterns[57397] = 25'b11100000_00110011_00010011_1;
      patterns[57398] = 25'b11100000_00110100_00010100_1;
      patterns[57399] = 25'b11100000_00110101_00010101_1;
      patterns[57400] = 25'b11100000_00110110_00010110_1;
      patterns[57401] = 25'b11100000_00110111_00010111_1;
      patterns[57402] = 25'b11100000_00111000_00011000_1;
      patterns[57403] = 25'b11100000_00111001_00011001_1;
      patterns[57404] = 25'b11100000_00111010_00011010_1;
      patterns[57405] = 25'b11100000_00111011_00011011_1;
      patterns[57406] = 25'b11100000_00111100_00011100_1;
      patterns[57407] = 25'b11100000_00111101_00011101_1;
      patterns[57408] = 25'b11100000_00111110_00011110_1;
      patterns[57409] = 25'b11100000_00111111_00011111_1;
      patterns[57410] = 25'b11100000_01000000_00100000_1;
      patterns[57411] = 25'b11100000_01000001_00100001_1;
      patterns[57412] = 25'b11100000_01000010_00100010_1;
      patterns[57413] = 25'b11100000_01000011_00100011_1;
      patterns[57414] = 25'b11100000_01000100_00100100_1;
      patterns[57415] = 25'b11100000_01000101_00100101_1;
      patterns[57416] = 25'b11100000_01000110_00100110_1;
      patterns[57417] = 25'b11100000_01000111_00100111_1;
      patterns[57418] = 25'b11100000_01001000_00101000_1;
      patterns[57419] = 25'b11100000_01001001_00101001_1;
      patterns[57420] = 25'b11100000_01001010_00101010_1;
      patterns[57421] = 25'b11100000_01001011_00101011_1;
      patterns[57422] = 25'b11100000_01001100_00101100_1;
      patterns[57423] = 25'b11100000_01001101_00101101_1;
      patterns[57424] = 25'b11100000_01001110_00101110_1;
      patterns[57425] = 25'b11100000_01001111_00101111_1;
      patterns[57426] = 25'b11100000_01010000_00110000_1;
      patterns[57427] = 25'b11100000_01010001_00110001_1;
      patterns[57428] = 25'b11100000_01010010_00110010_1;
      patterns[57429] = 25'b11100000_01010011_00110011_1;
      patterns[57430] = 25'b11100000_01010100_00110100_1;
      patterns[57431] = 25'b11100000_01010101_00110101_1;
      patterns[57432] = 25'b11100000_01010110_00110110_1;
      patterns[57433] = 25'b11100000_01010111_00110111_1;
      patterns[57434] = 25'b11100000_01011000_00111000_1;
      patterns[57435] = 25'b11100000_01011001_00111001_1;
      patterns[57436] = 25'b11100000_01011010_00111010_1;
      patterns[57437] = 25'b11100000_01011011_00111011_1;
      patterns[57438] = 25'b11100000_01011100_00111100_1;
      patterns[57439] = 25'b11100000_01011101_00111101_1;
      patterns[57440] = 25'b11100000_01011110_00111110_1;
      patterns[57441] = 25'b11100000_01011111_00111111_1;
      patterns[57442] = 25'b11100000_01100000_01000000_1;
      patterns[57443] = 25'b11100000_01100001_01000001_1;
      patterns[57444] = 25'b11100000_01100010_01000010_1;
      patterns[57445] = 25'b11100000_01100011_01000011_1;
      patterns[57446] = 25'b11100000_01100100_01000100_1;
      patterns[57447] = 25'b11100000_01100101_01000101_1;
      patterns[57448] = 25'b11100000_01100110_01000110_1;
      patterns[57449] = 25'b11100000_01100111_01000111_1;
      patterns[57450] = 25'b11100000_01101000_01001000_1;
      patterns[57451] = 25'b11100000_01101001_01001001_1;
      patterns[57452] = 25'b11100000_01101010_01001010_1;
      patterns[57453] = 25'b11100000_01101011_01001011_1;
      patterns[57454] = 25'b11100000_01101100_01001100_1;
      patterns[57455] = 25'b11100000_01101101_01001101_1;
      patterns[57456] = 25'b11100000_01101110_01001110_1;
      patterns[57457] = 25'b11100000_01101111_01001111_1;
      patterns[57458] = 25'b11100000_01110000_01010000_1;
      patterns[57459] = 25'b11100000_01110001_01010001_1;
      patterns[57460] = 25'b11100000_01110010_01010010_1;
      patterns[57461] = 25'b11100000_01110011_01010011_1;
      patterns[57462] = 25'b11100000_01110100_01010100_1;
      patterns[57463] = 25'b11100000_01110101_01010101_1;
      patterns[57464] = 25'b11100000_01110110_01010110_1;
      patterns[57465] = 25'b11100000_01110111_01010111_1;
      patterns[57466] = 25'b11100000_01111000_01011000_1;
      patterns[57467] = 25'b11100000_01111001_01011001_1;
      patterns[57468] = 25'b11100000_01111010_01011010_1;
      patterns[57469] = 25'b11100000_01111011_01011011_1;
      patterns[57470] = 25'b11100000_01111100_01011100_1;
      patterns[57471] = 25'b11100000_01111101_01011101_1;
      patterns[57472] = 25'b11100000_01111110_01011110_1;
      patterns[57473] = 25'b11100000_01111111_01011111_1;
      patterns[57474] = 25'b11100000_10000000_01100000_1;
      patterns[57475] = 25'b11100000_10000001_01100001_1;
      patterns[57476] = 25'b11100000_10000010_01100010_1;
      patterns[57477] = 25'b11100000_10000011_01100011_1;
      patterns[57478] = 25'b11100000_10000100_01100100_1;
      patterns[57479] = 25'b11100000_10000101_01100101_1;
      patterns[57480] = 25'b11100000_10000110_01100110_1;
      patterns[57481] = 25'b11100000_10000111_01100111_1;
      patterns[57482] = 25'b11100000_10001000_01101000_1;
      patterns[57483] = 25'b11100000_10001001_01101001_1;
      patterns[57484] = 25'b11100000_10001010_01101010_1;
      patterns[57485] = 25'b11100000_10001011_01101011_1;
      patterns[57486] = 25'b11100000_10001100_01101100_1;
      patterns[57487] = 25'b11100000_10001101_01101101_1;
      patterns[57488] = 25'b11100000_10001110_01101110_1;
      patterns[57489] = 25'b11100000_10001111_01101111_1;
      patterns[57490] = 25'b11100000_10010000_01110000_1;
      patterns[57491] = 25'b11100000_10010001_01110001_1;
      patterns[57492] = 25'b11100000_10010010_01110010_1;
      patterns[57493] = 25'b11100000_10010011_01110011_1;
      patterns[57494] = 25'b11100000_10010100_01110100_1;
      patterns[57495] = 25'b11100000_10010101_01110101_1;
      patterns[57496] = 25'b11100000_10010110_01110110_1;
      patterns[57497] = 25'b11100000_10010111_01110111_1;
      patterns[57498] = 25'b11100000_10011000_01111000_1;
      patterns[57499] = 25'b11100000_10011001_01111001_1;
      patterns[57500] = 25'b11100000_10011010_01111010_1;
      patterns[57501] = 25'b11100000_10011011_01111011_1;
      patterns[57502] = 25'b11100000_10011100_01111100_1;
      patterns[57503] = 25'b11100000_10011101_01111101_1;
      patterns[57504] = 25'b11100000_10011110_01111110_1;
      patterns[57505] = 25'b11100000_10011111_01111111_1;
      patterns[57506] = 25'b11100000_10100000_10000000_1;
      patterns[57507] = 25'b11100000_10100001_10000001_1;
      patterns[57508] = 25'b11100000_10100010_10000010_1;
      patterns[57509] = 25'b11100000_10100011_10000011_1;
      patterns[57510] = 25'b11100000_10100100_10000100_1;
      patterns[57511] = 25'b11100000_10100101_10000101_1;
      patterns[57512] = 25'b11100000_10100110_10000110_1;
      patterns[57513] = 25'b11100000_10100111_10000111_1;
      patterns[57514] = 25'b11100000_10101000_10001000_1;
      patterns[57515] = 25'b11100000_10101001_10001001_1;
      patterns[57516] = 25'b11100000_10101010_10001010_1;
      patterns[57517] = 25'b11100000_10101011_10001011_1;
      patterns[57518] = 25'b11100000_10101100_10001100_1;
      patterns[57519] = 25'b11100000_10101101_10001101_1;
      patterns[57520] = 25'b11100000_10101110_10001110_1;
      patterns[57521] = 25'b11100000_10101111_10001111_1;
      patterns[57522] = 25'b11100000_10110000_10010000_1;
      patterns[57523] = 25'b11100000_10110001_10010001_1;
      patterns[57524] = 25'b11100000_10110010_10010010_1;
      patterns[57525] = 25'b11100000_10110011_10010011_1;
      patterns[57526] = 25'b11100000_10110100_10010100_1;
      patterns[57527] = 25'b11100000_10110101_10010101_1;
      patterns[57528] = 25'b11100000_10110110_10010110_1;
      patterns[57529] = 25'b11100000_10110111_10010111_1;
      patterns[57530] = 25'b11100000_10111000_10011000_1;
      patterns[57531] = 25'b11100000_10111001_10011001_1;
      patterns[57532] = 25'b11100000_10111010_10011010_1;
      patterns[57533] = 25'b11100000_10111011_10011011_1;
      patterns[57534] = 25'b11100000_10111100_10011100_1;
      patterns[57535] = 25'b11100000_10111101_10011101_1;
      patterns[57536] = 25'b11100000_10111110_10011110_1;
      patterns[57537] = 25'b11100000_10111111_10011111_1;
      patterns[57538] = 25'b11100000_11000000_10100000_1;
      patterns[57539] = 25'b11100000_11000001_10100001_1;
      patterns[57540] = 25'b11100000_11000010_10100010_1;
      patterns[57541] = 25'b11100000_11000011_10100011_1;
      patterns[57542] = 25'b11100000_11000100_10100100_1;
      patterns[57543] = 25'b11100000_11000101_10100101_1;
      patterns[57544] = 25'b11100000_11000110_10100110_1;
      patterns[57545] = 25'b11100000_11000111_10100111_1;
      patterns[57546] = 25'b11100000_11001000_10101000_1;
      patterns[57547] = 25'b11100000_11001001_10101001_1;
      patterns[57548] = 25'b11100000_11001010_10101010_1;
      patterns[57549] = 25'b11100000_11001011_10101011_1;
      patterns[57550] = 25'b11100000_11001100_10101100_1;
      patterns[57551] = 25'b11100000_11001101_10101101_1;
      patterns[57552] = 25'b11100000_11001110_10101110_1;
      patterns[57553] = 25'b11100000_11001111_10101111_1;
      patterns[57554] = 25'b11100000_11010000_10110000_1;
      patterns[57555] = 25'b11100000_11010001_10110001_1;
      patterns[57556] = 25'b11100000_11010010_10110010_1;
      patterns[57557] = 25'b11100000_11010011_10110011_1;
      patterns[57558] = 25'b11100000_11010100_10110100_1;
      patterns[57559] = 25'b11100000_11010101_10110101_1;
      patterns[57560] = 25'b11100000_11010110_10110110_1;
      patterns[57561] = 25'b11100000_11010111_10110111_1;
      patterns[57562] = 25'b11100000_11011000_10111000_1;
      patterns[57563] = 25'b11100000_11011001_10111001_1;
      patterns[57564] = 25'b11100000_11011010_10111010_1;
      patterns[57565] = 25'b11100000_11011011_10111011_1;
      patterns[57566] = 25'b11100000_11011100_10111100_1;
      patterns[57567] = 25'b11100000_11011101_10111101_1;
      patterns[57568] = 25'b11100000_11011110_10111110_1;
      patterns[57569] = 25'b11100000_11011111_10111111_1;
      patterns[57570] = 25'b11100000_11100000_11000000_1;
      patterns[57571] = 25'b11100000_11100001_11000001_1;
      patterns[57572] = 25'b11100000_11100010_11000010_1;
      patterns[57573] = 25'b11100000_11100011_11000011_1;
      patterns[57574] = 25'b11100000_11100100_11000100_1;
      patterns[57575] = 25'b11100000_11100101_11000101_1;
      patterns[57576] = 25'b11100000_11100110_11000110_1;
      patterns[57577] = 25'b11100000_11100111_11000111_1;
      patterns[57578] = 25'b11100000_11101000_11001000_1;
      patterns[57579] = 25'b11100000_11101001_11001001_1;
      patterns[57580] = 25'b11100000_11101010_11001010_1;
      patterns[57581] = 25'b11100000_11101011_11001011_1;
      patterns[57582] = 25'b11100000_11101100_11001100_1;
      patterns[57583] = 25'b11100000_11101101_11001101_1;
      patterns[57584] = 25'b11100000_11101110_11001110_1;
      patterns[57585] = 25'b11100000_11101111_11001111_1;
      patterns[57586] = 25'b11100000_11110000_11010000_1;
      patterns[57587] = 25'b11100000_11110001_11010001_1;
      patterns[57588] = 25'b11100000_11110010_11010010_1;
      patterns[57589] = 25'b11100000_11110011_11010011_1;
      patterns[57590] = 25'b11100000_11110100_11010100_1;
      patterns[57591] = 25'b11100000_11110101_11010101_1;
      patterns[57592] = 25'b11100000_11110110_11010110_1;
      patterns[57593] = 25'b11100000_11110111_11010111_1;
      patterns[57594] = 25'b11100000_11111000_11011000_1;
      patterns[57595] = 25'b11100000_11111001_11011001_1;
      patterns[57596] = 25'b11100000_11111010_11011010_1;
      patterns[57597] = 25'b11100000_11111011_11011011_1;
      patterns[57598] = 25'b11100000_11111100_11011100_1;
      patterns[57599] = 25'b11100000_11111101_11011101_1;
      patterns[57600] = 25'b11100000_11111110_11011110_1;
      patterns[57601] = 25'b11100000_11111111_11011111_1;
      patterns[57602] = 25'b11100001_00000000_11100001_0;
      patterns[57603] = 25'b11100001_00000001_11100010_0;
      patterns[57604] = 25'b11100001_00000010_11100011_0;
      patterns[57605] = 25'b11100001_00000011_11100100_0;
      patterns[57606] = 25'b11100001_00000100_11100101_0;
      patterns[57607] = 25'b11100001_00000101_11100110_0;
      patterns[57608] = 25'b11100001_00000110_11100111_0;
      patterns[57609] = 25'b11100001_00000111_11101000_0;
      patterns[57610] = 25'b11100001_00001000_11101001_0;
      patterns[57611] = 25'b11100001_00001001_11101010_0;
      patterns[57612] = 25'b11100001_00001010_11101011_0;
      patterns[57613] = 25'b11100001_00001011_11101100_0;
      patterns[57614] = 25'b11100001_00001100_11101101_0;
      patterns[57615] = 25'b11100001_00001101_11101110_0;
      patterns[57616] = 25'b11100001_00001110_11101111_0;
      patterns[57617] = 25'b11100001_00001111_11110000_0;
      patterns[57618] = 25'b11100001_00010000_11110001_0;
      patterns[57619] = 25'b11100001_00010001_11110010_0;
      patterns[57620] = 25'b11100001_00010010_11110011_0;
      patterns[57621] = 25'b11100001_00010011_11110100_0;
      patterns[57622] = 25'b11100001_00010100_11110101_0;
      patterns[57623] = 25'b11100001_00010101_11110110_0;
      patterns[57624] = 25'b11100001_00010110_11110111_0;
      patterns[57625] = 25'b11100001_00010111_11111000_0;
      patterns[57626] = 25'b11100001_00011000_11111001_0;
      patterns[57627] = 25'b11100001_00011001_11111010_0;
      patterns[57628] = 25'b11100001_00011010_11111011_0;
      patterns[57629] = 25'b11100001_00011011_11111100_0;
      patterns[57630] = 25'b11100001_00011100_11111101_0;
      patterns[57631] = 25'b11100001_00011101_11111110_0;
      patterns[57632] = 25'b11100001_00011110_11111111_0;
      patterns[57633] = 25'b11100001_00011111_00000000_1;
      patterns[57634] = 25'b11100001_00100000_00000001_1;
      patterns[57635] = 25'b11100001_00100001_00000010_1;
      patterns[57636] = 25'b11100001_00100010_00000011_1;
      patterns[57637] = 25'b11100001_00100011_00000100_1;
      patterns[57638] = 25'b11100001_00100100_00000101_1;
      patterns[57639] = 25'b11100001_00100101_00000110_1;
      patterns[57640] = 25'b11100001_00100110_00000111_1;
      patterns[57641] = 25'b11100001_00100111_00001000_1;
      patterns[57642] = 25'b11100001_00101000_00001001_1;
      patterns[57643] = 25'b11100001_00101001_00001010_1;
      patterns[57644] = 25'b11100001_00101010_00001011_1;
      patterns[57645] = 25'b11100001_00101011_00001100_1;
      patterns[57646] = 25'b11100001_00101100_00001101_1;
      patterns[57647] = 25'b11100001_00101101_00001110_1;
      patterns[57648] = 25'b11100001_00101110_00001111_1;
      patterns[57649] = 25'b11100001_00101111_00010000_1;
      patterns[57650] = 25'b11100001_00110000_00010001_1;
      patterns[57651] = 25'b11100001_00110001_00010010_1;
      patterns[57652] = 25'b11100001_00110010_00010011_1;
      patterns[57653] = 25'b11100001_00110011_00010100_1;
      patterns[57654] = 25'b11100001_00110100_00010101_1;
      patterns[57655] = 25'b11100001_00110101_00010110_1;
      patterns[57656] = 25'b11100001_00110110_00010111_1;
      patterns[57657] = 25'b11100001_00110111_00011000_1;
      patterns[57658] = 25'b11100001_00111000_00011001_1;
      patterns[57659] = 25'b11100001_00111001_00011010_1;
      patterns[57660] = 25'b11100001_00111010_00011011_1;
      patterns[57661] = 25'b11100001_00111011_00011100_1;
      patterns[57662] = 25'b11100001_00111100_00011101_1;
      patterns[57663] = 25'b11100001_00111101_00011110_1;
      patterns[57664] = 25'b11100001_00111110_00011111_1;
      patterns[57665] = 25'b11100001_00111111_00100000_1;
      patterns[57666] = 25'b11100001_01000000_00100001_1;
      patterns[57667] = 25'b11100001_01000001_00100010_1;
      patterns[57668] = 25'b11100001_01000010_00100011_1;
      patterns[57669] = 25'b11100001_01000011_00100100_1;
      patterns[57670] = 25'b11100001_01000100_00100101_1;
      patterns[57671] = 25'b11100001_01000101_00100110_1;
      patterns[57672] = 25'b11100001_01000110_00100111_1;
      patterns[57673] = 25'b11100001_01000111_00101000_1;
      patterns[57674] = 25'b11100001_01001000_00101001_1;
      patterns[57675] = 25'b11100001_01001001_00101010_1;
      patterns[57676] = 25'b11100001_01001010_00101011_1;
      patterns[57677] = 25'b11100001_01001011_00101100_1;
      patterns[57678] = 25'b11100001_01001100_00101101_1;
      patterns[57679] = 25'b11100001_01001101_00101110_1;
      patterns[57680] = 25'b11100001_01001110_00101111_1;
      patterns[57681] = 25'b11100001_01001111_00110000_1;
      patterns[57682] = 25'b11100001_01010000_00110001_1;
      patterns[57683] = 25'b11100001_01010001_00110010_1;
      patterns[57684] = 25'b11100001_01010010_00110011_1;
      patterns[57685] = 25'b11100001_01010011_00110100_1;
      patterns[57686] = 25'b11100001_01010100_00110101_1;
      patterns[57687] = 25'b11100001_01010101_00110110_1;
      patterns[57688] = 25'b11100001_01010110_00110111_1;
      patterns[57689] = 25'b11100001_01010111_00111000_1;
      patterns[57690] = 25'b11100001_01011000_00111001_1;
      patterns[57691] = 25'b11100001_01011001_00111010_1;
      patterns[57692] = 25'b11100001_01011010_00111011_1;
      patterns[57693] = 25'b11100001_01011011_00111100_1;
      patterns[57694] = 25'b11100001_01011100_00111101_1;
      patterns[57695] = 25'b11100001_01011101_00111110_1;
      patterns[57696] = 25'b11100001_01011110_00111111_1;
      patterns[57697] = 25'b11100001_01011111_01000000_1;
      patterns[57698] = 25'b11100001_01100000_01000001_1;
      patterns[57699] = 25'b11100001_01100001_01000010_1;
      patterns[57700] = 25'b11100001_01100010_01000011_1;
      patterns[57701] = 25'b11100001_01100011_01000100_1;
      patterns[57702] = 25'b11100001_01100100_01000101_1;
      patterns[57703] = 25'b11100001_01100101_01000110_1;
      patterns[57704] = 25'b11100001_01100110_01000111_1;
      patterns[57705] = 25'b11100001_01100111_01001000_1;
      patterns[57706] = 25'b11100001_01101000_01001001_1;
      patterns[57707] = 25'b11100001_01101001_01001010_1;
      patterns[57708] = 25'b11100001_01101010_01001011_1;
      patterns[57709] = 25'b11100001_01101011_01001100_1;
      patterns[57710] = 25'b11100001_01101100_01001101_1;
      patterns[57711] = 25'b11100001_01101101_01001110_1;
      patterns[57712] = 25'b11100001_01101110_01001111_1;
      patterns[57713] = 25'b11100001_01101111_01010000_1;
      patterns[57714] = 25'b11100001_01110000_01010001_1;
      patterns[57715] = 25'b11100001_01110001_01010010_1;
      patterns[57716] = 25'b11100001_01110010_01010011_1;
      patterns[57717] = 25'b11100001_01110011_01010100_1;
      patterns[57718] = 25'b11100001_01110100_01010101_1;
      patterns[57719] = 25'b11100001_01110101_01010110_1;
      patterns[57720] = 25'b11100001_01110110_01010111_1;
      patterns[57721] = 25'b11100001_01110111_01011000_1;
      patterns[57722] = 25'b11100001_01111000_01011001_1;
      patterns[57723] = 25'b11100001_01111001_01011010_1;
      patterns[57724] = 25'b11100001_01111010_01011011_1;
      patterns[57725] = 25'b11100001_01111011_01011100_1;
      patterns[57726] = 25'b11100001_01111100_01011101_1;
      patterns[57727] = 25'b11100001_01111101_01011110_1;
      patterns[57728] = 25'b11100001_01111110_01011111_1;
      patterns[57729] = 25'b11100001_01111111_01100000_1;
      patterns[57730] = 25'b11100001_10000000_01100001_1;
      patterns[57731] = 25'b11100001_10000001_01100010_1;
      patterns[57732] = 25'b11100001_10000010_01100011_1;
      patterns[57733] = 25'b11100001_10000011_01100100_1;
      patterns[57734] = 25'b11100001_10000100_01100101_1;
      patterns[57735] = 25'b11100001_10000101_01100110_1;
      patterns[57736] = 25'b11100001_10000110_01100111_1;
      patterns[57737] = 25'b11100001_10000111_01101000_1;
      patterns[57738] = 25'b11100001_10001000_01101001_1;
      patterns[57739] = 25'b11100001_10001001_01101010_1;
      patterns[57740] = 25'b11100001_10001010_01101011_1;
      patterns[57741] = 25'b11100001_10001011_01101100_1;
      patterns[57742] = 25'b11100001_10001100_01101101_1;
      patterns[57743] = 25'b11100001_10001101_01101110_1;
      patterns[57744] = 25'b11100001_10001110_01101111_1;
      patterns[57745] = 25'b11100001_10001111_01110000_1;
      patterns[57746] = 25'b11100001_10010000_01110001_1;
      patterns[57747] = 25'b11100001_10010001_01110010_1;
      patterns[57748] = 25'b11100001_10010010_01110011_1;
      patterns[57749] = 25'b11100001_10010011_01110100_1;
      patterns[57750] = 25'b11100001_10010100_01110101_1;
      patterns[57751] = 25'b11100001_10010101_01110110_1;
      patterns[57752] = 25'b11100001_10010110_01110111_1;
      patterns[57753] = 25'b11100001_10010111_01111000_1;
      patterns[57754] = 25'b11100001_10011000_01111001_1;
      patterns[57755] = 25'b11100001_10011001_01111010_1;
      patterns[57756] = 25'b11100001_10011010_01111011_1;
      patterns[57757] = 25'b11100001_10011011_01111100_1;
      patterns[57758] = 25'b11100001_10011100_01111101_1;
      patterns[57759] = 25'b11100001_10011101_01111110_1;
      patterns[57760] = 25'b11100001_10011110_01111111_1;
      patterns[57761] = 25'b11100001_10011111_10000000_1;
      patterns[57762] = 25'b11100001_10100000_10000001_1;
      patterns[57763] = 25'b11100001_10100001_10000010_1;
      patterns[57764] = 25'b11100001_10100010_10000011_1;
      patterns[57765] = 25'b11100001_10100011_10000100_1;
      patterns[57766] = 25'b11100001_10100100_10000101_1;
      patterns[57767] = 25'b11100001_10100101_10000110_1;
      patterns[57768] = 25'b11100001_10100110_10000111_1;
      patterns[57769] = 25'b11100001_10100111_10001000_1;
      patterns[57770] = 25'b11100001_10101000_10001001_1;
      patterns[57771] = 25'b11100001_10101001_10001010_1;
      patterns[57772] = 25'b11100001_10101010_10001011_1;
      patterns[57773] = 25'b11100001_10101011_10001100_1;
      patterns[57774] = 25'b11100001_10101100_10001101_1;
      patterns[57775] = 25'b11100001_10101101_10001110_1;
      patterns[57776] = 25'b11100001_10101110_10001111_1;
      patterns[57777] = 25'b11100001_10101111_10010000_1;
      patterns[57778] = 25'b11100001_10110000_10010001_1;
      patterns[57779] = 25'b11100001_10110001_10010010_1;
      patterns[57780] = 25'b11100001_10110010_10010011_1;
      patterns[57781] = 25'b11100001_10110011_10010100_1;
      patterns[57782] = 25'b11100001_10110100_10010101_1;
      patterns[57783] = 25'b11100001_10110101_10010110_1;
      patterns[57784] = 25'b11100001_10110110_10010111_1;
      patterns[57785] = 25'b11100001_10110111_10011000_1;
      patterns[57786] = 25'b11100001_10111000_10011001_1;
      patterns[57787] = 25'b11100001_10111001_10011010_1;
      patterns[57788] = 25'b11100001_10111010_10011011_1;
      patterns[57789] = 25'b11100001_10111011_10011100_1;
      patterns[57790] = 25'b11100001_10111100_10011101_1;
      patterns[57791] = 25'b11100001_10111101_10011110_1;
      patterns[57792] = 25'b11100001_10111110_10011111_1;
      patterns[57793] = 25'b11100001_10111111_10100000_1;
      patterns[57794] = 25'b11100001_11000000_10100001_1;
      patterns[57795] = 25'b11100001_11000001_10100010_1;
      patterns[57796] = 25'b11100001_11000010_10100011_1;
      patterns[57797] = 25'b11100001_11000011_10100100_1;
      patterns[57798] = 25'b11100001_11000100_10100101_1;
      patterns[57799] = 25'b11100001_11000101_10100110_1;
      patterns[57800] = 25'b11100001_11000110_10100111_1;
      patterns[57801] = 25'b11100001_11000111_10101000_1;
      patterns[57802] = 25'b11100001_11001000_10101001_1;
      patterns[57803] = 25'b11100001_11001001_10101010_1;
      patterns[57804] = 25'b11100001_11001010_10101011_1;
      patterns[57805] = 25'b11100001_11001011_10101100_1;
      patterns[57806] = 25'b11100001_11001100_10101101_1;
      patterns[57807] = 25'b11100001_11001101_10101110_1;
      patterns[57808] = 25'b11100001_11001110_10101111_1;
      patterns[57809] = 25'b11100001_11001111_10110000_1;
      patterns[57810] = 25'b11100001_11010000_10110001_1;
      patterns[57811] = 25'b11100001_11010001_10110010_1;
      patterns[57812] = 25'b11100001_11010010_10110011_1;
      patterns[57813] = 25'b11100001_11010011_10110100_1;
      patterns[57814] = 25'b11100001_11010100_10110101_1;
      patterns[57815] = 25'b11100001_11010101_10110110_1;
      patterns[57816] = 25'b11100001_11010110_10110111_1;
      patterns[57817] = 25'b11100001_11010111_10111000_1;
      patterns[57818] = 25'b11100001_11011000_10111001_1;
      patterns[57819] = 25'b11100001_11011001_10111010_1;
      patterns[57820] = 25'b11100001_11011010_10111011_1;
      patterns[57821] = 25'b11100001_11011011_10111100_1;
      patterns[57822] = 25'b11100001_11011100_10111101_1;
      patterns[57823] = 25'b11100001_11011101_10111110_1;
      patterns[57824] = 25'b11100001_11011110_10111111_1;
      patterns[57825] = 25'b11100001_11011111_11000000_1;
      patterns[57826] = 25'b11100001_11100000_11000001_1;
      patterns[57827] = 25'b11100001_11100001_11000010_1;
      patterns[57828] = 25'b11100001_11100010_11000011_1;
      patterns[57829] = 25'b11100001_11100011_11000100_1;
      patterns[57830] = 25'b11100001_11100100_11000101_1;
      patterns[57831] = 25'b11100001_11100101_11000110_1;
      patterns[57832] = 25'b11100001_11100110_11000111_1;
      patterns[57833] = 25'b11100001_11100111_11001000_1;
      patterns[57834] = 25'b11100001_11101000_11001001_1;
      patterns[57835] = 25'b11100001_11101001_11001010_1;
      patterns[57836] = 25'b11100001_11101010_11001011_1;
      patterns[57837] = 25'b11100001_11101011_11001100_1;
      patterns[57838] = 25'b11100001_11101100_11001101_1;
      patterns[57839] = 25'b11100001_11101101_11001110_1;
      patterns[57840] = 25'b11100001_11101110_11001111_1;
      patterns[57841] = 25'b11100001_11101111_11010000_1;
      patterns[57842] = 25'b11100001_11110000_11010001_1;
      patterns[57843] = 25'b11100001_11110001_11010010_1;
      patterns[57844] = 25'b11100001_11110010_11010011_1;
      patterns[57845] = 25'b11100001_11110011_11010100_1;
      patterns[57846] = 25'b11100001_11110100_11010101_1;
      patterns[57847] = 25'b11100001_11110101_11010110_1;
      patterns[57848] = 25'b11100001_11110110_11010111_1;
      patterns[57849] = 25'b11100001_11110111_11011000_1;
      patterns[57850] = 25'b11100001_11111000_11011001_1;
      patterns[57851] = 25'b11100001_11111001_11011010_1;
      patterns[57852] = 25'b11100001_11111010_11011011_1;
      patterns[57853] = 25'b11100001_11111011_11011100_1;
      patterns[57854] = 25'b11100001_11111100_11011101_1;
      patterns[57855] = 25'b11100001_11111101_11011110_1;
      patterns[57856] = 25'b11100001_11111110_11011111_1;
      patterns[57857] = 25'b11100001_11111111_11100000_1;
      patterns[57858] = 25'b11100010_00000000_11100010_0;
      patterns[57859] = 25'b11100010_00000001_11100011_0;
      patterns[57860] = 25'b11100010_00000010_11100100_0;
      patterns[57861] = 25'b11100010_00000011_11100101_0;
      patterns[57862] = 25'b11100010_00000100_11100110_0;
      patterns[57863] = 25'b11100010_00000101_11100111_0;
      patterns[57864] = 25'b11100010_00000110_11101000_0;
      patterns[57865] = 25'b11100010_00000111_11101001_0;
      patterns[57866] = 25'b11100010_00001000_11101010_0;
      patterns[57867] = 25'b11100010_00001001_11101011_0;
      patterns[57868] = 25'b11100010_00001010_11101100_0;
      patterns[57869] = 25'b11100010_00001011_11101101_0;
      patterns[57870] = 25'b11100010_00001100_11101110_0;
      patterns[57871] = 25'b11100010_00001101_11101111_0;
      patterns[57872] = 25'b11100010_00001110_11110000_0;
      patterns[57873] = 25'b11100010_00001111_11110001_0;
      patterns[57874] = 25'b11100010_00010000_11110010_0;
      patterns[57875] = 25'b11100010_00010001_11110011_0;
      patterns[57876] = 25'b11100010_00010010_11110100_0;
      patterns[57877] = 25'b11100010_00010011_11110101_0;
      patterns[57878] = 25'b11100010_00010100_11110110_0;
      patterns[57879] = 25'b11100010_00010101_11110111_0;
      patterns[57880] = 25'b11100010_00010110_11111000_0;
      patterns[57881] = 25'b11100010_00010111_11111001_0;
      patterns[57882] = 25'b11100010_00011000_11111010_0;
      patterns[57883] = 25'b11100010_00011001_11111011_0;
      patterns[57884] = 25'b11100010_00011010_11111100_0;
      patterns[57885] = 25'b11100010_00011011_11111101_0;
      patterns[57886] = 25'b11100010_00011100_11111110_0;
      patterns[57887] = 25'b11100010_00011101_11111111_0;
      patterns[57888] = 25'b11100010_00011110_00000000_1;
      patterns[57889] = 25'b11100010_00011111_00000001_1;
      patterns[57890] = 25'b11100010_00100000_00000010_1;
      patterns[57891] = 25'b11100010_00100001_00000011_1;
      patterns[57892] = 25'b11100010_00100010_00000100_1;
      patterns[57893] = 25'b11100010_00100011_00000101_1;
      patterns[57894] = 25'b11100010_00100100_00000110_1;
      patterns[57895] = 25'b11100010_00100101_00000111_1;
      patterns[57896] = 25'b11100010_00100110_00001000_1;
      patterns[57897] = 25'b11100010_00100111_00001001_1;
      patterns[57898] = 25'b11100010_00101000_00001010_1;
      patterns[57899] = 25'b11100010_00101001_00001011_1;
      patterns[57900] = 25'b11100010_00101010_00001100_1;
      patterns[57901] = 25'b11100010_00101011_00001101_1;
      patterns[57902] = 25'b11100010_00101100_00001110_1;
      patterns[57903] = 25'b11100010_00101101_00001111_1;
      patterns[57904] = 25'b11100010_00101110_00010000_1;
      patterns[57905] = 25'b11100010_00101111_00010001_1;
      patterns[57906] = 25'b11100010_00110000_00010010_1;
      patterns[57907] = 25'b11100010_00110001_00010011_1;
      patterns[57908] = 25'b11100010_00110010_00010100_1;
      patterns[57909] = 25'b11100010_00110011_00010101_1;
      patterns[57910] = 25'b11100010_00110100_00010110_1;
      patterns[57911] = 25'b11100010_00110101_00010111_1;
      patterns[57912] = 25'b11100010_00110110_00011000_1;
      patterns[57913] = 25'b11100010_00110111_00011001_1;
      patterns[57914] = 25'b11100010_00111000_00011010_1;
      patterns[57915] = 25'b11100010_00111001_00011011_1;
      patterns[57916] = 25'b11100010_00111010_00011100_1;
      patterns[57917] = 25'b11100010_00111011_00011101_1;
      patterns[57918] = 25'b11100010_00111100_00011110_1;
      patterns[57919] = 25'b11100010_00111101_00011111_1;
      patterns[57920] = 25'b11100010_00111110_00100000_1;
      patterns[57921] = 25'b11100010_00111111_00100001_1;
      patterns[57922] = 25'b11100010_01000000_00100010_1;
      patterns[57923] = 25'b11100010_01000001_00100011_1;
      patterns[57924] = 25'b11100010_01000010_00100100_1;
      patterns[57925] = 25'b11100010_01000011_00100101_1;
      patterns[57926] = 25'b11100010_01000100_00100110_1;
      patterns[57927] = 25'b11100010_01000101_00100111_1;
      patterns[57928] = 25'b11100010_01000110_00101000_1;
      patterns[57929] = 25'b11100010_01000111_00101001_1;
      patterns[57930] = 25'b11100010_01001000_00101010_1;
      patterns[57931] = 25'b11100010_01001001_00101011_1;
      patterns[57932] = 25'b11100010_01001010_00101100_1;
      patterns[57933] = 25'b11100010_01001011_00101101_1;
      patterns[57934] = 25'b11100010_01001100_00101110_1;
      patterns[57935] = 25'b11100010_01001101_00101111_1;
      patterns[57936] = 25'b11100010_01001110_00110000_1;
      patterns[57937] = 25'b11100010_01001111_00110001_1;
      patterns[57938] = 25'b11100010_01010000_00110010_1;
      patterns[57939] = 25'b11100010_01010001_00110011_1;
      patterns[57940] = 25'b11100010_01010010_00110100_1;
      patterns[57941] = 25'b11100010_01010011_00110101_1;
      patterns[57942] = 25'b11100010_01010100_00110110_1;
      patterns[57943] = 25'b11100010_01010101_00110111_1;
      patterns[57944] = 25'b11100010_01010110_00111000_1;
      patterns[57945] = 25'b11100010_01010111_00111001_1;
      patterns[57946] = 25'b11100010_01011000_00111010_1;
      patterns[57947] = 25'b11100010_01011001_00111011_1;
      patterns[57948] = 25'b11100010_01011010_00111100_1;
      patterns[57949] = 25'b11100010_01011011_00111101_1;
      patterns[57950] = 25'b11100010_01011100_00111110_1;
      patterns[57951] = 25'b11100010_01011101_00111111_1;
      patterns[57952] = 25'b11100010_01011110_01000000_1;
      patterns[57953] = 25'b11100010_01011111_01000001_1;
      patterns[57954] = 25'b11100010_01100000_01000010_1;
      patterns[57955] = 25'b11100010_01100001_01000011_1;
      patterns[57956] = 25'b11100010_01100010_01000100_1;
      patterns[57957] = 25'b11100010_01100011_01000101_1;
      patterns[57958] = 25'b11100010_01100100_01000110_1;
      patterns[57959] = 25'b11100010_01100101_01000111_1;
      patterns[57960] = 25'b11100010_01100110_01001000_1;
      patterns[57961] = 25'b11100010_01100111_01001001_1;
      patterns[57962] = 25'b11100010_01101000_01001010_1;
      patterns[57963] = 25'b11100010_01101001_01001011_1;
      patterns[57964] = 25'b11100010_01101010_01001100_1;
      patterns[57965] = 25'b11100010_01101011_01001101_1;
      patterns[57966] = 25'b11100010_01101100_01001110_1;
      patterns[57967] = 25'b11100010_01101101_01001111_1;
      patterns[57968] = 25'b11100010_01101110_01010000_1;
      patterns[57969] = 25'b11100010_01101111_01010001_1;
      patterns[57970] = 25'b11100010_01110000_01010010_1;
      patterns[57971] = 25'b11100010_01110001_01010011_1;
      patterns[57972] = 25'b11100010_01110010_01010100_1;
      patterns[57973] = 25'b11100010_01110011_01010101_1;
      patterns[57974] = 25'b11100010_01110100_01010110_1;
      patterns[57975] = 25'b11100010_01110101_01010111_1;
      patterns[57976] = 25'b11100010_01110110_01011000_1;
      patterns[57977] = 25'b11100010_01110111_01011001_1;
      patterns[57978] = 25'b11100010_01111000_01011010_1;
      patterns[57979] = 25'b11100010_01111001_01011011_1;
      patterns[57980] = 25'b11100010_01111010_01011100_1;
      patterns[57981] = 25'b11100010_01111011_01011101_1;
      patterns[57982] = 25'b11100010_01111100_01011110_1;
      patterns[57983] = 25'b11100010_01111101_01011111_1;
      patterns[57984] = 25'b11100010_01111110_01100000_1;
      patterns[57985] = 25'b11100010_01111111_01100001_1;
      patterns[57986] = 25'b11100010_10000000_01100010_1;
      patterns[57987] = 25'b11100010_10000001_01100011_1;
      patterns[57988] = 25'b11100010_10000010_01100100_1;
      patterns[57989] = 25'b11100010_10000011_01100101_1;
      patterns[57990] = 25'b11100010_10000100_01100110_1;
      patterns[57991] = 25'b11100010_10000101_01100111_1;
      patterns[57992] = 25'b11100010_10000110_01101000_1;
      patterns[57993] = 25'b11100010_10000111_01101001_1;
      patterns[57994] = 25'b11100010_10001000_01101010_1;
      patterns[57995] = 25'b11100010_10001001_01101011_1;
      patterns[57996] = 25'b11100010_10001010_01101100_1;
      patterns[57997] = 25'b11100010_10001011_01101101_1;
      patterns[57998] = 25'b11100010_10001100_01101110_1;
      patterns[57999] = 25'b11100010_10001101_01101111_1;
      patterns[58000] = 25'b11100010_10001110_01110000_1;
      patterns[58001] = 25'b11100010_10001111_01110001_1;
      patterns[58002] = 25'b11100010_10010000_01110010_1;
      patterns[58003] = 25'b11100010_10010001_01110011_1;
      patterns[58004] = 25'b11100010_10010010_01110100_1;
      patterns[58005] = 25'b11100010_10010011_01110101_1;
      patterns[58006] = 25'b11100010_10010100_01110110_1;
      patterns[58007] = 25'b11100010_10010101_01110111_1;
      patterns[58008] = 25'b11100010_10010110_01111000_1;
      patterns[58009] = 25'b11100010_10010111_01111001_1;
      patterns[58010] = 25'b11100010_10011000_01111010_1;
      patterns[58011] = 25'b11100010_10011001_01111011_1;
      patterns[58012] = 25'b11100010_10011010_01111100_1;
      patterns[58013] = 25'b11100010_10011011_01111101_1;
      patterns[58014] = 25'b11100010_10011100_01111110_1;
      patterns[58015] = 25'b11100010_10011101_01111111_1;
      patterns[58016] = 25'b11100010_10011110_10000000_1;
      patterns[58017] = 25'b11100010_10011111_10000001_1;
      patterns[58018] = 25'b11100010_10100000_10000010_1;
      patterns[58019] = 25'b11100010_10100001_10000011_1;
      patterns[58020] = 25'b11100010_10100010_10000100_1;
      patterns[58021] = 25'b11100010_10100011_10000101_1;
      patterns[58022] = 25'b11100010_10100100_10000110_1;
      patterns[58023] = 25'b11100010_10100101_10000111_1;
      patterns[58024] = 25'b11100010_10100110_10001000_1;
      patterns[58025] = 25'b11100010_10100111_10001001_1;
      patterns[58026] = 25'b11100010_10101000_10001010_1;
      patterns[58027] = 25'b11100010_10101001_10001011_1;
      patterns[58028] = 25'b11100010_10101010_10001100_1;
      patterns[58029] = 25'b11100010_10101011_10001101_1;
      patterns[58030] = 25'b11100010_10101100_10001110_1;
      patterns[58031] = 25'b11100010_10101101_10001111_1;
      patterns[58032] = 25'b11100010_10101110_10010000_1;
      patterns[58033] = 25'b11100010_10101111_10010001_1;
      patterns[58034] = 25'b11100010_10110000_10010010_1;
      patterns[58035] = 25'b11100010_10110001_10010011_1;
      patterns[58036] = 25'b11100010_10110010_10010100_1;
      patterns[58037] = 25'b11100010_10110011_10010101_1;
      patterns[58038] = 25'b11100010_10110100_10010110_1;
      patterns[58039] = 25'b11100010_10110101_10010111_1;
      patterns[58040] = 25'b11100010_10110110_10011000_1;
      patterns[58041] = 25'b11100010_10110111_10011001_1;
      patterns[58042] = 25'b11100010_10111000_10011010_1;
      patterns[58043] = 25'b11100010_10111001_10011011_1;
      patterns[58044] = 25'b11100010_10111010_10011100_1;
      patterns[58045] = 25'b11100010_10111011_10011101_1;
      patterns[58046] = 25'b11100010_10111100_10011110_1;
      patterns[58047] = 25'b11100010_10111101_10011111_1;
      patterns[58048] = 25'b11100010_10111110_10100000_1;
      patterns[58049] = 25'b11100010_10111111_10100001_1;
      patterns[58050] = 25'b11100010_11000000_10100010_1;
      patterns[58051] = 25'b11100010_11000001_10100011_1;
      patterns[58052] = 25'b11100010_11000010_10100100_1;
      patterns[58053] = 25'b11100010_11000011_10100101_1;
      patterns[58054] = 25'b11100010_11000100_10100110_1;
      patterns[58055] = 25'b11100010_11000101_10100111_1;
      patterns[58056] = 25'b11100010_11000110_10101000_1;
      patterns[58057] = 25'b11100010_11000111_10101001_1;
      patterns[58058] = 25'b11100010_11001000_10101010_1;
      patterns[58059] = 25'b11100010_11001001_10101011_1;
      patterns[58060] = 25'b11100010_11001010_10101100_1;
      patterns[58061] = 25'b11100010_11001011_10101101_1;
      patterns[58062] = 25'b11100010_11001100_10101110_1;
      patterns[58063] = 25'b11100010_11001101_10101111_1;
      patterns[58064] = 25'b11100010_11001110_10110000_1;
      patterns[58065] = 25'b11100010_11001111_10110001_1;
      patterns[58066] = 25'b11100010_11010000_10110010_1;
      patterns[58067] = 25'b11100010_11010001_10110011_1;
      patterns[58068] = 25'b11100010_11010010_10110100_1;
      patterns[58069] = 25'b11100010_11010011_10110101_1;
      patterns[58070] = 25'b11100010_11010100_10110110_1;
      patterns[58071] = 25'b11100010_11010101_10110111_1;
      patterns[58072] = 25'b11100010_11010110_10111000_1;
      patterns[58073] = 25'b11100010_11010111_10111001_1;
      patterns[58074] = 25'b11100010_11011000_10111010_1;
      patterns[58075] = 25'b11100010_11011001_10111011_1;
      patterns[58076] = 25'b11100010_11011010_10111100_1;
      patterns[58077] = 25'b11100010_11011011_10111101_1;
      patterns[58078] = 25'b11100010_11011100_10111110_1;
      patterns[58079] = 25'b11100010_11011101_10111111_1;
      patterns[58080] = 25'b11100010_11011110_11000000_1;
      patterns[58081] = 25'b11100010_11011111_11000001_1;
      patterns[58082] = 25'b11100010_11100000_11000010_1;
      patterns[58083] = 25'b11100010_11100001_11000011_1;
      patterns[58084] = 25'b11100010_11100010_11000100_1;
      patterns[58085] = 25'b11100010_11100011_11000101_1;
      patterns[58086] = 25'b11100010_11100100_11000110_1;
      patterns[58087] = 25'b11100010_11100101_11000111_1;
      patterns[58088] = 25'b11100010_11100110_11001000_1;
      patterns[58089] = 25'b11100010_11100111_11001001_1;
      patterns[58090] = 25'b11100010_11101000_11001010_1;
      patterns[58091] = 25'b11100010_11101001_11001011_1;
      patterns[58092] = 25'b11100010_11101010_11001100_1;
      patterns[58093] = 25'b11100010_11101011_11001101_1;
      patterns[58094] = 25'b11100010_11101100_11001110_1;
      patterns[58095] = 25'b11100010_11101101_11001111_1;
      patterns[58096] = 25'b11100010_11101110_11010000_1;
      patterns[58097] = 25'b11100010_11101111_11010001_1;
      patterns[58098] = 25'b11100010_11110000_11010010_1;
      patterns[58099] = 25'b11100010_11110001_11010011_1;
      patterns[58100] = 25'b11100010_11110010_11010100_1;
      patterns[58101] = 25'b11100010_11110011_11010101_1;
      patterns[58102] = 25'b11100010_11110100_11010110_1;
      patterns[58103] = 25'b11100010_11110101_11010111_1;
      patterns[58104] = 25'b11100010_11110110_11011000_1;
      patterns[58105] = 25'b11100010_11110111_11011001_1;
      patterns[58106] = 25'b11100010_11111000_11011010_1;
      patterns[58107] = 25'b11100010_11111001_11011011_1;
      patterns[58108] = 25'b11100010_11111010_11011100_1;
      patterns[58109] = 25'b11100010_11111011_11011101_1;
      patterns[58110] = 25'b11100010_11111100_11011110_1;
      patterns[58111] = 25'b11100010_11111101_11011111_1;
      patterns[58112] = 25'b11100010_11111110_11100000_1;
      patterns[58113] = 25'b11100010_11111111_11100001_1;
      patterns[58114] = 25'b11100011_00000000_11100011_0;
      patterns[58115] = 25'b11100011_00000001_11100100_0;
      patterns[58116] = 25'b11100011_00000010_11100101_0;
      patterns[58117] = 25'b11100011_00000011_11100110_0;
      patterns[58118] = 25'b11100011_00000100_11100111_0;
      patterns[58119] = 25'b11100011_00000101_11101000_0;
      patterns[58120] = 25'b11100011_00000110_11101001_0;
      patterns[58121] = 25'b11100011_00000111_11101010_0;
      patterns[58122] = 25'b11100011_00001000_11101011_0;
      patterns[58123] = 25'b11100011_00001001_11101100_0;
      patterns[58124] = 25'b11100011_00001010_11101101_0;
      patterns[58125] = 25'b11100011_00001011_11101110_0;
      patterns[58126] = 25'b11100011_00001100_11101111_0;
      patterns[58127] = 25'b11100011_00001101_11110000_0;
      patterns[58128] = 25'b11100011_00001110_11110001_0;
      patterns[58129] = 25'b11100011_00001111_11110010_0;
      patterns[58130] = 25'b11100011_00010000_11110011_0;
      patterns[58131] = 25'b11100011_00010001_11110100_0;
      patterns[58132] = 25'b11100011_00010010_11110101_0;
      patterns[58133] = 25'b11100011_00010011_11110110_0;
      patterns[58134] = 25'b11100011_00010100_11110111_0;
      patterns[58135] = 25'b11100011_00010101_11111000_0;
      patterns[58136] = 25'b11100011_00010110_11111001_0;
      patterns[58137] = 25'b11100011_00010111_11111010_0;
      patterns[58138] = 25'b11100011_00011000_11111011_0;
      patterns[58139] = 25'b11100011_00011001_11111100_0;
      patterns[58140] = 25'b11100011_00011010_11111101_0;
      patterns[58141] = 25'b11100011_00011011_11111110_0;
      patterns[58142] = 25'b11100011_00011100_11111111_0;
      patterns[58143] = 25'b11100011_00011101_00000000_1;
      patterns[58144] = 25'b11100011_00011110_00000001_1;
      patterns[58145] = 25'b11100011_00011111_00000010_1;
      patterns[58146] = 25'b11100011_00100000_00000011_1;
      patterns[58147] = 25'b11100011_00100001_00000100_1;
      patterns[58148] = 25'b11100011_00100010_00000101_1;
      patterns[58149] = 25'b11100011_00100011_00000110_1;
      patterns[58150] = 25'b11100011_00100100_00000111_1;
      patterns[58151] = 25'b11100011_00100101_00001000_1;
      patterns[58152] = 25'b11100011_00100110_00001001_1;
      patterns[58153] = 25'b11100011_00100111_00001010_1;
      patterns[58154] = 25'b11100011_00101000_00001011_1;
      patterns[58155] = 25'b11100011_00101001_00001100_1;
      patterns[58156] = 25'b11100011_00101010_00001101_1;
      patterns[58157] = 25'b11100011_00101011_00001110_1;
      patterns[58158] = 25'b11100011_00101100_00001111_1;
      patterns[58159] = 25'b11100011_00101101_00010000_1;
      patterns[58160] = 25'b11100011_00101110_00010001_1;
      patterns[58161] = 25'b11100011_00101111_00010010_1;
      patterns[58162] = 25'b11100011_00110000_00010011_1;
      patterns[58163] = 25'b11100011_00110001_00010100_1;
      patterns[58164] = 25'b11100011_00110010_00010101_1;
      patterns[58165] = 25'b11100011_00110011_00010110_1;
      patterns[58166] = 25'b11100011_00110100_00010111_1;
      patterns[58167] = 25'b11100011_00110101_00011000_1;
      patterns[58168] = 25'b11100011_00110110_00011001_1;
      patterns[58169] = 25'b11100011_00110111_00011010_1;
      patterns[58170] = 25'b11100011_00111000_00011011_1;
      patterns[58171] = 25'b11100011_00111001_00011100_1;
      patterns[58172] = 25'b11100011_00111010_00011101_1;
      patterns[58173] = 25'b11100011_00111011_00011110_1;
      patterns[58174] = 25'b11100011_00111100_00011111_1;
      patterns[58175] = 25'b11100011_00111101_00100000_1;
      patterns[58176] = 25'b11100011_00111110_00100001_1;
      patterns[58177] = 25'b11100011_00111111_00100010_1;
      patterns[58178] = 25'b11100011_01000000_00100011_1;
      patterns[58179] = 25'b11100011_01000001_00100100_1;
      patterns[58180] = 25'b11100011_01000010_00100101_1;
      patterns[58181] = 25'b11100011_01000011_00100110_1;
      patterns[58182] = 25'b11100011_01000100_00100111_1;
      patterns[58183] = 25'b11100011_01000101_00101000_1;
      patterns[58184] = 25'b11100011_01000110_00101001_1;
      patterns[58185] = 25'b11100011_01000111_00101010_1;
      patterns[58186] = 25'b11100011_01001000_00101011_1;
      patterns[58187] = 25'b11100011_01001001_00101100_1;
      patterns[58188] = 25'b11100011_01001010_00101101_1;
      patterns[58189] = 25'b11100011_01001011_00101110_1;
      patterns[58190] = 25'b11100011_01001100_00101111_1;
      patterns[58191] = 25'b11100011_01001101_00110000_1;
      patterns[58192] = 25'b11100011_01001110_00110001_1;
      patterns[58193] = 25'b11100011_01001111_00110010_1;
      patterns[58194] = 25'b11100011_01010000_00110011_1;
      patterns[58195] = 25'b11100011_01010001_00110100_1;
      patterns[58196] = 25'b11100011_01010010_00110101_1;
      patterns[58197] = 25'b11100011_01010011_00110110_1;
      patterns[58198] = 25'b11100011_01010100_00110111_1;
      patterns[58199] = 25'b11100011_01010101_00111000_1;
      patterns[58200] = 25'b11100011_01010110_00111001_1;
      patterns[58201] = 25'b11100011_01010111_00111010_1;
      patterns[58202] = 25'b11100011_01011000_00111011_1;
      patterns[58203] = 25'b11100011_01011001_00111100_1;
      patterns[58204] = 25'b11100011_01011010_00111101_1;
      patterns[58205] = 25'b11100011_01011011_00111110_1;
      patterns[58206] = 25'b11100011_01011100_00111111_1;
      patterns[58207] = 25'b11100011_01011101_01000000_1;
      patterns[58208] = 25'b11100011_01011110_01000001_1;
      patterns[58209] = 25'b11100011_01011111_01000010_1;
      patterns[58210] = 25'b11100011_01100000_01000011_1;
      patterns[58211] = 25'b11100011_01100001_01000100_1;
      patterns[58212] = 25'b11100011_01100010_01000101_1;
      patterns[58213] = 25'b11100011_01100011_01000110_1;
      patterns[58214] = 25'b11100011_01100100_01000111_1;
      patterns[58215] = 25'b11100011_01100101_01001000_1;
      patterns[58216] = 25'b11100011_01100110_01001001_1;
      patterns[58217] = 25'b11100011_01100111_01001010_1;
      patterns[58218] = 25'b11100011_01101000_01001011_1;
      patterns[58219] = 25'b11100011_01101001_01001100_1;
      patterns[58220] = 25'b11100011_01101010_01001101_1;
      patterns[58221] = 25'b11100011_01101011_01001110_1;
      patterns[58222] = 25'b11100011_01101100_01001111_1;
      patterns[58223] = 25'b11100011_01101101_01010000_1;
      patterns[58224] = 25'b11100011_01101110_01010001_1;
      patterns[58225] = 25'b11100011_01101111_01010010_1;
      patterns[58226] = 25'b11100011_01110000_01010011_1;
      patterns[58227] = 25'b11100011_01110001_01010100_1;
      patterns[58228] = 25'b11100011_01110010_01010101_1;
      patterns[58229] = 25'b11100011_01110011_01010110_1;
      patterns[58230] = 25'b11100011_01110100_01010111_1;
      patterns[58231] = 25'b11100011_01110101_01011000_1;
      patterns[58232] = 25'b11100011_01110110_01011001_1;
      patterns[58233] = 25'b11100011_01110111_01011010_1;
      patterns[58234] = 25'b11100011_01111000_01011011_1;
      patterns[58235] = 25'b11100011_01111001_01011100_1;
      patterns[58236] = 25'b11100011_01111010_01011101_1;
      patterns[58237] = 25'b11100011_01111011_01011110_1;
      patterns[58238] = 25'b11100011_01111100_01011111_1;
      patterns[58239] = 25'b11100011_01111101_01100000_1;
      patterns[58240] = 25'b11100011_01111110_01100001_1;
      patterns[58241] = 25'b11100011_01111111_01100010_1;
      patterns[58242] = 25'b11100011_10000000_01100011_1;
      patterns[58243] = 25'b11100011_10000001_01100100_1;
      patterns[58244] = 25'b11100011_10000010_01100101_1;
      patterns[58245] = 25'b11100011_10000011_01100110_1;
      patterns[58246] = 25'b11100011_10000100_01100111_1;
      patterns[58247] = 25'b11100011_10000101_01101000_1;
      patterns[58248] = 25'b11100011_10000110_01101001_1;
      patterns[58249] = 25'b11100011_10000111_01101010_1;
      patterns[58250] = 25'b11100011_10001000_01101011_1;
      patterns[58251] = 25'b11100011_10001001_01101100_1;
      patterns[58252] = 25'b11100011_10001010_01101101_1;
      patterns[58253] = 25'b11100011_10001011_01101110_1;
      patterns[58254] = 25'b11100011_10001100_01101111_1;
      patterns[58255] = 25'b11100011_10001101_01110000_1;
      patterns[58256] = 25'b11100011_10001110_01110001_1;
      patterns[58257] = 25'b11100011_10001111_01110010_1;
      patterns[58258] = 25'b11100011_10010000_01110011_1;
      patterns[58259] = 25'b11100011_10010001_01110100_1;
      patterns[58260] = 25'b11100011_10010010_01110101_1;
      patterns[58261] = 25'b11100011_10010011_01110110_1;
      patterns[58262] = 25'b11100011_10010100_01110111_1;
      patterns[58263] = 25'b11100011_10010101_01111000_1;
      patterns[58264] = 25'b11100011_10010110_01111001_1;
      patterns[58265] = 25'b11100011_10010111_01111010_1;
      patterns[58266] = 25'b11100011_10011000_01111011_1;
      patterns[58267] = 25'b11100011_10011001_01111100_1;
      patterns[58268] = 25'b11100011_10011010_01111101_1;
      patterns[58269] = 25'b11100011_10011011_01111110_1;
      patterns[58270] = 25'b11100011_10011100_01111111_1;
      patterns[58271] = 25'b11100011_10011101_10000000_1;
      patterns[58272] = 25'b11100011_10011110_10000001_1;
      patterns[58273] = 25'b11100011_10011111_10000010_1;
      patterns[58274] = 25'b11100011_10100000_10000011_1;
      patterns[58275] = 25'b11100011_10100001_10000100_1;
      patterns[58276] = 25'b11100011_10100010_10000101_1;
      patterns[58277] = 25'b11100011_10100011_10000110_1;
      patterns[58278] = 25'b11100011_10100100_10000111_1;
      patterns[58279] = 25'b11100011_10100101_10001000_1;
      patterns[58280] = 25'b11100011_10100110_10001001_1;
      patterns[58281] = 25'b11100011_10100111_10001010_1;
      patterns[58282] = 25'b11100011_10101000_10001011_1;
      patterns[58283] = 25'b11100011_10101001_10001100_1;
      patterns[58284] = 25'b11100011_10101010_10001101_1;
      patterns[58285] = 25'b11100011_10101011_10001110_1;
      patterns[58286] = 25'b11100011_10101100_10001111_1;
      patterns[58287] = 25'b11100011_10101101_10010000_1;
      patterns[58288] = 25'b11100011_10101110_10010001_1;
      patterns[58289] = 25'b11100011_10101111_10010010_1;
      patterns[58290] = 25'b11100011_10110000_10010011_1;
      patterns[58291] = 25'b11100011_10110001_10010100_1;
      patterns[58292] = 25'b11100011_10110010_10010101_1;
      patterns[58293] = 25'b11100011_10110011_10010110_1;
      patterns[58294] = 25'b11100011_10110100_10010111_1;
      patterns[58295] = 25'b11100011_10110101_10011000_1;
      patterns[58296] = 25'b11100011_10110110_10011001_1;
      patterns[58297] = 25'b11100011_10110111_10011010_1;
      patterns[58298] = 25'b11100011_10111000_10011011_1;
      patterns[58299] = 25'b11100011_10111001_10011100_1;
      patterns[58300] = 25'b11100011_10111010_10011101_1;
      patterns[58301] = 25'b11100011_10111011_10011110_1;
      patterns[58302] = 25'b11100011_10111100_10011111_1;
      patterns[58303] = 25'b11100011_10111101_10100000_1;
      patterns[58304] = 25'b11100011_10111110_10100001_1;
      patterns[58305] = 25'b11100011_10111111_10100010_1;
      patterns[58306] = 25'b11100011_11000000_10100011_1;
      patterns[58307] = 25'b11100011_11000001_10100100_1;
      patterns[58308] = 25'b11100011_11000010_10100101_1;
      patterns[58309] = 25'b11100011_11000011_10100110_1;
      patterns[58310] = 25'b11100011_11000100_10100111_1;
      patterns[58311] = 25'b11100011_11000101_10101000_1;
      patterns[58312] = 25'b11100011_11000110_10101001_1;
      patterns[58313] = 25'b11100011_11000111_10101010_1;
      patterns[58314] = 25'b11100011_11001000_10101011_1;
      patterns[58315] = 25'b11100011_11001001_10101100_1;
      patterns[58316] = 25'b11100011_11001010_10101101_1;
      patterns[58317] = 25'b11100011_11001011_10101110_1;
      patterns[58318] = 25'b11100011_11001100_10101111_1;
      patterns[58319] = 25'b11100011_11001101_10110000_1;
      patterns[58320] = 25'b11100011_11001110_10110001_1;
      patterns[58321] = 25'b11100011_11001111_10110010_1;
      patterns[58322] = 25'b11100011_11010000_10110011_1;
      patterns[58323] = 25'b11100011_11010001_10110100_1;
      patterns[58324] = 25'b11100011_11010010_10110101_1;
      patterns[58325] = 25'b11100011_11010011_10110110_1;
      patterns[58326] = 25'b11100011_11010100_10110111_1;
      patterns[58327] = 25'b11100011_11010101_10111000_1;
      patterns[58328] = 25'b11100011_11010110_10111001_1;
      patterns[58329] = 25'b11100011_11010111_10111010_1;
      patterns[58330] = 25'b11100011_11011000_10111011_1;
      patterns[58331] = 25'b11100011_11011001_10111100_1;
      patterns[58332] = 25'b11100011_11011010_10111101_1;
      patterns[58333] = 25'b11100011_11011011_10111110_1;
      patterns[58334] = 25'b11100011_11011100_10111111_1;
      patterns[58335] = 25'b11100011_11011101_11000000_1;
      patterns[58336] = 25'b11100011_11011110_11000001_1;
      patterns[58337] = 25'b11100011_11011111_11000010_1;
      patterns[58338] = 25'b11100011_11100000_11000011_1;
      patterns[58339] = 25'b11100011_11100001_11000100_1;
      patterns[58340] = 25'b11100011_11100010_11000101_1;
      patterns[58341] = 25'b11100011_11100011_11000110_1;
      patterns[58342] = 25'b11100011_11100100_11000111_1;
      patterns[58343] = 25'b11100011_11100101_11001000_1;
      patterns[58344] = 25'b11100011_11100110_11001001_1;
      patterns[58345] = 25'b11100011_11100111_11001010_1;
      patterns[58346] = 25'b11100011_11101000_11001011_1;
      patterns[58347] = 25'b11100011_11101001_11001100_1;
      patterns[58348] = 25'b11100011_11101010_11001101_1;
      patterns[58349] = 25'b11100011_11101011_11001110_1;
      patterns[58350] = 25'b11100011_11101100_11001111_1;
      patterns[58351] = 25'b11100011_11101101_11010000_1;
      patterns[58352] = 25'b11100011_11101110_11010001_1;
      patterns[58353] = 25'b11100011_11101111_11010010_1;
      patterns[58354] = 25'b11100011_11110000_11010011_1;
      patterns[58355] = 25'b11100011_11110001_11010100_1;
      patterns[58356] = 25'b11100011_11110010_11010101_1;
      patterns[58357] = 25'b11100011_11110011_11010110_1;
      patterns[58358] = 25'b11100011_11110100_11010111_1;
      patterns[58359] = 25'b11100011_11110101_11011000_1;
      patterns[58360] = 25'b11100011_11110110_11011001_1;
      patterns[58361] = 25'b11100011_11110111_11011010_1;
      patterns[58362] = 25'b11100011_11111000_11011011_1;
      patterns[58363] = 25'b11100011_11111001_11011100_1;
      patterns[58364] = 25'b11100011_11111010_11011101_1;
      patterns[58365] = 25'b11100011_11111011_11011110_1;
      patterns[58366] = 25'b11100011_11111100_11011111_1;
      patterns[58367] = 25'b11100011_11111101_11100000_1;
      patterns[58368] = 25'b11100011_11111110_11100001_1;
      patterns[58369] = 25'b11100011_11111111_11100010_1;
      patterns[58370] = 25'b11100100_00000000_11100100_0;
      patterns[58371] = 25'b11100100_00000001_11100101_0;
      patterns[58372] = 25'b11100100_00000010_11100110_0;
      patterns[58373] = 25'b11100100_00000011_11100111_0;
      patterns[58374] = 25'b11100100_00000100_11101000_0;
      patterns[58375] = 25'b11100100_00000101_11101001_0;
      patterns[58376] = 25'b11100100_00000110_11101010_0;
      patterns[58377] = 25'b11100100_00000111_11101011_0;
      patterns[58378] = 25'b11100100_00001000_11101100_0;
      patterns[58379] = 25'b11100100_00001001_11101101_0;
      patterns[58380] = 25'b11100100_00001010_11101110_0;
      patterns[58381] = 25'b11100100_00001011_11101111_0;
      patterns[58382] = 25'b11100100_00001100_11110000_0;
      patterns[58383] = 25'b11100100_00001101_11110001_0;
      patterns[58384] = 25'b11100100_00001110_11110010_0;
      patterns[58385] = 25'b11100100_00001111_11110011_0;
      patterns[58386] = 25'b11100100_00010000_11110100_0;
      patterns[58387] = 25'b11100100_00010001_11110101_0;
      patterns[58388] = 25'b11100100_00010010_11110110_0;
      patterns[58389] = 25'b11100100_00010011_11110111_0;
      patterns[58390] = 25'b11100100_00010100_11111000_0;
      patterns[58391] = 25'b11100100_00010101_11111001_0;
      patterns[58392] = 25'b11100100_00010110_11111010_0;
      patterns[58393] = 25'b11100100_00010111_11111011_0;
      patterns[58394] = 25'b11100100_00011000_11111100_0;
      patterns[58395] = 25'b11100100_00011001_11111101_0;
      patterns[58396] = 25'b11100100_00011010_11111110_0;
      patterns[58397] = 25'b11100100_00011011_11111111_0;
      patterns[58398] = 25'b11100100_00011100_00000000_1;
      patterns[58399] = 25'b11100100_00011101_00000001_1;
      patterns[58400] = 25'b11100100_00011110_00000010_1;
      patterns[58401] = 25'b11100100_00011111_00000011_1;
      patterns[58402] = 25'b11100100_00100000_00000100_1;
      patterns[58403] = 25'b11100100_00100001_00000101_1;
      patterns[58404] = 25'b11100100_00100010_00000110_1;
      patterns[58405] = 25'b11100100_00100011_00000111_1;
      patterns[58406] = 25'b11100100_00100100_00001000_1;
      patterns[58407] = 25'b11100100_00100101_00001001_1;
      patterns[58408] = 25'b11100100_00100110_00001010_1;
      patterns[58409] = 25'b11100100_00100111_00001011_1;
      patterns[58410] = 25'b11100100_00101000_00001100_1;
      patterns[58411] = 25'b11100100_00101001_00001101_1;
      patterns[58412] = 25'b11100100_00101010_00001110_1;
      patterns[58413] = 25'b11100100_00101011_00001111_1;
      patterns[58414] = 25'b11100100_00101100_00010000_1;
      patterns[58415] = 25'b11100100_00101101_00010001_1;
      patterns[58416] = 25'b11100100_00101110_00010010_1;
      patterns[58417] = 25'b11100100_00101111_00010011_1;
      patterns[58418] = 25'b11100100_00110000_00010100_1;
      patterns[58419] = 25'b11100100_00110001_00010101_1;
      patterns[58420] = 25'b11100100_00110010_00010110_1;
      patterns[58421] = 25'b11100100_00110011_00010111_1;
      patterns[58422] = 25'b11100100_00110100_00011000_1;
      patterns[58423] = 25'b11100100_00110101_00011001_1;
      patterns[58424] = 25'b11100100_00110110_00011010_1;
      patterns[58425] = 25'b11100100_00110111_00011011_1;
      patterns[58426] = 25'b11100100_00111000_00011100_1;
      patterns[58427] = 25'b11100100_00111001_00011101_1;
      patterns[58428] = 25'b11100100_00111010_00011110_1;
      patterns[58429] = 25'b11100100_00111011_00011111_1;
      patterns[58430] = 25'b11100100_00111100_00100000_1;
      patterns[58431] = 25'b11100100_00111101_00100001_1;
      patterns[58432] = 25'b11100100_00111110_00100010_1;
      patterns[58433] = 25'b11100100_00111111_00100011_1;
      patterns[58434] = 25'b11100100_01000000_00100100_1;
      patterns[58435] = 25'b11100100_01000001_00100101_1;
      patterns[58436] = 25'b11100100_01000010_00100110_1;
      patterns[58437] = 25'b11100100_01000011_00100111_1;
      patterns[58438] = 25'b11100100_01000100_00101000_1;
      patterns[58439] = 25'b11100100_01000101_00101001_1;
      patterns[58440] = 25'b11100100_01000110_00101010_1;
      patterns[58441] = 25'b11100100_01000111_00101011_1;
      patterns[58442] = 25'b11100100_01001000_00101100_1;
      patterns[58443] = 25'b11100100_01001001_00101101_1;
      patterns[58444] = 25'b11100100_01001010_00101110_1;
      patterns[58445] = 25'b11100100_01001011_00101111_1;
      patterns[58446] = 25'b11100100_01001100_00110000_1;
      patterns[58447] = 25'b11100100_01001101_00110001_1;
      patterns[58448] = 25'b11100100_01001110_00110010_1;
      patterns[58449] = 25'b11100100_01001111_00110011_1;
      patterns[58450] = 25'b11100100_01010000_00110100_1;
      patterns[58451] = 25'b11100100_01010001_00110101_1;
      patterns[58452] = 25'b11100100_01010010_00110110_1;
      patterns[58453] = 25'b11100100_01010011_00110111_1;
      patterns[58454] = 25'b11100100_01010100_00111000_1;
      patterns[58455] = 25'b11100100_01010101_00111001_1;
      patterns[58456] = 25'b11100100_01010110_00111010_1;
      patterns[58457] = 25'b11100100_01010111_00111011_1;
      patterns[58458] = 25'b11100100_01011000_00111100_1;
      patterns[58459] = 25'b11100100_01011001_00111101_1;
      patterns[58460] = 25'b11100100_01011010_00111110_1;
      patterns[58461] = 25'b11100100_01011011_00111111_1;
      patterns[58462] = 25'b11100100_01011100_01000000_1;
      patterns[58463] = 25'b11100100_01011101_01000001_1;
      patterns[58464] = 25'b11100100_01011110_01000010_1;
      patterns[58465] = 25'b11100100_01011111_01000011_1;
      patterns[58466] = 25'b11100100_01100000_01000100_1;
      patterns[58467] = 25'b11100100_01100001_01000101_1;
      patterns[58468] = 25'b11100100_01100010_01000110_1;
      patterns[58469] = 25'b11100100_01100011_01000111_1;
      patterns[58470] = 25'b11100100_01100100_01001000_1;
      patterns[58471] = 25'b11100100_01100101_01001001_1;
      patterns[58472] = 25'b11100100_01100110_01001010_1;
      patterns[58473] = 25'b11100100_01100111_01001011_1;
      patterns[58474] = 25'b11100100_01101000_01001100_1;
      patterns[58475] = 25'b11100100_01101001_01001101_1;
      patterns[58476] = 25'b11100100_01101010_01001110_1;
      patterns[58477] = 25'b11100100_01101011_01001111_1;
      patterns[58478] = 25'b11100100_01101100_01010000_1;
      patterns[58479] = 25'b11100100_01101101_01010001_1;
      patterns[58480] = 25'b11100100_01101110_01010010_1;
      patterns[58481] = 25'b11100100_01101111_01010011_1;
      patterns[58482] = 25'b11100100_01110000_01010100_1;
      patterns[58483] = 25'b11100100_01110001_01010101_1;
      patterns[58484] = 25'b11100100_01110010_01010110_1;
      patterns[58485] = 25'b11100100_01110011_01010111_1;
      patterns[58486] = 25'b11100100_01110100_01011000_1;
      patterns[58487] = 25'b11100100_01110101_01011001_1;
      patterns[58488] = 25'b11100100_01110110_01011010_1;
      patterns[58489] = 25'b11100100_01110111_01011011_1;
      patterns[58490] = 25'b11100100_01111000_01011100_1;
      patterns[58491] = 25'b11100100_01111001_01011101_1;
      patterns[58492] = 25'b11100100_01111010_01011110_1;
      patterns[58493] = 25'b11100100_01111011_01011111_1;
      patterns[58494] = 25'b11100100_01111100_01100000_1;
      patterns[58495] = 25'b11100100_01111101_01100001_1;
      patterns[58496] = 25'b11100100_01111110_01100010_1;
      patterns[58497] = 25'b11100100_01111111_01100011_1;
      patterns[58498] = 25'b11100100_10000000_01100100_1;
      patterns[58499] = 25'b11100100_10000001_01100101_1;
      patterns[58500] = 25'b11100100_10000010_01100110_1;
      patterns[58501] = 25'b11100100_10000011_01100111_1;
      patterns[58502] = 25'b11100100_10000100_01101000_1;
      patterns[58503] = 25'b11100100_10000101_01101001_1;
      patterns[58504] = 25'b11100100_10000110_01101010_1;
      patterns[58505] = 25'b11100100_10000111_01101011_1;
      patterns[58506] = 25'b11100100_10001000_01101100_1;
      patterns[58507] = 25'b11100100_10001001_01101101_1;
      patterns[58508] = 25'b11100100_10001010_01101110_1;
      patterns[58509] = 25'b11100100_10001011_01101111_1;
      patterns[58510] = 25'b11100100_10001100_01110000_1;
      patterns[58511] = 25'b11100100_10001101_01110001_1;
      patterns[58512] = 25'b11100100_10001110_01110010_1;
      patterns[58513] = 25'b11100100_10001111_01110011_1;
      patterns[58514] = 25'b11100100_10010000_01110100_1;
      patterns[58515] = 25'b11100100_10010001_01110101_1;
      patterns[58516] = 25'b11100100_10010010_01110110_1;
      patterns[58517] = 25'b11100100_10010011_01110111_1;
      patterns[58518] = 25'b11100100_10010100_01111000_1;
      patterns[58519] = 25'b11100100_10010101_01111001_1;
      patterns[58520] = 25'b11100100_10010110_01111010_1;
      patterns[58521] = 25'b11100100_10010111_01111011_1;
      patterns[58522] = 25'b11100100_10011000_01111100_1;
      patterns[58523] = 25'b11100100_10011001_01111101_1;
      patterns[58524] = 25'b11100100_10011010_01111110_1;
      patterns[58525] = 25'b11100100_10011011_01111111_1;
      patterns[58526] = 25'b11100100_10011100_10000000_1;
      patterns[58527] = 25'b11100100_10011101_10000001_1;
      patterns[58528] = 25'b11100100_10011110_10000010_1;
      patterns[58529] = 25'b11100100_10011111_10000011_1;
      patterns[58530] = 25'b11100100_10100000_10000100_1;
      patterns[58531] = 25'b11100100_10100001_10000101_1;
      patterns[58532] = 25'b11100100_10100010_10000110_1;
      patterns[58533] = 25'b11100100_10100011_10000111_1;
      patterns[58534] = 25'b11100100_10100100_10001000_1;
      patterns[58535] = 25'b11100100_10100101_10001001_1;
      patterns[58536] = 25'b11100100_10100110_10001010_1;
      patterns[58537] = 25'b11100100_10100111_10001011_1;
      patterns[58538] = 25'b11100100_10101000_10001100_1;
      patterns[58539] = 25'b11100100_10101001_10001101_1;
      patterns[58540] = 25'b11100100_10101010_10001110_1;
      patterns[58541] = 25'b11100100_10101011_10001111_1;
      patterns[58542] = 25'b11100100_10101100_10010000_1;
      patterns[58543] = 25'b11100100_10101101_10010001_1;
      patterns[58544] = 25'b11100100_10101110_10010010_1;
      patterns[58545] = 25'b11100100_10101111_10010011_1;
      patterns[58546] = 25'b11100100_10110000_10010100_1;
      patterns[58547] = 25'b11100100_10110001_10010101_1;
      patterns[58548] = 25'b11100100_10110010_10010110_1;
      patterns[58549] = 25'b11100100_10110011_10010111_1;
      patterns[58550] = 25'b11100100_10110100_10011000_1;
      patterns[58551] = 25'b11100100_10110101_10011001_1;
      patterns[58552] = 25'b11100100_10110110_10011010_1;
      patterns[58553] = 25'b11100100_10110111_10011011_1;
      patterns[58554] = 25'b11100100_10111000_10011100_1;
      patterns[58555] = 25'b11100100_10111001_10011101_1;
      patterns[58556] = 25'b11100100_10111010_10011110_1;
      patterns[58557] = 25'b11100100_10111011_10011111_1;
      patterns[58558] = 25'b11100100_10111100_10100000_1;
      patterns[58559] = 25'b11100100_10111101_10100001_1;
      patterns[58560] = 25'b11100100_10111110_10100010_1;
      patterns[58561] = 25'b11100100_10111111_10100011_1;
      patterns[58562] = 25'b11100100_11000000_10100100_1;
      patterns[58563] = 25'b11100100_11000001_10100101_1;
      patterns[58564] = 25'b11100100_11000010_10100110_1;
      patterns[58565] = 25'b11100100_11000011_10100111_1;
      patterns[58566] = 25'b11100100_11000100_10101000_1;
      patterns[58567] = 25'b11100100_11000101_10101001_1;
      patterns[58568] = 25'b11100100_11000110_10101010_1;
      patterns[58569] = 25'b11100100_11000111_10101011_1;
      patterns[58570] = 25'b11100100_11001000_10101100_1;
      patterns[58571] = 25'b11100100_11001001_10101101_1;
      patterns[58572] = 25'b11100100_11001010_10101110_1;
      patterns[58573] = 25'b11100100_11001011_10101111_1;
      patterns[58574] = 25'b11100100_11001100_10110000_1;
      patterns[58575] = 25'b11100100_11001101_10110001_1;
      patterns[58576] = 25'b11100100_11001110_10110010_1;
      patterns[58577] = 25'b11100100_11001111_10110011_1;
      patterns[58578] = 25'b11100100_11010000_10110100_1;
      patterns[58579] = 25'b11100100_11010001_10110101_1;
      patterns[58580] = 25'b11100100_11010010_10110110_1;
      patterns[58581] = 25'b11100100_11010011_10110111_1;
      patterns[58582] = 25'b11100100_11010100_10111000_1;
      patterns[58583] = 25'b11100100_11010101_10111001_1;
      patterns[58584] = 25'b11100100_11010110_10111010_1;
      patterns[58585] = 25'b11100100_11010111_10111011_1;
      patterns[58586] = 25'b11100100_11011000_10111100_1;
      patterns[58587] = 25'b11100100_11011001_10111101_1;
      patterns[58588] = 25'b11100100_11011010_10111110_1;
      patterns[58589] = 25'b11100100_11011011_10111111_1;
      patterns[58590] = 25'b11100100_11011100_11000000_1;
      patterns[58591] = 25'b11100100_11011101_11000001_1;
      patterns[58592] = 25'b11100100_11011110_11000010_1;
      patterns[58593] = 25'b11100100_11011111_11000011_1;
      patterns[58594] = 25'b11100100_11100000_11000100_1;
      patterns[58595] = 25'b11100100_11100001_11000101_1;
      patterns[58596] = 25'b11100100_11100010_11000110_1;
      patterns[58597] = 25'b11100100_11100011_11000111_1;
      patterns[58598] = 25'b11100100_11100100_11001000_1;
      patterns[58599] = 25'b11100100_11100101_11001001_1;
      patterns[58600] = 25'b11100100_11100110_11001010_1;
      patterns[58601] = 25'b11100100_11100111_11001011_1;
      patterns[58602] = 25'b11100100_11101000_11001100_1;
      patterns[58603] = 25'b11100100_11101001_11001101_1;
      patterns[58604] = 25'b11100100_11101010_11001110_1;
      patterns[58605] = 25'b11100100_11101011_11001111_1;
      patterns[58606] = 25'b11100100_11101100_11010000_1;
      patterns[58607] = 25'b11100100_11101101_11010001_1;
      patterns[58608] = 25'b11100100_11101110_11010010_1;
      patterns[58609] = 25'b11100100_11101111_11010011_1;
      patterns[58610] = 25'b11100100_11110000_11010100_1;
      patterns[58611] = 25'b11100100_11110001_11010101_1;
      patterns[58612] = 25'b11100100_11110010_11010110_1;
      patterns[58613] = 25'b11100100_11110011_11010111_1;
      patterns[58614] = 25'b11100100_11110100_11011000_1;
      patterns[58615] = 25'b11100100_11110101_11011001_1;
      patterns[58616] = 25'b11100100_11110110_11011010_1;
      patterns[58617] = 25'b11100100_11110111_11011011_1;
      patterns[58618] = 25'b11100100_11111000_11011100_1;
      patterns[58619] = 25'b11100100_11111001_11011101_1;
      patterns[58620] = 25'b11100100_11111010_11011110_1;
      patterns[58621] = 25'b11100100_11111011_11011111_1;
      patterns[58622] = 25'b11100100_11111100_11100000_1;
      patterns[58623] = 25'b11100100_11111101_11100001_1;
      patterns[58624] = 25'b11100100_11111110_11100010_1;
      patterns[58625] = 25'b11100100_11111111_11100011_1;
      patterns[58626] = 25'b11100101_00000000_11100101_0;
      patterns[58627] = 25'b11100101_00000001_11100110_0;
      patterns[58628] = 25'b11100101_00000010_11100111_0;
      patterns[58629] = 25'b11100101_00000011_11101000_0;
      patterns[58630] = 25'b11100101_00000100_11101001_0;
      patterns[58631] = 25'b11100101_00000101_11101010_0;
      patterns[58632] = 25'b11100101_00000110_11101011_0;
      patterns[58633] = 25'b11100101_00000111_11101100_0;
      patterns[58634] = 25'b11100101_00001000_11101101_0;
      patterns[58635] = 25'b11100101_00001001_11101110_0;
      patterns[58636] = 25'b11100101_00001010_11101111_0;
      patterns[58637] = 25'b11100101_00001011_11110000_0;
      patterns[58638] = 25'b11100101_00001100_11110001_0;
      patterns[58639] = 25'b11100101_00001101_11110010_0;
      patterns[58640] = 25'b11100101_00001110_11110011_0;
      patterns[58641] = 25'b11100101_00001111_11110100_0;
      patterns[58642] = 25'b11100101_00010000_11110101_0;
      patterns[58643] = 25'b11100101_00010001_11110110_0;
      patterns[58644] = 25'b11100101_00010010_11110111_0;
      patterns[58645] = 25'b11100101_00010011_11111000_0;
      patterns[58646] = 25'b11100101_00010100_11111001_0;
      patterns[58647] = 25'b11100101_00010101_11111010_0;
      patterns[58648] = 25'b11100101_00010110_11111011_0;
      patterns[58649] = 25'b11100101_00010111_11111100_0;
      patterns[58650] = 25'b11100101_00011000_11111101_0;
      patterns[58651] = 25'b11100101_00011001_11111110_0;
      patterns[58652] = 25'b11100101_00011010_11111111_0;
      patterns[58653] = 25'b11100101_00011011_00000000_1;
      patterns[58654] = 25'b11100101_00011100_00000001_1;
      patterns[58655] = 25'b11100101_00011101_00000010_1;
      patterns[58656] = 25'b11100101_00011110_00000011_1;
      patterns[58657] = 25'b11100101_00011111_00000100_1;
      patterns[58658] = 25'b11100101_00100000_00000101_1;
      patterns[58659] = 25'b11100101_00100001_00000110_1;
      patterns[58660] = 25'b11100101_00100010_00000111_1;
      patterns[58661] = 25'b11100101_00100011_00001000_1;
      patterns[58662] = 25'b11100101_00100100_00001001_1;
      patterns[58663] = 25'b11100101_00100101_00001010_1;
      patterns[58664] = 25'b11100101_00100110_00001011_1;
      patterns[58665] = 25'b11100101_00100111_00001100_1;
      patterns[58666] = 25'b11100101_00101000_00001101_1;
      patterns[58667] = 25'b11100101_00101001_00001110_1;
      patterns[58668] = 25'b11100101_00101010_00001111_1;
      patterns[58669] = 25'b11100101_00101011_00010000_1;
      patterns[58670] = 25'b11100101_00101100_00010001_1;
      patterns[58671] = 25'b11100101_00101101_00010010_1;
      patterns[58672] = 25'b11100101_00101110_00010011_1;
      patterns[58673] = 25'b11100101_00101111_00010100_1;
      patterns[58674] = 25'b11100101_00110000_00010101_1;
      patterns[58675] = 25'b11100101_00110001_00010110_1;
      patterns[58676] = 25'b11100101_00110010_00010111_1;
      patterns[58677] = 25'b11100101_00110011_00011000_1;
      patterns[58678] = 25'b11100101_00110100_00011001_1;
      patterns[58679] = 25'b11100101_00110101_00011010_1;
      patterns[58680] = 25'b11100101_00110110_00011011_1;
      patterns[58681] = 25'b11100101_00110111_00011100_1;
      patterns[58682] = 25'b11100101_00111000_00011101_1;
      patterns[58683] = 25'b11100101_00111001_00011110_1;
      patterns[58684] = 25'b11100101_00111010_00011111_1;
      patterns[58685] = 25'b11100101_00111011_00100000_1;
      patterns[58686] = 25'b11100101_00111100_00100001_1;
      patterns[58687] = 25'b11100101_00111101_00100010_1;
      patterns[58688] = 25'b11100101_00111110_00100011_1;
      patterns[58689] = 25'b11100101_00111111_00100100_1;
      patterns[58690] = 25'b11100101_01000000_00100101_1;
      patterns[58691] = 25'b11100101_01000001_00100110_1;
      patterns[58692] = 25'b11100101_01000010_00100111_1;
      patterns[58693] = 25'b11100101_01000011_00101000_1;
      patterns[58694] = 25'b11100101_01000100_00101001_1;
      patterns[58695] = 25'b11100101_01000101_00101010_1;
      patterns[58696] = 25'b11100101_01000110_00101011_1;
      patterns[58697] = 25'b11100101_01000111_00101100_1;
      patterns[58698] = 25'b11100101_01001000_00101101_1;
      patterns[58699] = 25'b11100101_01001001_00101110_1;
      patterns[58700] = 25'b11100101_01001010_00101111_1;
      patterns[58701] = 25'b11100101_01001011_00110000_1;
      patterns[58702] = 25'b11100101_01001100_00110001_1;
      patterns[58703] = 25'b11100101_01001101_00110010_1;
      patterns[58704] = 25'b11100101_01001110_00110011_1;
      patterns[58705] = 25'b11100101_01001111_00110100_1;
      patterns[58706] = 25'b11100101_01010000_00110101_1;
      patterns[58707] = 25'b11100101_01010001_00110110_1;
      patterns[58708] = 25'b11100101_01010010_00110111_1;
      patterns[58709] = 25'b11100101_01010011_00111000_1;
      patterns[58710] = 25'b11100101_01010100_00111001_1;
      patterns[58711] = 25'b11100101_01010101_00111010_1;
      patterns[58712] = 25'b11100101_01010110_00111011_1;
      patterns[58713] = 25'b11100101_01010111_00111100_1;
      patterns[58714] = 25'b11100101_01011000_00111101_1;
      patterns[58715] = 25'b11100101_01011001_00111110_1;
      patterns[58716] = 25'b11100101_01011010_00111111_1;
      patterns[58717] = 25'b11100101_01011011_01000000_1;
      patterns[58718] = 25'b11100101_01011100_01000001_1;
      patterns[58719] = 25'b11100101_01011101_01000010_1;
      patterns[58720] = 25'b11100101_01011110_01000011_1;
      patterns[58721] = 25'b11100101_01011111_01000100_1;
      patterns[58722] = 25'b11100101_01100000_01000101_1;
      patterns[58723] = 25'b11100101_01100001_01000110_1;
      patterns[58724] = 25'b11100101_01100010_01000111_1;
      patterns[58725] = 25'b11100101_01100011_01001000_1;
      patterns[58726] = 25'b11100101_01100100_01001001_1;
      patterns[58727] = 25'b11100101_01100101_01001010_1;
      patterns[58728] = 25'b11100101_01100110_01001011_1;
      patterns[58729] = 25'b11100101_01100111_01001100_1;
      patterns[58730] = 25'b11100101_01101000_01001101_1;
      patterns[58731] = 25'b11100101_01101001_01001110_1;
      patterns[58732] = 25'b11100101_01101010_01001111_1;
      patterns[58733] = 25'b11100101_01101011_01010000_1;
      patterns[58734] = 25'b11100101_01101100_01010001_1;
      patterns[58735] = 25'b11100101_01101101_01010010_1;
      patterns[58736] = 25'b11100101_01101110_01010011_1;
      patterns[58737] = 25'b11100101_01101111_01010100_1;
      patterns[58738] = 25'b11100101_01110000_01010101_1;
      patterns[58739] = 25'b11100101_01110001_01010110_1;
      patterns[58740] = 25'b11100101_01110010_01010111_1;
      patterns[58741] = 25'b11100101_01110011_01011000_1;
      patterns[58742] = 25'b11100101_01110100_01011001_1;
      patterns[58743] = 25'b11100101_01110101_01011010_1;
      patterns[58744] = 25'b11100101_01110110_01011011_1;
      patterns[58745] = 25'b11100101_01110111_01011100_1;
      patterns[58746] = 25'b11100101_01111000_01011101_1;
      patterns[58747] = 25'b11100101_01111001_01011110_1;
      patterns[58748] = 25'b11100101_01111010_01011111_1;
      patterns[58749] = 25'b11100101_01111011_01100000_1;
      patterns[58750] = 25'b11100101_01111100_01100001_1;
      patterns[58751] = 25'b11100101_01111101_01100010_1;
      patterns[58752] = 25'b11100101_01111110_01100011_1;
      patterns[58753] = 25'b11100101_01111111_01100100_1;
      patterns[58754] = 25'b11100101_10000000_01100101_1;
      patterns[58755] = 25'b11100101_10000001_01100110_1;
      patterns[58756] = 25'b11100101_10000010_01100111_1;
      patterns[58757] = 25'b11100101_10000011_01101000_1;
      patterns[58758] = 25'b11100101_10000100_01101001_1;
      patterns[58759] = 25'b11100101_10000101_01101010_1;
      patterns[58760] = 25'b11100101_10000110_01101011_1;
      patterns[58761] = 25'b11100101_10000111_01101100_1;
      patterns[58762] = 25'b11100101_10001000_01101101_1;
      patterns[58763] = 25'b11100101_10001001_01101110_1;
      patterns[58764] = 25'b11100101_10001010_01101111_1;
      patterns[58765] = 25'b11100101_10001011_01110000_1;
      patterns[58766] = 25'b11100101_10001100_01110001_1;
      patterns[58767] = 25'b11100101_10001101_01110010_1;
      patterns[58768] = 25'b11100101_10001110_01110011_1;
      patterns[58769] = 25'b11100101_10001111_01110100_1;
      patterns[58770] = 25'b11100101_10010000_01110101_1;
      patterns[58771] = 25'b11100101_10010001_01110110_1;
      patterns[58772] = 25'b11100101_10010010_01110111_1;
      patterns[58773] = 25'b11100101_10010011_01111000_1;
      patterns[58774] = 25'b11100101_10010100_01111001_1;
      patterns[58775] = 25'b11100101_10010101_01111010_1;
      patterns[58776] = 25'b11100101_10010110_01111011_1;
      patterns[58777] = 25'b11100101_10010111_01111100_1;
      patterns[58778] = 25'b11100101_10011000_01111101_1;
      patterns[58779] = 25'b11100101_10011001_01111110_1;
      patterns[58780] = 25'b11100101_10011010_01111111_1;
      patterns[58781] = 25'b11100101_10011011_10000000_1;
      patterns[58782] = 25'b11100101_10011100_10000001_1;
      patterns[58783] = 25'b11100101_10011101_10000010_1;
      patterns[58784] = 25'b11100101_10011110_10000011_1;
      patterns[58785] = 25'b11100101_10011111_10000100_1;
      patterns[58786] = 25'b11100101_10100000_10000101_1;
      patterns[58787] = 25'b11100101_10100001_10000110_1;
      patterns[58788] = 25'b11100101_10100010_10000111_1;
      patterns[58789] = 25'b11100101_10100011_10001000_1;
      patterns[58790] = 25'b11100101_10100100_10001001_1;
      patterns[58791] = 25'b11100101_10100101_10001010_1;
      patterns[58792] = 25'b11100101_10100110_10001011_1;
      patterns[58793] = 25'b11100101_10100111_10001100_1;
      patterns[58794] = 25'b11100101_10101000_10001101_1;
      patterns[58795] = 25'b11100101_10101001_10001110_1;
      patterns[58796] = 25'b11100101_10101010_10001111_1;
      patterns[58797] = 25'b11100101_10101011_10010000_1;
      patterns[58798] = 25'b11100101_10101100_10010001_1;
      patterns[58799] = 25'b11100101_10101101_10010010_1;
      patterns[58800] = 25'b11100101_10101110_10010011_1;
      patterns[58801] = 25'b11100101_10101111_10010100_1;
      patterns[58802] = 25'b11100101_10110000_10010101_1;
      patterns[58803] = 25'b11100101_10110001_10010110_1;
      patterns[58804] = 25'b11100101_10110010_10010111_1;
      patterns[58805] = 25'b11100101_10110011_10011000_1;
      patterns[58806] = 25'b11100101_10110100_10011001_1;
      patterns[58807] = 25'b11100101_10110101_10011010_1;
      patterns[58808] = 25'b11100101_10110110_10011011_1;
      patterns[58809] = 25'b11100101_10110111_10011100_1;
      patterns[58810] = 25'b11100101_10111000_10011101_1;
      patterns[58811] = 25'b11100101_10111001_10011110_1;
      patterns[58812] = 25'b11100101_10111010_10011111_1;
      patterns[58813] = 25'b11100101_10111011_10100000_1;
      patterns[58814] = 25'b11100101_10111100_10100001_1;
      patterns[58815] = 25'b11100101_10111101_10100010_1;
      patterns[58816] = 25'b11100101_10111110_10100011_1;
      patterns[58817] = 25'b11100101_10111111_10100100_1;
      patterns[58818] = 25'b11100101_11000000_10100101_1;
      patterns[58819] = 25'b11100101_11000001_10100110_1;
      patterns[58820] = 25'b11100101_11000010_10100111_1;
      patterns[58821] = 25'b11100101_11000011_10101000_1;
      patterns[58822] = 25'b11100101_11000100_10101001_1;
      patterns[58823] = 25'b11100101_11000101_10101010_1;
      patterns[58824] = 25'b11100101_11000110_10101011_1;
      patterns[58825] = 25'b11100101_11000111_10101100_1;
      patterns[58826] = 25'b11100101_11001000_10101101_1;
      patterns[58827] = 25'b11100101_11001001_10101110_1;
      patterns[58828] = 25'b11100101_11001010_10101111_1;
      patterns[58829] = 25'b11100101_11001011_10110000_1;
      patterns[58830] = 25'b11100101_11001100_10110001_1;
      patterns[58831] = 25'b11100101_11001101_10110010_1;
      patterns[58832] = 25'b11100101_11001110_10110011_1;
      patterns[58833] = 25'b11100101_11001111_10110100_1;
      patterns[58834] = 25'b11100101_11010000_10110101_1;
      patterns[58835] = 25'b11100101_11010001_10110110_1;
      patterns[58836] = 25'b11100101_11010010_10110111_1;
      patterns[58837] = 25'b11100101_11010011_10111000_1;
      patterns[58838] = 25'b11100101_11010100_10111001_1;
      patterns[58839] = 25'b11100101_11010101_10111010_1;
      patterns[58840] = 25'b11100101_11010110_10111011_1;
      patterns[58841] = 25'b11100101_11010111_10111100_1;
      patterns[58842] = 25'b11100101_11011000_10111101_1;
      patterns[58843] = 25'b11100101_11011001_10111110_1;
      patterns[58844] = 25'b11100101_11011010_10111111_1;
      patterns[58845] = 25'b11100101_11011011_11000000_1;
      patterns[58846] = 25'b11100101_11011100_11000001_1;
      patterns[58847] = 25'b11100101_11011101_11000010_1;
      patterns[58848] = 25'b11100101_11011110_11000011_1;
      patterns[58849] = 25'b11100101_11011111_11000100_1;
      patterns[58850] = 25'b11100101_11100000_11000101_1;
      patterns[58851] = 25'b11100101_11100001_11000110_1;
      patterns[58852] = 25'b11100101_11100010_11000111_1;
      patterns[58853] = 25'b11100101_11100011_11001000_1;
      patterns[58854] = 25'b11100101_11100100_11001001_1;
      patterns[58855] = 25'b11100101_11100101_11001010_1;
      patterns[58856] = 25'b11100101_11100110_11001011_1;
      patterns[58857] = 25'b11100101_11100111_11001100_1;
      patterns[58858] = 25'b11100101_11101000_11001101_1;
      patterns[58859] = 25'b11100101_11101001_11001110_1;
      patterns[58860] = 25'b11100101_11101010_11001111_1;
      patterns[58861] = 25'b11100101_11101011_11010000_1;
      patterns[58862] = 25'b11100101_11101100_11010001_1;
      patterns[58863] = 25'b11100101_11101101_11010010_1;
      patterns[58864] = 25'b11100101_11101110_11010011_1;
      patterns[58865] = 25'b11100101_11101111_11010100_1;
      patterns[58866] = 25'b11100101_11110000_11010101_1;
      patterns[58867] = 25'b11100101_11110001_11010110_1;
      patterns[58868] = 25'b11100101_11110010_11010111_1;
      patterns[58869] = 25'b11100101_11110011_11011000_1;
      patterns[58870] = 25'b11100101_11110100_11011001_1;
      patterns[58871] = 25'b11100101_11110101_11011010_1;
      patterns[58872] = 25'b11100101_11110110_11011011_1;
      patterns[58873] = 25'b11100101_11110111_11011100_1;
      patterns[58874] = 25'b11100101_11111000_11011101_1;
      patterns[58875] = 25'b11100101_11111001_11011110_1;
      patterns[58876] = 25'b11100101_11111010_11011111_1;
      patterns[58877] = 25'b11100101_11111011_11100000_1;
      patterns[58878] = 25'b11100101_11111100_11100001_1;
      patterns[58879] = 25'b11100101_11111101_11100010_1;
      patterns[58880] = 25'b11100101_11111110_11100011_1;
      patterns[58881] = 25'b11100101_11111111_11100100_1;
      patterns[58882] = 25'b11100110_00000000_11100110_0;
      patterns[58883] = 25'b11100110_00000001_11100111_0;
      patterns[58884] = 25'b11100110_00000010_11101000_0;
      patterns[58885] = 25'b11100110_00000011_11101001_0;
      patterns[58886] = 25'b11100110_00000100_11101010_0;
      patterns[58887] = 25'b11100110_00000101_11101011_0;
      patterns[58888] = 25'b11100110_00000110_11101100_0;
      patterns[58889] = 25'b11100110_00000111_11101101_0;
      patterns[58890] = 25'b11100110_00001000_11101110_0;
      patterns[58891] = 25'b11100110_00001001_11101111_0;
      patterns[58892] = 25'b11100110_00001010_11110000_0;
      patterns[58893] = 25'b11100110_00001011_11110001_0;
      patterns[58894] = 25'b11100110_00001100_11110010_0;
      patterns[58895] = 25'b11100110_00001101_11110011_0;
      patterns[58896] = 25'b11100110_00001110_11110100_0;
      patterns[58897] = 25'b11100110_00001111_11110101_0;
      patterns[58898] = 25'b11100110_00010000_11110110_0;
      patterns[58899] = 25'b11100110_00010001_11110111_0;
      patterns[58900] = 25'b11100110_00010010_11111000_0;
      patterns[58901] = 25'b11100110_00010011_11111001_0;
      patterns[58902] = 25'b11100110_00010100_11111010_0;
      patterns[58903] = 25'b11100110_00010101_11111011_0;
      patterns[58904] = 25'b11100110_00010110_11111100_0;
      patterns[58905] = 25'b11100110_00010111_11111101_0;
      patterns[58906] = 25'b11100110_00011000_11111110_0;
      patterns[58907] = 25'b11100110_00011001_11111111_0;
      patterns[58908] = 25'b11100110_00011010_00000000_1;
      patterns[58909] = 25'b11100110_00011011_00000001_1;
      patterns[58910] = 25'b11100110_00011100_00000010_1;
      patterns[58911] = 25'b11100110_00011101_00000011_1;
      patterns[58912] = 25'b11100110_00011110_00000100_1;
      patterns[58913] = 25'b11100110_00011111_00000101_1;
      patterns[58914] = 25'b11100110_00100000_00000110_1;
      patterns[58915] = 25'b11100110_00100001_00000111_1;
      patterns[58916] = 25'b11100110_00100010_00001000_1;
      patterns[58917] = 25'b11100110_00100011_00001001_1;
      patterns[58918] = 25'b11100110_00100100_00001010_1;
      patterns[58919] = 25'b11100110_00100101_00001011_1;
      patterns[58920] = 25'b11100110_00100110_00001100_1;
      patterns[58921] = 25'b11100110_00100111_00001101_1;
      patterns[58922] = 25'b11100110_00101000_00001110_1;
      patterns[58923] = 25'b11100110_00101001_00001111_1;
      patterns[58924] = 25'b11100110_00101010_00010000_1;
      patterns[58925] = 25'b11100110_00101011_00010001_1;
      patterns[58926] = 25'b11100110_00101100_00010010_1;
      patterns[58927] = 25'b11100110_00101101_00010011_1;
      patterns[58928] = 25'b11100110_00101110_00010100_1;
      patterns[58929] = 25'b11100110_00101111_00010101_1;
      patterns[58930] = 25'b11100110_00110000_00010110_1;
      patterns[58931] = 25'b11100110_00110001_00010111_1;
      patterns[58932] = 25'b11100110_00110010_00011000_1;
      patterns[58933] = 25'b11100110_00110011_00011001_1;
      patterns[58934] = 25'b11100110_00110100_00011010_1;
      patterns[58935] = 25'b11100110_00110101_00011011_1;
      patterns[58936] = 25'b11100110_00110110_00011100_1;
      patterns[58937] = 25'b11100110_00110111_00011101_1;
      patterns[58938] = 25'b11100110_00111000_00011110_1;
      patterns[58939] = 25'b11100110_00111001_00011111_1;
      patterns[58940] = 25'b11100110_00111010_00100000_1;
      patterns[58941] = 25'b11100110_00111011_00100001_1;
      patterns[58942] = 25'b11100110_00111100_00100010_1;
      patterns[58943] = 25'b11100110_00111101_00100011_1;
      patterns[58944] = 25'b11100110_00111110_00100100_1;
      patterns[58945] = 25'b11100110_00111111_00100101_1;
      patterns[58946] = 25'b11100110_01000000_00100110_1;
      patterns[58947] = 25'b11100110_01000001_00100111_1;
      patterns[58948] = 25'b11100110_01000010_00101000_1;
      patterns[58949] = 25'b11100110_01000011_00101001_1;
      patterns[58950] = 25'b11100110_01000100_00101010_1;
      patterns[58951] = 25'b11100110_01000101_00101011_1;
      patterns[58952] = 25'b11100110_01000110_00101100_1;
      patterns[58953] = 25'b11100110_01000111_00101101_1;
      patterns[58954] = 25'b11100110_01001000_00101110_1;
      patterns[58955] = 25'b11100110_01001001_00101111_1;
      patterns[58956] = 25'b11100110_01001010_00110000_1;
      patterns[58957] = 25'b11100110_01001011_00110001_1;
      patterns[58958] = 25'b11100110_01001100_00110010_1;
      patterns[58959] = 25'b11100110_01001101_00110011_1;
      patterns[58960] = 25'b11100110_01001110_00110100_1;
      patterns[58961] = 25'b11100110_01001111_00110101_1;
      patterns[58962] = 25'b11100110_01010000_00110110_1;
      patterns[58963] = 25'b11100110_01010001_00110111_1;
      patterns[58964] = 25'b11100110_01010010_00111000_1;
      patterns[58965] = 25'b11100110_01010011_00111001_1;
      patterns[58966] = 25'b11100110_01010100_00111010_1;
      patterns[58967] = 25'b11100110_01010101_00111011_1;
      patterns[58968] = 25'b11100110_01010110_00111100_1;
      patterns[58969] = 25'b11100110_01010111_00111101_1;
      patterns[58970] = 25'b11100110_01011000_00111110_1;
      patterns[58971] = 25'b11100110_01011001_00111111_1;
      patterns[58972] = 25'b11100110_01011010_01000000_1;
      patterns[58973] = 25'b11100110_01011011_01000001_1;
      patterns[58974] = 25'b11100110_01011100_01000010_1;
      patterns[58975] = 25'b11100110_01011101_01000011_1;
      patterns[58976] = 25'b11100110_01011110_01000100_1;
      patterns[58977] = 25'b11100110_01011111_01000101_1;
      patterns[58978] = 25'b11100110_01100000_01000110_1;
      patterns[58979] = 25'b11100110_01100001_01000111_1;
      patterns[58980] = 25'b11100110_01100010_01001000_1;
      patterns[58981] = 25'b11100110_01100011_01001001_1;
      patterns[58982] = 25'b11100110_01100100_01001010_1;
      patterns[58983] = 25'b11100110_01100101_01001011_1;
      patterns[58984] = 25'b11100110_01100110_01001100_1;
      patterns[58985] = 25'b11100110_01100111_01001101_1;
      patterns[58986] = 25'b11100110_01101000_01001110_1;
      patterns[58987] = 25'b11100110_01101001_01001111_1;
      patterns[58988] = 25'b11100110_01101010_01010000_1;
      patterns[58989] = 25'b11100110_01101011_01010001_1;
      patterns[58990] = 25'b11100110_01101100_01010010_1;
      patterns[58991] = 25'b11100110_01101101_01010011_1;
      patterns[58992] = 25'b11100110_01101110_01010100_1;
      patterns[58993] = 25'b11100110_01101111_01010101_1;
      patterns[58994] = 25'b11100110_01110000_01010110_1;
      patterns[58995] = 25'b11100110_01110001_01010111_1;
      patterns[58996] = 25'b11100110_01110010_01011000_1;
      patterns[58997] = 25'b11100110_01110011_01011001_1;
      patterns[58998] = 25'b11100110_01110100_01011010_1;
      patterns[58999] = 25'b11100110_01110101_01011011_1;
      patterns[59000] = 25'b11100110_01110110_01011100_1;
      patterns[59001] = 25'b11100110_01110111_01011101_1;
      patterns[59002] = 25'b11100110_01111000_01011110_1;
      patterns[59003] = 25'b11100110_01111001_01011111_1;
      patterns[59004] = 25'b11100110_01111010_01100000_1;
      patterns[59005] = 25'b11100110_01111011_01100001_1;
      patterns[59006] = 25'b11100110_01111100_01100010_1;
      patterns[59007] = 25'b11100110_01111101_01100011_1;
      patterns[59008] = 25'b11100110_01111110_01100100_1;
      patterns[59009] = 25'b11100110_01111111_01100101_1;
      patterns[59010] = 25'b11100110_10000000_01100110_1;
      patterns[59011] = 25'b11100110_10000001_01100111_1;
      patterns[59012] = 25'b11100110_10000010_01101000_1;
      patterns[59013] = 25'b11100110_10000011_01101001_1;
      patterns[59014] = 25'b11100110_10000100_01101010_1;
      patterns[59015] = 25'b11100110_10000101_01101011_1;
      patterns[59016] = 25'b11100110_10000110_01101100_1;
      patterns[59017] = 25'b11100110_10000111_01101101_1;
      patterns[59018] = 25'b11100110_10001000_01101110_1;
      patterns[59019] = 25'b11100110_10001001_01101111_1;
      patterns[59020] = 25'b11100110_10001010_01110000_1;
      patterns[59021] = 25'b11100110_10001011_01110001_1;
      patterns[59022] = 25'b11100110_10001100_01110010_1;
      patterns[59023] = 25'b11100110_10001101_01110011_1;
      patterns[59024] = 25'b11100110_10001110_01110100_1;
      patterns[59025] = 25'b11100110_10001111_01110101_1;
      patterns[59026] = 25'b11100110_10010000_01110110_1;
      patterns[59027] = 25'b11100110_10010001_01110111_1;
      patterns[59028] = 25'b11100110_10010010_01111000_1;
      patterns[59029] = 25'b11100110_10010011_01111001_1;
      patterns[59030] = 25'b11100110_10010100_01111010_1;
      patterns[59031] = 25'b11100110_10010101_01111011_1;
      patterns[59032] = 25'b11100110_10010110_01111100_1;
      patterns[59033] = 25'b11100110_10010111_01111101_1;
      patterns[59034] = 25'b11100110_10011000_01111110_1;
      patterns[59035] = 25'b11100110_10011001_01111111_1;
      patterns[59036] = 25'b11100110_10011010_10000000_1;
      patterns[59037] = 25'b11100110_10011011_10000001_1;
      patterns[59038] = 25'b11100110_10011100_10000010_1;
      patterns[59039] = 25'b11100110_10011101_10000011_1;
      patterns[59040] = 25'b11100110_10011110_10000100_1;
      patterns[59041] = 25'b11100110_10011111_10000101_1;
      patterns[59042] = 25'b11100110_10100000_10000110_1;
      patterns[59043] = 25'b11100110_10100001_10000111_1;
      patterns[59044] = 25'b11100110_10100010_10001000_1;
      patterns[59045] = 25'b11100110_10100011_10001001_1;
      patterns[59046] = 25'b11100110_10100100_10001010_1;
      patterns[59047] = 25'b11100110_10100101_10001011_1;
      patterns[59048] = 25'b11100110_10100110_10001100_1;
      patterns[59049] = 25'b11100110_10100111_10001101_1;
      patterns[59050] = 25'b11100110_10101000_10001110_1;
      patterns[59051] = 25'b11100110_10101001_10001111_1;
      patterns[59052] = 25'b11100110_10101010_10010000_1;
      patterns[59053] = 25'b11100110_10101011_10010001_1;
      patterns[59054] = 25'b11100110_10101100_10010010_1;
      patterns[59055] = 25'b11100110_10101101_10010011_1;
      patterns[59056] = 25'b11100110_10101110_10010100_1;
      patterns[59057] = 25'b11100110_10101111_10010101_1;
      patterns[59058] = 25'b11100110_10110000_10010110_1;
      patterns[59059] = 25'b11100110_10110001_10010111_1;
      patterns[59060] = 25'b11100110_10110010_10011000_1;
      patterns[59061] = 25'b11100110_10110011_10011001_1;
      patterns[59062] = 25'b11100110_10110100_10011010_1;
      patterns[59063] = 25'b11100110_10110101_10011011_1;
      patterns[59064] = 25'b11100110_10110110_10011100_1;
      patterns[59065] = 25'b11100110_10110111_10011101_1;
      patterns[59066] = 25'b11100110_10111000_10011110_1;
      patterns[59067] = 25'b11100110_10111001_10011111_1;
      patterns[59068] = 25'b11100110_10111010_10100000_1;
      patterns[59069] = 25'b11100110_10111011_10100001_1;
      patterns[59070] = 25'b11100110_10111100_10100010_1;
      patterns[59071] = 25'b11100110_10111101_10100011_1;
      patterns[59072] = 25'b11100110_10111110_10100100_1;
      patterns[59073] = 25'b11100110_10111111_10100101_1;
      patterns[59074] = 25'b11100110_11000000_10100110_1;
      patterns[59075] = 25'b11100110_11000001_10100111_1;
      patterns[59076] = 25'b11100110_11000010_10101000_1;
      patterns[59077] = 25'b11100110_11000011_10101001_1;
      patterns[59078] = 25'b11100110_11000100_10101010_1;
      patterns[59079] = 25'b11100110_11000101_10101011_1;
      patterns[59080] = 25'b11100110_11000110_10101100_1;
      patterns[59081] = 25'b11100110_11000111_10101101_1;
      patterns[59082] = 25'b11100110_11001000_10101110_1;
      patterns[59083] = 25'b11100110_11001001_10101111_1;
      patterns[59084] = 25'b11100110_11001010_10110000_1;
      patterns[59085] = 25'b11100110_11001011_10110001_1;
      patterns[59086] = 25'b11100110_11001100_10110010_1;
      patterns[59087] = 25'b11100110_11001101_10110011_1;
      patterns[59088] = 25'b11100110_11001110_10110100_1;
      patterns[59089] = 25'b11100110_11001111_10110101_1;
      patterns[59090] = 25'b11100110_11010000_10110110_1;
      patterns[59091] = 25'b11100110_11010001_10110111_1;
      patterns[59092] = 25'b11100110_11010010_10111000_1;
      patterns[59093] = 25'b11100110_11010011_10111001_1;
      patterns[59094] = 25'b11100110_11010100_10111010_1;
      patterns[59095] = 25'b11100110_11010101_10111011_1;
      patterns[59096] = 25'b11100110_11010110_10111100_1;
      patterns[59097] = 25'b11100110_11010111_10111101_1;
      patterns[59098] = 25'b11100110_11011000_10111110_1;
      patterns[59099] = 25'b11100110_11011001_10111111_1;
      patterns[59100] = 25'b11100110_11011010_11000000_1;
      patterns[59101] = 25'b11100110_11011011_11000001_1;
      patterns[59102] = 25'b11100110_11011100_11000010_1;
      patterns[59103] = 25'b11100110_11011101_11000011_1;
      patterns[59104] = 25'b11100110_11011110_11000100_1;
      patterns[59105] = 25'b11100110_11011111_11000101_1;
      patterns[59106] = 25'b11100110_11100000_11000110_1;
      patterns[59107] = 25'b11100110_11100001_11000111_1;
      patterns[59108] = 25'b11100110_11100010_11001000_1;
      patterns[59109] = 25'b11100110_11100011_11001001_1;
      patterns[59110] = 25'b11100110_11100100_11001010_1;
      patterns[59111] = 25'b11100110_11100101_11001011_1;
      patterns[59112] = 25'b11100110_11100110_11001100_1;
      patterns[59113] = 25'b11100110_11100111_11001101_1;
      patterns[59114] = 25'b11100110_11101000_11001110_1;
      patterns[59115] = 25'b11100110_11101001_11001111_1;
      patterns[59116] = 25'b11100110_11101010_11010000_1;
      patterns[59117] = 25'b11100110_11101011_11010001_1;
      patterns[59118] = 25'b11100110_11101100_11010010_1;
      patterns[59119] = 25'b11100110_11101101_11010011_1;
      patterns[59120] = 25'b11100110_11101110_11010100_1;
      patterns[59121] = 25'b11100110_11101111_11010101_1;
      patterns[59122] = 25'b11100110_11110000_11010110_1;
      patterns[59123] = 25'b11100110_11110001_11010111_1;
      patterns[59124] = 25'b11100110_11110010_11011000_1;
      patterns[59125] = 25'b11100110_11110011_11011001_1;
      patterns[59126] = 25'b11100110_11110100_11011010_1;
      patterns[59127] = 25'b11100110_11110101_11011011_1;
      patterns[59128] = 25'b11100110_11110110_11011100_1;
      patterns[59129] = 25'b11100110_11110111_11011101_1;
      patterns[59130] = 25'b11100110_11111000_11011110_1;
      patterns[59131] = 25'b11100110_11111001_11011111_1;
      patterns[59132] = 25'b11100110_11111010_11100000_1;
      patterns[59133] = 25'b11100110_11111011_11100001_1;
      patterns[59134] = 25'b11100110_11111100_11100010_1;
      patterns[59135] = 25'b11100110_11111101_11100011_1;
      patterns[59136] = 25'b11100110_11111110_11100100_1;
      patterns[59137] = 25'b11100110_11111111_11100101_1;
      patterns[59138] = 25'b11100111_00000000_11100111_0;
      patterns[59139] = 25'b11100111_00000001_11101000_0;
      patterns[59140] = 25'b11100111_00000010_11101001_0;
      patterns[59141] = 25'b11100111_00000011_11101010_0;
      patterns[59142] = 25'b11100111_00000100_11101011_0;
      patterns[59143] = 25'b11100111_00000101_11101100_0;
      patterns[59144] = 25'b11100111_00000110_11101101_0;
      patterns[59145] = 25'b11100111_00000111_11101110_0;
      patterns[59146] = 25'b11100111_00001000_11101111_0;
      patterns[59147] = 25'b11100111_00001001_11110000_0;
      patterns[59148] = 25'b11100111_00001010_11110001_0;
      patterns[59149] = 25'b11100111_00001011_11110010_0;
      patterns[59150] = 25'b11100111_00001100_11110011_0;
      patterns[59151] = 25'b11100111_00001101_11110100_0;
      patterns[59152] = 25'b11100111_00001110_11110101_0;
      patterns[59153] = 25'b11100111_00001111_11110110_0;
      patterns[59154] = 25'b11100111_00010000_11110111_0;
      patterns[59155] = 25'b11100111_00010001_11111000_0;
      patterns[59156] = 25'b11100111_00010010_11111001_0;
      patterns[59157] = 25'b11100111_00010011_11111010_0;
      patterns[59158] = 25'b11100111_00010100_11111011_0;
      patterns[59159] = 25'b11100111_00010101_11111100_0;
      patterns[59160] = 25'b11100111_00010110_11111101_0;
      patterns[59161] = 25'b11100111_00010111_11111110_0;
      patterns[59162] = 25'b11100111_00011000_11111111_0;
      patterns[59163] = 25'b11100111_00011001_00000000_1;
      patterns[59164] = 25'b11100111_00011010_00000001_1;
      patterns[59165] = 25'b11100111_00011011_00000010_1;
      patterns[59166] = 25'b11100111_00011100_00000011_1;
      patterns[59167] = 25'b11100111_00011101_00000100_1;
      patterns[59168] = 25'b11100111_00011110_00000101_1;
      patterns[59169] = 25'b11100111_00011111_00000110_1;
      patterns[59170] = 25'b11100111_00100000_00000111_1;
      patterns[59171] = 25'b11100111_00100001_00001000_1;
      patterns[59172] = 25'b11100111_00100010_00001001_1;
      patterns[59173] = 25'b11100111_00100011_00001010_1;
      patterns[59174] = 25'b11100111_00100100_00001011_1;
      patterns[59175] = 25'b11100111_00100101_00001100_1;
      patterns[59176] = 25'b11100111_00100110_00001101_1;
      patterns[59177] = 25'b11100111_00100111_00001110_1;
      patterns[59178] = 25'b11100111_00101000_00001111_1;
      patterns[59179] = 25'b11100111_00101001_00010000_1;
      patterns[59180] = 25'b11100111_00101010_00010001_1;
      patterns[59181] = 25'b11100111_00101011_00010010_1;
      patterns[59182] = 25'b11100111_00101100_00010011_1;
      patterns[59183] = 25'b11100111_00101101_00010100_1;
      patterns[59184] = 25'b11100111_00101110_00010101_1;
      patterns[59185] = 25'b11100111_00101111_00010110_1;
      patterns[59186] = 25'b11100111_00110000_00010111_1;
      patterns[59187] = 25'b11100111_00110001_00011000_1;
      patterns[59188] = 25'b11100111_00110010_00011001_1;
      patterns[59189] = 25'b11100111_00110011_00011010_1;
      patterns[59190] = 25'b11100111_00110100_00011011_1;
      patterns[59191] = 25'b11100111_00110101_00011100_1;
      patterns[59192] = 25'b11100111_00110110_00011101_1;
      patterns[59193] = 25'b11100111_00110111_00011110_1;
      patterns[59194] = 25'b11100111_00111000_00011111_1;
      patterns[59195] = 25'b11100111_00111001_00100000_1;
      patterns[59196] = 25'b11100111_00111010_00100001_1;
      patterns[59197] = 25'b11100111_00111011_00100010_1;
      patterns[59198] = 25'b11100111_00111100_00100011_1;
      patterns[59199] = 25'b11100111_00111101_00100100_1;
      patterns[59200] = 25'b11100111_00111110_00100101_1;
      patterns[59201] = 25'b11100111_00111111_00100110_1;
      patterns[59202] = 25'b11100111_01000000_00100111_1;
      patterns[59203] = 25'b11100111_01000001_00101000_1;
      patterns[59204] = 25'b11100111_01000010_00101001_1;
      patterns[59205] = 25'b11100111_01000011_00101010_1;
      patterns[59206] = 25'b11100111_01000100_00101011_1;
      patterns[59207] = 25'b11100111_01000101_00101100_1;
      patterns[59208] = 25'b11100111_01000110_00101101_1;
      patterns[59209] = 25'b11100111_01000111_00101110_1;
      patterns[59210] = 25'b11100111_01001000_00101111_1;
      patterns[59211] = 25'b11100111_01001001_00110000_1;
      patterns[59212] = 25'b11100111_01001010_00110001_1;
      patterns[59213] = 25'b11100111_01001011_00110010_1;
      patterns[59214] = 25'b11100111_01001100_00110011_1;
      patterns[59215] = 25'b11100111_01001101_00110100_1;
      patterns[59216] = 25'b11100111_01001110_00110101_1;
      patterns[59217] = 25'b11100111_01001111_00110110_1;
      patterns[59218] = 25'b11100111_01010000_00110111_1;
      patterns[59219] = 25'b11100111_01010001_00111000_1;
      patterns[59220] = 25'b11100111_01010010_00111001_1;
      patterns[59221] = 25'b11100111_01010011_00111010_1;
      patterns[59222] = 25'b11100111_01010100_00111011_1;
      patterns[59223] = 25'b11100111_01010101_00111100_1;
      patterns[59224] = 25'b11100111_01010110_00111101_1;
      patterns[59225] = 25'b11100111_01010111_00111110_1;
      patterns[59226] = 25'b11100111_01011000_00111111_1;
      patterns[59227] = 25'b11100111_01011001_01000000_1;
      patterns[59228] = 25'b11100111_01011010_01000001_1;
      patterns[59229] = 25'b11100111_01011011_01000010_1;
      patterns[59230] = 25'b11100111_01011100_01000011_1;
      patterns[59231] = 25'b11100111_01011101_01000100_1;
      patterns[59232] = 25'b11100111_01011110_01000101_1;
      patterns[59233] = 25'b11100111_01011111_01000110_1;
      patterns[59234] = 25'b11100111_01100000_01000111_1;
      patterns[59235] = 25'b11100111_01100001_01001000_1;
      patterns[59236] = 25'b11100111_01100010_01001001_1;
      patterns[59237] = 25'b11100111_01100011_01001010_1;
      patterns[59238] = 25'b11100111_01100100_01001011_1;
      patterns[59239] = 25'b11100111_01100101_01001100_1;
      patterns[59240] = 25'b11100111_01100110_01001101_1;
      patterns[59241] = 25'b11100111_01100111_01001110_1;
      patterns[59242] = 25'b11100111_01101000_01001111_1;
      patterns[59243] = 25'b11100111_01101001_01010000_1;
      patterns[59244] = 25'b11100111_01101010_01010001_1;
      patterns[59245] = 25'b11100111_01101011_01010010_1;
      patterns[59246] = 25'b11100111_01101100_01010011_1;
      patterns[59247] = 25'b11100111_01101101_01010100_1;
      patterns[59248] = 25'b11100111_01101110_01010101_1;
      patterns[59249] = 25'b11100111_01101111_01010110_1;
      patterns[59250] = 25'b11100111_01110000_01010111_1;
      patterns[59251] = 25'b11100111_01110001_01011000_1;
      patterns[59252] = 25'b11100111_01110010_01011001_1;
      patterns[59253] = 25'b11100111_01110011_01011010_1;
      patterns[59254] = 25'b11100111_01110100_01011011_1;
      patterns[59255] = 25'b11100111_01110101_01011100_1;
      patterns[59256] = 25'b11100111_01110110_01011101_1;
      patterns[59257] = 25'b11100111_01110111_01011110_1;
      patterns[59258] = 25'b11100111_01111000_01011111_1;
      patterns[59259] = 25'b11100111_01111001_01100000_1;
      patterns[59260] = 25'b11100111_01111010_01100001_1;
      patterns[59261] = 25'b11100111_01111011_01100010_1;
      patterns[59262] = 25'b11100111_01111100_01100011_1;
      patterns[59263] = 25'b11100111_01111101_01100100_1;
      patterns[59264] = 25'b11100111_01111110_01100101_1;
      patterns[59265] = 25'b11100111_01111111_01100110_1;
      patterns[59266] = 25'b11100111_10000000_01100111_1;
      patterns[59267] = 25'b11100111_10000001_01101000_1;
      patterns[59268] = 25'b11100111_10000010_01101001_1;
      patterns[59269] = 25'b11100111_10000011_01101010_1;
      patterns[59270] = 25'b11100111_10000100_01101011_1;
      patterns[59271] = 25'b11100111_10000101_01101100_1;
      patterns[59272] = 25'b11100111_10000110_01101101_1;
      patterns[59273] = 25'b11100111_10000111_01101110_1;
      patterns[59274] = 25'b11100111_10001000_01101111_1;
      patterns[59275] = 25'b11100111_10001001_01110000_1;
      patterns[59276] = 25'b11100111_10001010_01110001_1;
      patterns[59277] = 25'b11100111_10001011_01110010_1;
      patterns[59278] = 25'b11100111_10001100_01110011_1;
      patterns[59279] = 25'b11100111_10001101_01110100_1;
      patterns[59280] = 25'b11100111_10001110_01110101_1;
      patterns[59281] = 25'b11100111_10001111_01110110_1;
      patterns[59282] = 25'b11100111_10010000_01110111_1;
      patterns[59283] = 25'b11100111_10010001_01111000_1;
      patterns[59284] = 25'b11100111_10010010_01111001_1;
      patterns[59285] = 25'b11100111_10010011_01111010_1;
      patterns[59286] = 25'b11100111_10010100_01111011_1;
      patterns[59287] = 25'b11100111_10010101_01111100_1;
      patterns[59288] = 25'b11100111_10010110_01111101_1;
      patterns[59289] = 25'b11100111_10010111_01111110_1;
      patterns[59290] = 25'b11100111_10011000_01111111_1;
      patterns[59291] = 25'b11100111_10011001_10000000_1;
      patterns[59292] = 25'b11100111_10011010_10000001_1;
      patterns[59293] = 25'b11100111_10011011_10000010_1;
      patterns[59294] = 25'b11100111_10011100_10000011_1;
      patterns[59295] = 25'b11100111_10011101_10000100_1;
      patterns[59296] = 25'b11100111_10011110_10000101_1;
      patterns[59297] = 25'b11100111_10011111_10000110_1;
      patterns[59298] = 25'b11100111_10100000_10000111_1;
      patterns[59299] = 25'b11100111_10100001_10001000_1;
      patterns[59300] = 25'b11100111_10100010_10001001_1;
      patterns[59301] = 25'b11100111_10100011_10001010_1;
      patterns[59302] = 25'b11100111_10100100_10001011_1;
      patterns[59303] = 25'b11100111_10100101_10001100_1;
      patterns[59304] = 25'b11100111_10100110_10001101_1;
      patterns[59305] = 25'b11100111_10100111_10001110_1;
      patterns[59306] = 25'b11100111_10101000_10001111_1;
      patterns[59307] = 25'b11100111_10101001_10010000_1;
      patterns[59308] = 25'b11100111_10101010_10010001_1;
      patterns[59309] = 25'b11100111_10101011_10010010_1;
      patterns[59310] = 25'b11100111_10101100_10010011_1;
      patterns[59311] = 25'b11100111_10101101_10010100_1;
      patterns[59312] = 25'b11100111_10101110_10010101_1;
      patterns[59313] = 25'b11100111_10101111_10010110_1;
      patterns[59314] = 25'b11100111_10110000_10010111_1;
      patterns[59315] = 25'b11100111_10110001_10011000_1;
      patterns[59316] = 25'b11100111_10110010_10011001_1;
      patterns[59317] = 25'b11100111_10110011_10011010_1;
      patterns[59318] = 25'b11100111_10110100_10011011_1;
      patterns[59319] = 25'b11100111_10110101_10011100_1;
      patterns[59320] = 25'b11100111_10110110_10011101_1;
      patterns[59321] = 25'b11100111_10110111_10011110_1;
      patterns[59322] = 25'b11100111_10111000_10011111_1;
      patterns[59323] = 25'b11100111_10111001_10100000_1;
      patterns[59324] = 25'b11100111_10111010_10100001_1;
      patterns[59325] = 25'b11100111_10111011_10100010_1;
      patterns[59326] = 25'b11100111_10111100_10100011_1;
      patterns[59327] = 25'b11100111_10111101_10100100_1;
      patterns[59328] = 25'b11100111_10111110_10100101_1;
      patterns[59329] = 25'b11100111_10111111_10100110_1;
      patterns[59330] = 25'b11100111_11000000_10100111_1;
      patterns[59331] = 25'b11100111_11000001_10101000_1;
      patterns[59332] = 25'b11100111_11000010_10101001_1;
      patterns[59333] = 25'b11100111_11000011_10101010_1;
      patterns[59334] = 25'b11100111_11000100_10101011_1;
      patterns[59335] = 25'b11100111_11000101_10101100_1;
      patterns[59336] = 25'b11100111_11000110_10101101_1;
      patterns[59337] = 25'b11100111_11000111_10101110_1;
      patterns[59338] = 25'b11100111_11001000_10101111_1;
      patterns[59339] = 25'b11100111_11001001_10110000_1;
      patterns[59340] = 25'b11100111_11001010_10110001_1;
      patterns[59341] = 25'b11100111_11001011_10110010_1;
      patterns[59342] = 25'b11100111_11001100_10110011_1;
      patterns[59343] = 25'b11100111_11001101_10110100_1;
      patterns[59344] = 25'b11100111_11001110_10110101_1;
      patterns[59345] = 25'b11100111_11001111_10110110_1;
      patterns[59346] = 25'b11100111_11010000_10110111_1;
      patterns[59347] = 25'b11100111_11010001_10111000_1;
      patterns[59348] = 25'b11100111_11010010_10111001_1;
      patterns[59349] = 25'b11100111_11010011_10111010_1;
      patterns[59350] = 25'b11100111_11010100_10111011_1;
      patterns[59351] = 25'b11100111_11010101_10111100_1;
      patterns[59352] = 25'b11100111_11010110_10111101_1;
      patterns[59353] = 25'b11100111_11010111_10111110_1;
      patterns[59354] = 25'b11100111_11011000_10111111_1;
      patterns[59355] = 25'b11100111_11011001_11000000_1;
      patterns[59356] = 25'b11100111_11011010_11000001_1;
      patterns[59357] = 25'b11100111_11011011_11000010_1;
      patterns[59358] = 25'b11100111_11011100_11000011_1;
      patterns[59359] = 25'b11100111_11011101_11000100_1;
      patterns[59360] = 25'b11100111_11011110_11000101_1;
      patterns[59361] = 25'b11100111_11011111_11000110_1;
      patterns[59362] = 25'b11100111_11100000_11000111_1;
      patterns[59363] = 25'b11100111_11100001_11001000_1;
      patterns[59364] = 25'b11100111_11100010_11001001_1;
      patterns[59365] = 25'b11100111_11100011_11001010_1;
      patterns[59366] = 25'b11100111_11100100_11001011_1;
      patterns[59367] = 25'b11100111_11100101_11001100_1;
      patterns[59368] = 25'b11100111_11100110_11001101_1;
      patterns[59369] = 25'b11100111_11100111_11001110_1;
      patterns[59370] = 25'b11100111_11101000_11001111_1;
      patterns[59371] = 25'b11100111_11101001_11010000_1;
      patterns[59372] = 25'b11100111_11101010_11010001_1;
      patterns[59373] = 25'b11100111_11101011_11010010_1;
      patterns[59374] = 25'b11100111_11101100_11010011_1;
      patterns[59375] = 25'b11100111_11101101_11010100_1;
      patterns[59376] = 25'b11100111_11101110_11010101_1;
      patterns[59377] = 25'b11100111_11101111_11010110_1;
      patterns[59378] = 25'b11100111_11110000_11010111_1;
      patterns[59379] = 25'b11100111_11110001_11011000_1;
      patterns[59380] = 25'b11100111_11110010_11011001_1;
      patterns[59381] = 25'b11100111_11110011_11011010_1;
      patterns[59382] = 25'b11100111_11110100_11011011_1;
      patterns[59383] = 25'b11100111_11110101_11011100_1;
      patterns[59384] = 25'b11100111_11110110_11011101_1;
      patterns[59385] = 25'b11100111_11110111_11011110_1;
      patterns[59386] = 25'b11100111_11111000_11011111_1;
      patterns[59387] = 25'b11100111_11111001_11100000_1;
      patterns[59388] = 25'b11100111_11111010_11100001_1;
      patterns[59389] = 25'b11100111_11111011_11100010_1;
      patterns[59390] = 25'b11100111_11111100_11100011_1;
      patterns[59391] = 25'b11100111_11111101_11100100_1;
      patterns[59392] = 25'b11100111_11111110_11100101_1;
      patterns[59393] = 25'b11100111_11111111_11100110_1;
      patterns[59394] = 25'b11101000_00000000_11101000_0;
      patterns[59395] = 25'b11101000_00000001_11101001_0;
      patterns[59396] = 25'b11101000_00000010_11101010_0;
      patterns[59397] = 25'b11101000_00000011_11101011_0;
      patterns[59398] = 25'b11101000_00000100_11101100_0;
      patterns[59399] = 25'b11101000_00000101_11101101_0;
      patterns[59400] = 25'b11101000_00000110_11101110_0;
      patterns[59401] = 25'b11101000_00000111_11101111_0;
      patterns[59402] = 25'b11101000_00001000_11110000_0;
      patterns[59403] = 25'b11101000_00001001_11110001_0;
      patterns[59404] = 25'b11101000_00001010_11110010_0;
      patterns[59405] = 25'b11101000_00001011_11110011_0;
      patterns[59406] = 25'b11101000_00001100_11110100_0;
      patterns[59407] = 25'b11101000_00001101_11110101_0;
      patterns[59408] = 25'b11101000_00001110_11110110_0;
      patterns[59409] = 25'b11101000_00001111_11110111_0;
      patterns[59410] = 25'b11101000_00010000_11111000_0;
      patterns[59411] = 25'b11101000_00010001_11111001_0;
      patterns[59412] = 25'b11101000_00010010_11111010_0;
      patterns[59413] = 25'b11101000_00010011_11111011_0;
      patterns[59414] = 25'b11101000_00010100_11111100_0;
      patterns[59415] = 25'b11101000_00010101_11111101_0;
      patterns[59416] = 25'b11101000_00010110_11111110_0;
      patterns[59417] = 25'b11101000_00010111_11111111_0;
      patterns[59418] = 25'b11101000_00011000_00000000_1;
      patterns[59419] = 25'b11101000_00011001_00000001_1;
      patterns[59420] = 25'b11101000_00011010_00000010_1;
      patterns[59421] = 25'b11101000_00011011_00000011_1;
      patterns[59422] = 25'b11101000_00011100_00000100_1;
      patterns[59423] = 25'b11101000_00011101_00000101_1;
      patterns[59424] = 25'b11101000_00011110_00000110_1;
      patterns[59425] = 25'b11101000_00011111_00000111_1;
      patterns[59426] = 25'b11101000_00100000_00001000_1;
      patterns[59427] = 25'b11101000_00100001_00001001_1;
      patterns[59428] = 25'b11101000_00100010_00001010_1;
      patterns[59429] = 25'b11101000_00100011_00001011_1;
      patterns[59430] = 25'b11101000_00100100_00001100_1;
      patterns[59431] = 25'b11101000_00100101_00001101_1;
      patterns[59432] = 25'b11101000_00100110_00001110_1;
      patterns[59433] = 25'b11101000_00100111_00001111_1;
      patterns[59434] = 25'b11101000_00101000_00010000_1;
      patterns[59435] = 25'b11101000_00101001_00010001_1;
      patterns[59436] = 25'b11101000_00101010_00010010_1;
      patterns[59437] = 25'b11101000_00101011_00010011_1;
      patterns[59438] = 25'b11101000_00101100_00010100_1;
      patterns[59439] = 25'b11101000_00101101_00010101_1;
      patterns[59440] = 25'b11101000_00101110_00010110_1;
      patterns[59441] = 25'b11101000_00101111_00010111_1;
      patterns[59442] = 25'b11101000_00110000_00011000_1;
      patterns[59443] = 25'b11101000_00110001_00011001_1;
      patterns[59444] = 25'b11101000_00110010_00011010_1;
      patterns[59445] = 25'b11101000_00110011_00011011_1;
      patterns[59446] = 25'b11101000_00110100_00011100_1;
      patterns[59447] = 25'b11101000_00110101_00011101_1;
      patterns[59448] = 25'b11101000_00110110_00011110_1;
      patterns[59449] = 25'b11101000_00110111_00011111_1;
      patterns[59450] = 25'b11101000_00111000_00100000_1;
      patterns[59451] = 25'b11101000_00111001_00100001_1;
      patterns[59452] = 25'b11101000_00111010_00100010_1;
      patterns[59453] = 25'b11101000_00111011_00100011_1;
      patterns[59454] = 25'b11101000_00111100_00100100_1;
      patterns[59455] = 25'b11101000_00111101_00100101_1;
      patterns[59456] = 25'b11101000_00111110_00100110_1;
      patterns[59457] = 25'b11101000_00111111_00100111_1;
      patterns[59458] = 25'b11101000_01000000_00101000_1;
      patterns[59459] = 25'b11101000_01000001_00101001_1;
      patterns[59460] = 25'b11101000_01000010_00101010_1;
      patterns[59461] = 25'b11101000_01000011_00101011_1;
      patterns[59462] = 25'b11101000_01000100_00101100_1;
      patterns[59463] = 25'b11101000_01000101_00101101_1;
      patterns[59464] = 25'b11101000_01000110_00101110_1;
      patterns[59465] = 25'b11101000_01000111_00101111_1;
      patterns[59466] = 25'b11101000_01001000_00110000_1;
      patterns[59467] = 25'b11101000_01001001_00110001_1;
      patterns[59468] = 25'b11101000_01001010_00110010_1;
      patterns[59469] = 25'b11101000_01001011_00110011_1;
      patterns[59470] = 25'b11101000_01001100_00110100_1;
      patterns[59471] = 25'b11101000_01001101_00110101_1;
      patterns[59472] = 25'b11101000_01001110_00110110_1;
      patterns[59473] = 25'b11101000_01001111_00110111_1;
      patterns[59474] = 25'b11101000_01010000_00111000_1;
      patterns[59475] = 25'b11101000_01010001_00111001_1;
      patterns[59476] = 25'b11101000_01010010_00111010_1;
      patterns[59477] = 25'b11101000_01010011_00111011_1;
      patterns[59478] = 25'b11101000_01010100_00111100_1;
      patterns[59479] = 25'b11101000_01010101_00111101_1;
      patterns[59480] = 25'b11101000_01010110_00111110_1;
      patterns[59481] = 25'b11101000_01010111_00111111_1;
      patterns[59482] = 25'b11101000_01011000_01000000_1;
      patterns[59483] = 25'b11101000_01011001_01000001_1;
      patterns[59484] = 25'b11101000_01011010_01000010_1;
      patterns[59485] = 25'b11101000_01011011_01000011_1;
      patterns[59486] = 25'b11101000_01011100_01000100_1;
      patterns[59487] = 25'b11101000_01011101_01000101_1;
      patterns[59488] = 25'b11101000_01011110_01000110_1;
      patterns[59489] = 25'b11101000_01011111_01000111_1;
      patterns[59490] = 25'b11101000_01100000_01001000_1;
      patterns[59491] = 25'b11101000_01100001_01001001_1;
      patterns[59492] = 25'b11101000_01100010_01001010_1;
      patterns[59493] = 25'b11101000_01100011_01001011_1;
      patterns[59494] = 25'b11101000_01100100_01001100_1;
      patterns[59495] = 25'b11101000_01100101_01001101_1;
      patterns[59496] = 25'b11101000_01100110_01001110_1;
      patterns[59497] = 25'b11101000_01100111_01001111_1;
      patterns[59498] = 25'b11101000_01101000_01010000_1;
      patterns[59499] = 25'b11101000_01101001_01010001_1;
      patterns[59500] = 25'b11101000_01101010_01010010_1;
      patterns[59501] = 25'b11101000_01101011_01010011_1;
      patterns[59502] = 25'b11101000_01101100_01010100_1;
      patterns[59503] = 25'b11101000_01101101_01010101_1;
      patterns[59504] = 25'b11101000_01101110_01010110_1;
      patterns[59505] = 25'b11101000_01101111_01010111_1;
      patterns[59506] = 25'b11101000_01110000_01011000_1;
      patterns[59507] = 25'b11101000_01110001_01011001_1;
      patterns[59508] = 25'b11101000_01110010_01011010_1;
      patterns[59509] = 25'b11101000_01110011_01011011_1;
      patterns[59510] = 25'b11101000_01110100_01011100_1;
      patterns[59511] = 25'b11101000_01110101_01011101_1;
      patterns[59512] = 25'b11101000_01110110_01011110_1;
      patterns[59513] = 25'b11101000_01110111_01011111_1;
      patterns[59514] = 25'b11101000_01111000_01100000_1;
      patterns[59515] = 25'b11101000_01111001_01100001_1;
      patterns[59516] = 25'b11101000_01111010_01100010_1;
      patterns[59517] = 25'b11101000_01111011_01100011_1;
      patterns[59518] = 25'b11101000_01111100_01100100_1;
      patterns[59519] = 25'b11101000_01111101_01100101_1;
      patterns[59520] = 25'b11101000_01111110_01100110_1;
      patterns[59521] = 25'b11101000_01111111_01100111_1;
      patterns[59522] = 25'b11101000_10000000_01101000_1;
      patterns[59523] = 25'b11101000_10000001_01101001_1;
      patterns[59524] = 25'b11101000_10000010_01101010_1;
      patterns[59525] = 25'b11101000_10000011_01101011_1;
      patterns[59526] = 25'b11101000_10000100_01101100_1;
      patterns[59527] = 25'b11101000_10000101_01101101_1;
      patterns[59528] = 25'b11101000_10000110_01101110_1;
      patterns[59529] = 25'b11101000_10000111_01101111_1;
      patterns[59530] = 25'b11101000_10001000_01110000_1;
      patterns[59531] = 25'b11101000_10001001_01110001_1;
      patterns[59532] = 25'b11101000_10001010_01110010_1;
      patterns[59533] = 25'b11101000_10001011_01110011_1;
      patterns[59534] = 25'b11101000_10001100_01110100_1;
      patterns[59535] = 25'b11101000_10001101_01110101_1;
      patterns[59536] = 25'b11101000_10001110_01110110_1;
      patterns[59537] = 25'b11101000_10001111_01110111_1;
      patterns[59538] = 25'b11101000_10010000_01111000_1;
      patterns[59539] = 25'b11101000_10010001_01111001_1;
      patterns[59540] = 25'b11101000_10010010_01111010_1;
      patterns[59541] = 25'b11101000_10010011_01111011_1;
      patterns[59542] = 25'b11101000_10010100_01111100_1;
      patterns[59543] = 25'b11101000_10010101_01111101_1;
      patterns[59544] = 25'b11101000_10010110_01111110_1;
      patterns[59545] = 25'b11101000_10010111_01111111_1;
      patterns[59546] = 25'b11101000_10011000_10000000_1;
      patterns[59547] = 25'b11101000_10011001_10000001_1;
      patterns[59548] = 25'b11101000_10011010_10000010_1;
      patterns[59549] = 25'b11101000_10011011_10000011_1;
      patterns[59550] = 25'b11101000_10011100_10000100_1;
      patterns[59551] = 25'b11101000_10011101_10000101_1;
      patterns[59552] = 25'b11101000_10011110_10000110_1;
      patterns[59553] = 25'b11101000_10011111_10000111_1;
      patterns[59554] = 25'b11101000_10100000_10001000_1;
      patterns[59555] = 25'b11101000_10100001_10001001_1;
      patterns[59556] = 25'b11101000_10100010_10001010_1;
      patterns[59557] = 25'b11101000_10100011_10001011_1;
      patterns[59558] = 25'b11101000_10100100_10001100_1;
      patterns[59559] = 25'b11101000_10100101_10001101_1;
      patterns[59560] = 25'b11101000_10100110_10001110_1;
      patterns[59561] = 25'b11101000_10100111_10001111_1;
      patterns[59562] = 25'b11101000_10101000_10010000_1;
      patterns[59563] = 25'b11101000_10101001_10010001_1;
      patterns[59564] = 25'b11101000_10101010_10010010_1;
      patterns[59565] = 25'b11101000_10101011_10010011_1;
      patterns[59566] = 25'b11101000_10101100_10010100_1;
      patterns[59567] = 25'b11101000_10101101_10010101_1;
      patterns[59568] = 25'b11101000_10101110_10010110_1;
      patterns[59569] = 25'b11101000_10101111_10010111_1;
      patterns[59570] = 25'b11101000_10110000_10011000_1;
      patterns[59571] = 25'b11101000_10110001_10011001_1;
      patterns[59572] = 25'b11101000_10110010_10011010_1;
      patterns[59573] = 25'b11101000_10110011_10011011_1;
      patterns[59574] = 25'b11101000_10110100_10011100_1;
      patterns[59575] = 25'b11101000_10110101_10011101_1;
      patterns[59576] = 25'b11101000_10110110_10011110_1;
      patterns[59577] = 25'b11101000_10110111_10011111_1;
      patterns[59578] = 25'b11101000_10111000_10100000_1;
      patterns[59579] = 25'b11101000_10111001_10100001_1;
      patterns[59580] = 25'b11101000_10111010_10100010_1;
      patterns[59581] = 25'b11101000_10111011_10100011_1;
      patterns[59582] = 25'b11101000_10111100_10100100_1;
      patterns[59583] = 25'b11101000_10111101_10100101_1;
      patterns[59584] = 25'b11101000_10111110_10100110_1;
      patterns[59585] = 25'b11101000_10111111_10100111_1;
      patterns[59586] = 25'b11101000_11000000_10101000_1;
      patterns[59587] = 25'b11101000_11000001_10101001_1;
      patterns[59588] = 25'b11101000_11000010_10101010_1;
      patterns[59589] = 25'b11101000_11000011_10101011_1;
      patterns[59590] = 25'b11101000_11000100_10101100_1;
      patterns[59591] = 25'b11101000_11000101_10101101_1;
      patterns[59592] = 25'b11101000_11000110_10101110_1;
      patterns[59593] = 25'b11101000_11000111_10101111_1;
      patterns[59594] = 25'b11101000_11001000_10110000_1;
      patterns[59595] = 25'b11101000_11001001_10110001_1;
      patterns[59596] = 25'b11101000_11001010_10110010_1;
      patterns[59597] = 25'b11101000_11001011_10110011_1;
      patterns[59598] = 25'b11101000_11001100_10110100_1;
      patterns[59599] = 25'b11101000_11001101_10110101_1;
      patterns[59600] = 25'b11101000_11001110_10110110_1;
      patterns[59601] = 25'b11101000_11001111_10110111_1;
      patterns[59602] = 25'b11101000_11010000_10111000_1;
      patterns[59603] = 25'b11101000_11010001_10111001_1;
      patterns[59604] = 25'b11101000_11010010_10111010_1;
      patterns[59605] = 25'b11101000_11010011_10111011_1;
      patterns[59606] = 25'b11101000_11010100_10111100_1;
      patterns[59607] = 25'b11101000_11010101_10111101_1;
      patterns[59608] = 25'b11101000_11010110_10111110_1;
      patterns[59609] = 25'b11101000_11010111_10111111_1;
      patterns[59610] = 25'b11101000_11011000_11000000_1;
      patterns[59611] = 25'b11101000_11011001_11000001_1;
      patterns[59612] = 25'b11101000_11011010_11000010_1;
      patterns[59613] = 25'b11101000_11011011_11000011_1;
      patterns[59614] = 25'b11101000_11011100_11000100_1;
      patterns[59615] = 25'b11101000_11011101_11000101_1;
      patterns[59616] = 25'b11101000_11011110_11000110_1;
      patterns[59617] = 25'b11101000_11011111_11000111_1;
      patterns[59618] = 25'b11101000_11100000_11001000_1;
      patterns[59619] = 25'b11101000_11100001_11001001_1;
      patterns[59620] = 25'b11101000_11100010_11001010_1;
      patterns[59621] = 25'b11101000_11100011_11001011_1;
      patterns[59622] = 25'b11101000_11100100_11001100_1;
      patterns[59623] = 25'b11101000_11100101_11001101_1;
      patterns[59624] = 25'b11101000_11100110_11001110_1;
      patterns[59625] = 25'b11101000_11100111_11001111_1;
      patterns[59626] = 25'b11101000_11101000_11010000_1;
      patterns[59627] = 25'b11101000_11101001_11010001_1;
      patterns[59628] = 25'b11101000_11101010_11010010_1;
      patterns[59629] = 25'b11101000_11101011_11010011_1;
      patterns[59630] = 25'b11101000_11101100_11010100_1;
      patterns[59631] = 25'b11101000_11101101_11010101_1;
      patterns[59632] = 25'b11101000_11101110_11010110_1;
      patterns[59633] = 25'b11101000_11101111_11010111_1;
      patterns[59634] = 25'b11101000_11110000_11011000_1;
      patterns[59635] = 25'b11101000_11110001_11011001_1;
      patterns[59636] = 25'b11101000_11110010_11011010_1;
      patterns[59637] = 25'b11101000_11110011_11011011_1;
      patterns[59638] = 25'b11101000_11110100_11011100_1;
      patterns[59639] = 25'b11101000_11110101_11011101_1;
      patterns[59640] = 25'b11101000_11110110_11011110_1;
      patterns[59641] = 25'b11101000_11110111_11011111_1;
      patterns[59642] = 25'b11101000_11111000_11100000_1;
      patterns[59643] = 25'b11101000_11111001_11100001_1;
      patterns[59644] = 25'b11101000_11111010_11100010_1;
      patterns[59645] = 25'b11101000_11111011_11100011_1;
      patterns[59646] = 25'b11101000_11111100_11100100_1;
      patterns[59647] = 25'b11101000_11111101_11100101_1;
      patterns[59648] = 25'b11101000_11111110_11100110_1;
      patterns[59649] = 25'b11101000_11111111_11100111_1;
      patterns[59650] = 25'b11101001_00000000_11101001_0;
      patterns[59651] = 25'b11101001_00000001_11101010_0;
      patterns[59652] = 25'b11101001_00000010_11101011_0;
      patterns[59653] = 25'b11101001_00000011_11101100_0;
      patterns[59654] = 25'b11101001_00000100_11101101_0;
      patterns[59655] = 25'b11101001_00000101_11101110_0;
      patterns[59656] = 25'b11101001_00000110_11101111_0;
      patterns[59657] = 25'b11101001_00000111_11110000_0;
      patterns[59658] = 25'b11101001_00001000_11110001_0;
      patterns[59659] = 25'b11101001_00001001_11110010_0;
      patterns[59660] = 25'b11101001_00001010_11110011_0;
      patterns[59661] = 25'b11101001_00001011_11110100_0;
      patterns[59662] = 25'b11101001_00001100_11110101_0;
      patterns[59663] = 25'b11101001_00001101_11110110_0;
      patterns[59664] = 25'b11101001_00001110_11110111_0;
      patterns[59665] = 25'b11101001_00001111_11111000_0;
      patterns[59666] = 25'b11101001_00010000_11111001_0;
      patterns[59667] = 25'b11101001_00010001_11111010_0;
      patterns[59668] = 25'b11101001_00010010_11111011_0;
      patterns[59669] = 25'b11101001_00010011_11111100_0;
      patterns[59670] = 25'b11101001_00010100_11111101_0;
      patterns[59671] = 25'b11101001_00010101_11111110_0;
      patterns[59672] = 25'b11101001_00010110_11111111_0;
      patterns[59673] = 25'b11101001_00010111_00000000_1;
      patterns[59674] = 25'b11101001_00011000_00000001_1;
      patterns[59675] = 25'b11101001_00011001_00000010_1;
      patterns[59676] = 25'b11101001_00011010_00000011_1;
      patterns[59677] = 25'b11101001_00011011_00000100_1;
      patterns[59678] = 25'b11101001_00011100_00000101_1;
      patterns[59679] = 25'b11101001_00011101_00000110_1;
      patterns[59680] = 25'b11101001_00011110_00000111_1;
      patterns[59681] = 25'b11101001_00011111_00001000_1;
      patterns[59682] = 25'b11101001_00100000_00001001_1;
      patterns[59683] = 25'b11101001_00100001_00001010_1;
      patterns[59684] = 25'b11101001_00100010_00001011_1;
      patterns[59685] = 25'b11101001_00100011_00001100_1;
      patterns[59686] = 25'b11101001_00100100_00001101_1;
      patterns[59687] = 25'b11101001_00100101_00001110_1;
      patterns[59688] = 25'b11101001_00100110_00001111_1;
      patterns[59689] = 25'b11101001_00100111_00010000_1;
      patterns[59690] = 25'b11101001_00101000_00010001_1;
      patterns[59691] = 25'b11101001_00101001_00010010_1;
      patterns[59692] = 25'b11101001_00101010_00010011_1;
      patterns[59693] = 25'b11101001_00101011_00010100_1;
      patterns[59694] = 25'b11101001_00101100_00010101_1;
      patterns[59695] = 25'b11101001_00101101_00010110_1;
      patterns[59696] = 25'b11101001_00101110_00010111_1;
      patterns[59697] = 25'b11101001_00101111_00011000_1;
      patterns[59698] = 25'b11101001_00110000_00011001_1;
      patterns[59699] = 25'b11101001_00110001_00011010_1;
      patterns[59700] = 25'b11101001_00110010_00011011_1;
      patterns[59701] = 25'b11101001_00110011_00011100_1;
      patterns[59702] = 25'b11101001_00110100_00011101_1;
      patterns[59703] = 25'b11101001_00110101_00011110_1;
      patterns[59704] = 25'b11101001_00110110_00011111_1;
      patterns[59705] = 25'b11101001_00110111_00100000_1;
      patterns[59706] = 25'b11101001_00111000_00100001_1;
      patterns[59707] = 25'b11101001_00111001_00100010_1;
      patterns[59708] = 25'b11101001_00111010_00100011_1;
      patterns[59709] = 25'b11101001_00111011_00100100_1;
      patterns[59710] = 25'b11101001_00111100_00100101_1;
      patterns[59711] = 25'b11101001_00111101_00100110_1;
      patterns[59712] = 25'b11101001_00111110_00100111_1;
      patterns[59713] = 25'b11101001_00111111_00101000_1;
      patterns[59714] = 25'b11101001_01000000_00101001_1;
      patterns[59715] = 25'b11101001_01000001_00101010_1;
      patterns[59716] = 25'b11101001_01000010_00101011_1;
      patterns[59717] = 25'b11101001_01000011_00101100_1;
      patterns[59718] = 25'b11101001_01000100_00101101_1;
      patterns[59719] = 25'b11101001_01000101_00101110_1;
      patterns[59720] = 25'b11101001_01000110_00101111_1;
      patterns[59721] = 25'b11101001_01000111_00110000_1;
      patterns[59722] = 25'b11101001_01001000_00110001_1;
      patterns[59723] = 25'b11101001_01001001_00110010_1;
      patterns[59724] = 25'b11101001_01001010_00110011_1;
      patterns[59725] = 25'b11101001_01001011_00110100_1;
      patterns[59726] = 25'b11101001_01001100_00110101_1;
      patterns[59727] = 25'b11101001_01001101_00110110_1;
      patterns[59728] = 25'b11101001_01001110_00110111_1;
      patterns[59729] = 25'b11101001_01001111_00111000_1;
      patterns[59730] = 25'b11101001_01010000_00111001_1;
      patterns[59731] = 25'b11101001_01010001_00111010_1;
      patterns[59732] = 25'b11101001_01010010_00111011_1;
      patterns[59733] = 25'b11101001_01010011_00111100_1;
      patterns[59734] = 25'b11101001_01010100_00111101_1;
      patterns[59735] = 25'b11101001_01010101_00111110_1;
      patterns[59736] = 25'b11101001_01010110_00111111_1;
      patterns[59737] = 25'b11101001_01010111_01000000_1;
      patterns[59738] = 25'b11101001_01011000_01000001_1;
      patterns[59739] = 25'b11101001_01011001_01000010_1;
      patterns[59740] = 25'b11101001_01011010_01000011_1;
      patterns[59741] = 25'b11101001_01011011_01000100_1;
      patterns[59742] = 25'b11101001_01011100_01000101_1;
      patterns[59743] = 25'b11101001_01011101_01000110_1;
      patterns[59744] = 25'b11101001_01011110_01000111_1;
      patterns[59745] = 25'b11101001_01011111_01001000_1;
      patterns[59746] = 25'b11101001_01100000_01001001_1;
      patterns[59747] = 25'b11101001_01100001_01001010_1;
      patterns[59748] = 25'b11101001_01100010_01001011_1;
      patterns[59749] = 25'b11101001_01100011_01001100_1;
      patterns[59750] = 25'b11101001_01100100_01001101_1;
      patterns[59751] = 25'b11101001_01100101_01001110_1;
      patterns[59752] = 25'b11101001_01100110_01001111_1;
      patterns[59753] = 25'b11101001_01100111_01010000_1;
      patterns[59754] = 25'b11101001_01101000_01010001_1;
      patterns[59755] = 25'b11101001_01101001_01010010_1;
      patterns[59756] = 25'b11101001_01101010_01010011_1;
      patterns[59757] = 25'b11101001_01101011_01010100_1;
      patterns[59758] = 25'b11101001_01101100_01010101_1;
      patterns[59759] = 25'b11101001_01101101_01010110_1;
      patterns[59760] = 25'b11101001_01101110_01010111_1;
      patterns[59761] = 25'b11101001_01101111_01011000_1;
      patterns[59762] = 25'b11101001_01110000_01011001_1;
      patterns[59763] = 25'b11101001_01110001_01011010_1;
      patterns[59764] = 25'b11101001_01110010_01011011_1;
      patterns[59765] = 25'b11101001_01110011_01011100_1;
      patterns[59766] = 25'b11101001_01110100_01011101_1;
      patterns[59767] = 25'b11101001_01110101_01011110_1;
      patterns[59768] = 25'b11101001_01110110_01011111_1;
      patterns[59769] = 25'b11101001_01110111_01100000_1;
      patterns[59770] = 25'b11101001_01111000_01100001_1;
      patterns[59771] = 25'b11101001_01111001_01100010_1;
      patterns[59772] = 25'b11101001_01111010_01100011_1;
      patterns[59773] = 25'b11101001_01111011_01100100_1;
      patterns[59774] = 25'b11101001_01111100_01100101_1;
      patterns[59775] = 25'b11101001_01111101_01100110_1;
      patterns[59776] = 25'b11101001_01111110_01100111_1;
      patterns[59777] = 25'b11101001_01111111_01101000_1;
      patterns[59778] = 25'b11101001_10000000_01101001_1;
      patterns[59779] = 25'b11101001_10000001_01101010_1;
      patterns[59780] = 25'b11101001_10000010_01101011_1;
      patterns[59781] = 25'b11101001_10000011_01101100_1;
      patterns[59782] = 25'b11101001_10000100_01101101_1;
      patterns[59783] = 25'b11101001_10000101_01101110_1;
      patterns[59784] = 25'b11101001_10000110_01101111_1;
      patterns[59785] = 25'b11101001_10000111_01110000_1;
      patterns[59786] = 25'b11101001_10001000_01110001_1;
      patterns[59787] = 25'b11101001_10001001_01110010_1;
      patterns[59788] = 25'b11101001_10001010_01110011_1;
      patterns[59789] = 25'b11101001_10001011_01110100_1;
      patterns[59790] = 25'b11101001_10001100_01110101_1;
      patterns[59791] = 25'b11101001_10001101_01110110_1;
      patterns[59792] = 25'b11101001_10001110_01110111_1;
      patterns[59793] = 25'b11101001_10001111_01111000_1;
      patterns[59794] = 25'b11101001_10010000_01111001_1;
      patterns[59795] = 25'b11101001_10010001_01111010_1;
      patterns[59796] = 25'b11101001_10010010_01111011_1;
      patterns[59797] = 25'b11101001_10010011_01111100_1;
      patterns[59798] = 25'b11101001_10010100_01111101_1;
      patterns[59799] = 25'b11101001_10010101_01111110_1;
      patterns[59800] = 25'b11101001_10010110_01111111_1;
      patterns[59801] = 25'b11101001_10010111_10000000_1;
      patterns[59802] = 25'b11101001_10011000_10000001_1;
      patterns[59803] = 25'b11101001_10011001_10000010_1;
      patterns[59804] = 25'b11101001_10011010_10000011_1;
      patterns[59805] = 25'b11101001_10011011_10000100_1;
      patterns[59806] = 25'b11101001_10011100_10000101_1;
      patterns[59807] = 25'b11101001_10011101_10000110_1;
      patterns[59808] = 25'b11101001_10011110_10000111_1;
      patterns[59809] = 25'b11101001_10011111_10001000_1;
      patterns[59810] = 25'b11101001_10100000_10001001_1;
      patterns[59811] = 25'b11101001_10100001_10001010_1;
      patterns[59812] = 25'b11101001_10100010_10001011_1;
      patterns[59813] = 25'b11101001_10100011_10001100_1;
      patterns[59814] = 25'b11101001_10100100_10001101_1;
      patterns[59815] = 25'b11101001_10100101_10001110_1;
      patterns[59816] = 25'b11101001_10100110_10001111_1;
      patterns[59817] = 25'b11101001_10100111_10010000_1;
      patterns[59818] = 25'b11101001_10101000_10010001_1;
      patterns[59819] = 25'b11101001_10101001_10010010_1;
      patterns[59820] = 25'b11101001_10101010_10010011_1;
      patterns[59821] = 25'b11101001_10101011_10010100_1;
      patterns[59822] = 25'b11101001_10101100_10010101_1;
      patterns[59823] = 25'b11101001_10101101_10010110_1;
      patterns[59824] = 25'b11101001_10101110_10010111_1;
      patterns[59825] = 25'b11101001_10101111_10011000_1;
      patterns[59826] = 25'b11101001_10110000_10011001_1;
      patterns[59827] = 25'b11101001_10110001_10011010_1;
      patterns[59828] = 25'b11101001_10110010_10011011_1;
      patterns[59829] = 25'b11101001_10110011_10011100_1;
      patterns[59830] = 25'b11101001_10110100_10011101_1;
      patterns[59831] = 25'b11101001_10110101_10011110_1;
      patterns[59832] = 25'b11101001_10110110_10011111_1;
      patterns[59833] = 25'b11101001_10110111_10100000_1;
      patterns[59834] = 25'b11101001_10111000_10100001_1;
      patterns[59835] = 25'b11101001_10111001_10100010_1;
      patterns[59836] = 25'b11101001_10111010_10100011_1;
      patterns[59837] = 25'b11101001_10111011_10100100_1;
      patterns[59838] = 25'b11101001_10111100_10100101_1;
      patterns[59839] = 25'b11101001_10111101_10100110_1;
      patterns[59840] = 25'b11101001_10111110_10100111_1;
      patterns[59841] = 25'b11101001_10111111_10101000_1;
      patterns[59842] = 25'b11101001_11000000_10101001_1;
      patterns[59843] = 25'b11101001_11000001_10101010_1;
      patterns[59844] = 25'b11101001_11000010_10101011_1;
      patterns[59845] = 25'b11101001_11000011_10101100_1;
      patterns[59846] = 25'b11101001_11000100_10101101_1;
      patterns[59847] = 25'b11101001_11000101_10101110_1;
      patterns[59848] = 25'b11101001_11000110_10101111_1;
      patterns[59849] = 25'b11101001_11000111_10110000_1;
      patterns[59850] = 25'b11101001_11001000_10110001_1;
      patterns[59851] = 25'b11101001_11001001_10110010_1;
      patterns[59852] = 25'b11101001_11001010_10110011_1;
      patterns[59853] = 25'b11101001_11001011_10110100_1;
      patterns[59854] = 25'b11101001_11001100_10110101_1;
      patterns[59855] = 25'b11101001_11001101_10110110_1;
      patterns[59856] = 25'b11101001_11001110_10110111_1;
      patterns[59857] = 25'b11101001_11001111_10111000_1;
      patterns[59858] = 25'b11101001_11010000_10111001_1;
      patterns[59859] = 25'b11101001_11010001_10111010_1;
      patterns[59860] = 25'b11101001_11010010_10111011_1;
      patterns[59861] = 25'b11101001_11010011_10111100_1;
      patterns[59862] = 25'b11101001_11010100_10111101_1;
      patterns[59863] = 25'b11101001_11010101_10111110_1;
      patterns[59864] = 25'b11101001_11010110_10111111_1;
      patterns[59865] = 25'b11101001_11010111_11000000_1;
      patterns[59866] = 25'b11101001_11011000_11000001_1;
      patterns[59867] = 25'b11101001_11011001_11000010_1;
      patterns[59868] = 25'b11101001_11011010_11000011_1;
      patterns[59869] = 25'b11101001_11011011_11000100_1;
      patterns[59870] = 25'b11101001_11011100_11000101_1;
      patterns[59871] = 25'b11101001_11011101_11000110_1;
      patterns[59872] = 25'b11101001_11011110_11000111_1;
      patterns[59873] = 25'b11101001_11011111_11001000_1;
      patterns[59874] = 25'b11101001_11100000_11001001_1;
      patterns[59875] = 25'b11101001_11100001_11001010_1;
      patterns[59876] = 25'b11101001_11100010_11001011_1;
      patterns[59877] = 25'b11101001_11100011_11001100_1;
      patterns[59878] = 25'b11101001_11100100_11001101_1;
      patterns[59879] = 25'b11101001_11100101_11001110_1;
      patterns[59880] = 25'b11101001_11100110_11001111_1;
      patterns[59881] = 25'b11101001_11100111_11010000_1;
      patterns[59882] = 25'b11101001_11101000_11010001_1;
      patterns[59883] = 25'b11101001_11101001_11010010_1;
      patterns[59884] = 25'b11101001_11101010_11010011_1;
      patterns[59885] = 25'b11101001_11101011_11010100_1;
      patterns[59886] = 25'b11101001_11101100_11010101_1;
      patterns[59887] = 25'b11101001_11101101_11010110_1;
      patterns[59888] = 25'b11101001_11101110_11010111_1;
      patterns[59889] = 25'b11101001_11101111_11011000_1;
      patterns[59890] = 25'b11101001_11110000_11011001_1;
      patterns[59891] = 25'b11101001_11110001_11011010_1;
      patterns[59892] = 25'b11101001_11110010_11011011_1;
      patterns[59893] = 25'b11101001_11110011_11011100_1;
      patterns[59894] = 25'b11101001_11110100_11011101_1;
      patterns[59895] = 25'b11101001_11110101_11011110_1;
      patterns[59896] = 25'b11101001_11110110_11011111_1;
      patterns[59897] = 25'b11101001_11110111_11100000_1;
      patterns[59898] = 25'b11101001_11111000_11100001_1;
      patterns[59899] = 25'b11101001_11111001_11100010_1;
      patterns[59900] = 25'b11101001_11111010_11100011_1;
      patterns[59901] = 25'b11101001_11111011_11100100_1;
      patterns[59902] = 25'b11101001_11111100_11100101_1;
      patterns[59903] = 25'b11101001_11111101_11100110_1;
      patterns[59904] = 25'b11101001_11111110_11100111_1;
      patterns[59905] = 25'b11101001_11111111_11101000_1;
      patterns[59906] = 25'b11101010_00000000_11101010_0;
      patterns[59907] = 25'b11101010_00000001_11101011_0;
      patterns[59908] = 25'b11101010_00000010_11101100_0;
      patterns[59909] = 25'b11101010_00000011_11101101_0;
      patterns[59910] = 25'b11101010_00000100_11101110_0;
      patterns[59911] = 25'b11101010_00000101_11101111_0;
      patterns[59912] = 25'b11101010_00000110_11110000_0;
      patterns[59913] = 25'b11101010_00000111_11110001_0;
      patterns[59914] = 25'b11101010_00001000_11110010_0;
      patterns[59915] = 25'b11101010_00001001_11110011_0;
      patterns[59916] = 25'b11101010_00001010_11110100_0;
      patterns[59917] = 25'b11101010_00001011_11110101_0;
      patterns[59918] = 25'b11101010_00001100_11110110_0;
      patterns[59919] = 25'b11101010_00001101_11110111_0;
      patterns[59920] = 25'b11101010_00001110_11111000_0;
      patterns[59921] = 25'b11101010_00001111_11111001_0;
      patterns[59922] = 25'b11101010_00010000_11111010_0;
      patterns[59923] = 25'b11101010_00010001_11111011_0;
      patterns[59924] = 25'b11101010_00010010_11111100_0;
      patterns[59925] = 25'b11101010_00010011_11111101_0;
      patterns[59926] = 25'b11101010_00010100_11111110_0;
      patterns[59927] = 25'b11101010_00010101_11111111_0;
      patterns[59928] = 25'b11101010_00010110_00000000_1;
      patterns[59929] = 25'b11101010_00010111_00000001_1;
      patterns[59930] = 25'b11101010_00011000_00000010_1;
      patterns[59931] = 25'b11101010_00011001_00000011_1;
      patterns[59932] = 25'b11101010_00011010_00000100_1;
      patterns[59933] = 25'b11101010_00011011_00000101_1;
      patterns[59934] = 25'b11101010_00011100_00000110_1;
      patterns[59935] = 25'b11101010_00011101_00000111_1;
      patterns[59936] = 25'b11101010_00011110_00001000_1;
      patterns[59937] = 25'b11101010_00011111_00001001_1;
      patterns[59938] = 25'b11101010_00100000_00001010_1;
      patterns[59939] = 25'b11101010_00100001_00001011_1;
      patterns[59940] = 25'b11101010_00100010_00001100_1;
      patterns[59941] = 25'b11101010_00100011_00001101_1;
      patterns[59942] = 25'b11101010_00100100_00001110_1;
      patterns[59943] = 25'b11101010_00100101_00001111_1;
      patterns[59944] = 25'b11101010_00100110_00010000_1;
      patterns[59945] = 25'b11101010_00100111_00010001_1;
      patterns[59946] = 25'b11101010_00101000_00010010_1;
      patterns[59947] = 25'b11101010_00101001_00010011_1;
      patterns[59948] = 25'b11101010_00101010_00010100_1;
      patterns[59949] = 25'b11101010_00101011_00010101_1;
      patterns[59950] = 25'b11101010_00101100_00010110_1;
      patterns[59951] = 25'b11101010_00101101_00010111_1;
      patterns[59952] = 25'b11101010_00101110_00011000_1;
      patterns[59953] = 25'b11101010_00101111_00011001_1;
      patterns[59954] = 25'b11101010_00110000_00011010_1;
      patterns[59955] = 25'b11101010_00110001_00011011_1;
      patterns[59956] = 25'b11101010_00110010_00011100_1;
      patterns[59957] = 25'b11101010_00110011_00011101_1;
      patterns[59958] = 25'b11101010_00110100_00011110_1;
      patterns[59959] = 25'b11101010_00110101_00011111_1;
      patterns[59960] = 25'b11101010_00110110_00100000_1;
      patterns[59961] = 25'b11101010_00110111_00100001_1;
      patterns[59962] = 25'b11101010_00111000_00100010_1;
      patterns[59963] = 25'b11101010_00111001_00100011_1;
      patterns[59964] = 25'b11101010_00111010_00100100_1;
      patterns[59965] = 25'b11101010_00111011_00100101_1;
      patterns[59966] = 25'b11101010_00111100_00100110_1;
      patterns[59967] = 25'b11101010_00111101_00100111_1;
      patterns[59968] = 25'b11101010_00111110_00101000_1;
      patterns[59969] = 25'b11101010_00111111_00101001_1;
      patterns[59970] = 25'b11101010_01000000_00101010_1;
      patterns[59971] = 25'b11101010_01000001_00101011_1;
      patterns[59972] = 25'b11101010_01000010_00101100_1;
      patterns[59973] = 25'b11101010_01000011_00101101_1;
      patterns[59974] = 25'b11101010_01000100_00101110_1;
      patterns[59975] = 25'b11101010_01000101_00101111_1;
      patterns[59976] = 25'b11101010_01000110_00110000_1;
      patterns[59977] = 25'b11101010_01000111_00110001_1;
      patterns[59978] = 25'b11101010_01001000_00110010_1;
      patterns[59979] = 25'b11101010_01001001_00110011_1;
      patterns[59980] = 25'b11101010_01001010_00110100_1;
      patterns[59981] = 25'b11101010_01001011_00110101_1;
      patterns[59982] = 25'b11101010_01001100_00110110_1;
      patterns[59983] = 25'b11101010_01001101_00110111_1;
      patterns[59984] = 25'b11101010_01001110_00111000_1;
      patterns[59985] = 25'b11101010_01001111_00111001_1;
      patterns[59986] = 25'b11101010_01010000_00111010_1;
      patterns[59987] = 25'b11101010_01010001_00111011_1;
      patterns[59988] = 25'b11101010_01010010_00111100_1;
      patterns[59989] = 25'b11101010_01010011_00111101_1;
      patterns[59990] = 25'b11101010_01010100_00111110_1;
      patterns[59991] = 25'b11101010_01010101_00111111_1;
      patterns[59992] = 25'b11101010_01010110_01000000_1;
      patterns[59993] = 25'b11101010_01010111_01000001_1;
      patterns[59994] = 25'b11101010_01011000_01000010_1;
      patterns[59995] = 25'b11101010_01011001_01000011_1;
      patterns[59996] = 25'b11101010_01011010_01000100_1;
      patterns[59997] = 25'b11101010_01011011_01000101_1;
      patterns[59998] = 25'b11101010_01011100_01000110_1;
      patterns[59999] = 25'b11101010_01011101_01000111_1;
      patterns[60000] = 25'b11101010_01011110_01001000_1;
      patterns[60001] = 25'b11101010_01011111_01001001_1;
      patterns[60002] = 25'b11101010_01100000_01001010_1;
      patterns[60003] = 25'b11101010_01100001_01001011_1;
      patterns[60004] = 25'b11101010_01100010_01001100_1;
      patterns[60005] = 25'b11101010_01100011_01001101_1;
      patterns[60006] = 25'b11101010_01100100_01001110_1;
      patterns[60007] = 25'b11101010_01100101_01001111_1;
      patterns[60008] = 25'b11101010_01100110_01010000_1;
      patterns[60009] = 25'b11101010_01100111_01010001_1;
      patterns[60010] = 25'b11101010_01101000_01010010_1;
      patterns[60011] = 25'b11101010_01101001_01010011_1;
      patterns[60012] = 25'b11101010_01101010_01010100_1;
      patterns[60013] = 25'b11101010_01101011_01010101_1;
      patterns[60014] = 25'b11101010_01101100_01010110_1;
      patterns[60015] = 25'b11101010_01101101_01010111_1;
      patterns[60016] = 25'b11101010_01101110_01011000_1;
      patterns[60017] = 25'b11101010_01101111_01011001_1;
      patterns[60018] = 25'b11101010_01110000_01011010_1;
      patterns[60019] = 25'b11101010_01110001_01011011_1;
      patterns[60020] = 25'b11101010_01110010_01011100_1;
      patterns[60021] = 25'b11101010_01110011_01011101_1;
      patterns[60022] = 25'b11101010_01110100_01011110_1;
      patterns[60023] = 25'b11101010_01110101_01011111_1;
      patterns[60024] = 25'b11101010_01110110_01100000_1;
      patterns[60025] = 25'b11101010_01110111_01100001_1;
      patterns[60026] = 25'b11101010_01111000_01100010_1;
      patterns[60027] = 25'b11101010_01111001_01100011_1;
      patterns[60028] = 25'b11101010_01111010_01100100_1;
      patterns[60029] = 25'b11101010_01111011_01100101_1;
      patterns[60030] = 25'b11101010_01111100_01100110_1;
      patterns[60031] = 25'b11101010_01111101_01100111_1;
      patterns[60032] = 25'b11101010_01111110_01101000_1;
      patterns[60033] = 25'b11101010_01111111_01101001_1;
      patterns[60034] = 25'b11101010_10000000_01101010_1;
      patterns[60035] = 25'b11101010_10000001_01101011_1;
      patterns[60036] = 25'b11101010_10000010_01101100_1;
      patterns[60037] = 25'b11101010_10000011_01101101_1;
      patterns[60038] = 25'b11101010_10000100_01101110_1;
      patterns[60039] = 25'b11101010_10000101_01101111_1;
      patterns[60040] = 25'b11101010_10000110_01110000_1;
      patterns[60041] = 25'b11101010_10000111_01110001_1;
      patterns[60042] = 25'b11101010_10001000_01110010_1;
      patterns[60043] = 25'b11101010_10001001_01110011_1;
      patterns[60044] = 25'b11101010_10001010_01110100_1;
      patterns[60045] = 25'b11101010_10001011_01110101_1;
      patterns[60046] = 25'b11101010_10001100_01110110_1;
      patterns[60047] = 25'b11101010_10001101_01110111_1;
      patterns[60048] = 25'b11101010_10001110_01111000_1;
      patterns[60049] = 25'b11101010_10001111_01111001_1;
      patterns[60050] = 25'b11101010_10010000_01111010_1;
      patterns[60051] = 25'b11101010_10010001_01111011_1;
      patterns[60052] = 25'b11101010_10010010_01111100_1;
      patterns[60053] = 25'b11101010_10010011_01111101_1;
      patterns[60054] = 25'b11101010_10010100_01111110_1;
      patterns[60055] = 25'b11101010_10010101_01111111_1;
      patterns[60056] = 25'b11101010_10010110_10000000_1;
      patterns[60057] = 25'b11101010_10010111_10000001_1;
      patterns[60058] = 25'b11101010_10011000_10000010_1;
      patterns[60059] = 25'b11101010_10011001_10000011_1;
      patterns[60060] = 25'b11101010_10011010_10000100_1;
      patterns[60061] = 25'b11101010_10011011_10000101_1;
      patterns[60062] = 25'b11101010_10011100_10000110_1;
      patterns[60063] = 25'b11101010_10011101_10000111_1;
      patterns[60064] = 25'b11101010_10011110_10001000_1;
      patterns[60065] = 25'b11101010_10011111_10001001_1;
      patterns[60066] = 25'b11101010_10100000_10001010_1;
      patterns[60067] = 25'b11101010_10100001_10001011_1;
      patterns[60068] = 25'b11101010_10100010_10001100_1;
      patterns[60069] = 25'b11101010_10100011_10001101_1;
      patterns[60070] = 25'b11101010_10100100_10001110_1;
      patterns[60071] = 25'b11101010_10100101_10001111_1;
      patterns[60072] = 25'b11101010_10100110_10010000_1;
      patterns[60073] = 25'b11101010_10100111_10010001_1;
      patterns[60074] = 25'b11101010_10101000_10010010_1;
      patterns[60075] = 25'b11101010_10101001_10010011_1;
      patterns[60076] = 25'b11101010_10101010_10010100_1;
      patterns[60077] = 25'b11101010_10101011_10010101_1;
      patterns[60078] = 25'b11101010_10101100_10010110_1;
      patterns[60079] = 25'b11101010_10101101_10010111_1;
      patterns[60080] = 25'b11101010_10101110_10011000_1;
      patterns[60081] = 25'b11101010_10101111_10011001_1;
      patterns[60082] = 25'b11101010_10110000_10011010_1;
      patterns[60083] = 25'b11101010_10110001_10011011_1;
      patterns[60084] = 25'b11101010_10110010_10011100_1;
      patterns[60085] = 25'b11101010_10110011_10011101_1;
      patterns[60086] = 25'b11101010_10110100_10011110_1;
      patterns[60087] = 25'b11101010_10110101_10011111_1;
      patterns[60088] = 25'b11101010_10110110_10100000_1;
      patterns[60089] = 25'b11101010_10110111_10100001_1;
      patterns[60090] = 25'b11101010_10111000_10100010_1;
      patterns[60091] = 25'b11101010_10111001_10100011_1;
      patterns[60092] = 25'b11101010_10111010_10100100_1;
      patterns[60093] = 25'b11101010_10111011_10100101_1;
      patterns[60094] = 25'b11101010_10111100_10100110_1;
      patterns[60095] = 25'b11101010_10111101_10100111_1;
      patterns[60096] = 25'b11101010_10111110_10101000_1;
      patterns[60097] = 25'b11101010_10111111_10101001_1;
      patterns[60098] = 25'b11101010_11000000_10101010_1;
      patterns[60099] = 25'b11101010_11000001_10101011_1;
      patterns[60100] = 25'b11101010_11000010_10101100_1;
      patterns[60101] = 25'b11101010_11000011_10101101_1;
      patterns[60102] = 25'b11101010_11000100_10101110_1;
      patterns[60103] = 25'b11101010_11000101_10101111_1;
      patterns[60104] = 25'b11101010_11000110_10110000_1;
      patterns[60105] = 25'b11101010_11000111_10110001_1;
      patterns[60106] = 25'b11101010_11001000_10110010_1;
      patterns[60107] = 25'b11101010_11001001_10110011_1;
      patterns[60108] = 25'b11101010_11001010_10110100_1;
      patterns[60109] = 25'b11101010_11001011_10110101_1;
      patterns[60110] = 25'b11101010_11001100_10110110_1;
      patterns[60111] = 25'b11101010_11001101_10110111_1;
      patterns[60112] = 25'b11101010_11001110_10111000_1;
      patterns[60113] = 25'b11101010_11001111_10111001_1;
      patterns[60114] = 25'b11101010_11010000_10111010_1;
      patterns[60115] = 25'b11101010_11010001_10111011_1;
      patterns[60116] = 25'b11101010_11010010_10111100_1;
      patterns[60117] = 25'b11101010_11010011_10111101_1;
      patterns[60118] = 25'b11101010_11010100_10111110_1;
      patterns[60119] = 25'b11101010_11010101_10111111_1;
      patterns[60120] = 25'b11101010_11010110_11000000_1;
      patterns[60121] = 25'b11101010_11010111_11000001_1;
      patterns[60122] = 25'b11101010_11011000_11000010_1;
      patterns[60123] = 25'b11101010_11011001_11000011_1;
      patterns[60124] = 25'b11101010_11011010_11000100_1;
      patterns[60125] = 25'b11101010_11011011_11000101_1;
      patterns[60126] = 25'b11101010_11011100_11000110_1;
      patterns[60127] = 25'b11101010_11011101_11000111_1;
      patterns[60128] = 25'b11101010_11011110_11001000_1;
      patterns[60129] = 25'b11101010_11011111_11001001_1;
      patterns[60130] = 25'b11101010_11100000_11001010_1;
      patterns[60131] = 25'b11101010_11100001_11001011_1;
      patterns[60132] = 25'b11101010_11100010_11001100_1;
      patterns[60133] = 25'b11101010_11100011_11001101_1;
      patterns[60134] = 25'b11101010_11100100_11001110_1;
      patterns[60135] = 25'b11101010_11100101_11001111_1;
      patterns[60136] = 25'b11101010_11100110_11010000_1;
      patterns[60137] = 25'b11101010_11100111_11010001_1;
      patterns[60138] = 25'b11101010_11101000_11010010_1;
      patterns[60139] = 25'b11101010_11101001_11010011_1;
      patterns[60140] = 25'b11101010_11101010_11010100_1;
      patterns[60141] = 25'b11101010_11101011_11010101_1;
      patterns[60142] = 25'b11101010_11101100_11010110_1;
      patterns[60143] = 25'b11101010_11101101_11010111_1;
      patterns[60144] = 25'b11101010_11101110_11011000_1;
      patterns[60145] = 25'b11101010_11101111_11011001_1;
      patterns[60146] = 25'b11101010_11110000_11011010_1;
      patterns[60147] = 25'b11101010_11110001_11011011_1;
      patterns[60148] = 25'b11101010_11110010_11011100_1;
      patterns[60149] = 25'b11101010_11110011_11011101_1;
      patterns[60150] = 25'b11101010_11110100_11011110_1;
      patterns[60151] = 25'b11101010_11110101_11011111_1;
      patterns[60152] = 25'b11101010_11110110_11100000_1;
      patterns[60153] = 25'b11101010_11110111_11100001_1;
      patterns[60154] = 25'b11101010_11111000_11100010_1;
      patterns[60155] = 25'b11101010_11111001_11100011_1;
      patterns[60156] = 25'b11101010_11111010_11100100_1;
      patterns[60157] = 25'b11101010_11111011_11100101_1;
      patterns[60158] = 25'b11101010_11111100_11100110_1;
      patterns[60159] = 25'b11101010_11111101_11100111_1;
      patterns[60160] = 25'b11101010_11111110_11101000_1;
      patterns[60161] = 25'b11101010_11111111_11101001_1;
      patterns[60162] = 25'b11101011_00000000_11101011_0;
      patterns[60163] = 25'b11101011_00000001_11101100_0;
      patterns[60164] = 25'b11101011_00000010_11101101_0;
      patterns[60165] = 25'b11101011_00000011_11101110_0;
      patterns[60166] = 25'b11101011_00000100_11101111_0;
      patterns[60167] = 25'b11101011_00000101_11110000_0;
      patterns[60168] = 25'b11101011_00000110_11110001_0;
      patterns[60169] = 25'b11101011_00000111_11110010_0;
      patterns[60170] = 25'b11101011_00001000_11110011_0;
      patterns[60171] = 25'b11101011_00001001_11110100_0;
      patterns[60172] = 25'b11101011_00001010_11110101_0;
      patterns[60173] = 25'b11101011_00001011_11110110_0;
      patterns[60174] = 25'b11101011_00001100_11110111_0;
      patterns[60175] = 25'b11101011_00001101_11111000_0;
      patterns[60176] = 25'b11101011_00001110_11111001_0;
      patterns[60177] = 25'b11101011_00001111_11111010_0;
      patterns[60178] = 25'b11101011_00010000_11111011_0;
      patterns[60179] = 25'b11101011_00010001_11111100_0;
      patterns[60180] = 25'b11101011_00010010_11111101_0;
      patterns[60181] = 25'b11101011_00010011_11111110_0;
      patterns[60182] = 25'b11101011_00010100_11111111_0;
      patterns[60183] = 25'b11101011_00010101_00000000_1;
      patterns[60184] = 25'b11101011_00010110_00000001_1;
      patterns[60185] = 25'b11101011_00010111_00000010_1;
      patterns[60186] = 25'b11101011_00011000_00000011_1;
      patterns[60187] = 25'b11101011_00011001_00000100_1;
      patterns[60188] = 25'b11101011_00011010_00000101_1;
      patterns[60189] = 25'b11101011_00011011_00000110_1;
      patterns[60190] = 25'b11101011_00011100_00000111_1;
      patterns[60191] = 25'b11101011_00011101_00001000_1;
      patterns[60192] = 25'b11101011_00011110_00001001_1;
      patterns[60193] = 25'b11101011_00011111_00001010_1;
      patterns[60194] = 25'b11101011_00100000_00001011_1;
      patterns[60195] = 25'b11101011_00100001_00001100_1;
      patterns[60196] = 25'b11101011_00100010_00001101_1;
      patterns[60197] = 25'b11101011_00100011_00001110_1;
      patterns[60198] = 25'b11101011_00100100_00001111_1;
      patterns[60199] = 25'b11101011_00100101_00010000_1;
      patterns[60200] = 25'b11101011_00100110_00010001_1;
      patterns[60201] = 25'b11101011_00100111_00010010_1;
      patterns[60202] = 25'b11101011_00101000_00010011_1;
      patterns[60203] = 25'b11101011_00101001_00010100_1;
      patterns[60204] = 25'b11101011_00101010_00010101_1;
      patterns[60205] = 25'b11101011_00101011_00010110_1;
      patterns[60206] = 25'b11101011_00101100_00010111_1;
      patterns[60207] = 25'b11101011_00101101_00011000_1;
      patterns[60208] = 25'b11101011_00101110_00011001_1;
      patterns[60209] = 25'b11101011_00101111_00011010_1;
      patterns[60210] = 25'b11101011_00110000_00011011_1;
      patterns[60211] = 25'b11101011_00110001_00011100_1;
      patterns[60212] = 25'b11101011_00110010_00011101_1;
      patterns[60213] = 25'b11101011_00110011_00011110_1;
      patterns[60214] = 25'b11101011_00110100_00011111_1;
      patterns[60215] = 25'b11101011_00110101_00100000_1;
      patterns[60216] = 25'b11101011_00110110_00100001_1;
      patterns[60217] = 25'b11101011_00110111_00100010_1;
      patterns[60218] = 25'b11101011_00111000_00100011_1;
      patterns[60219] = 25'b11101011_00111001_00100100_1;
      patterns[60220] = 25'b11101011_00111010_00100101_1;
      patterns[60221] = 25'b11101011_00111011_00100110_1;
      patterns[60222] = 25'b11101011_00111100_00100111_1;
      patterns[60223] = 25'b11101011_00111101_00101000_1;
      patterns[60224] = 25'b11101011_00111110_00101001_1;
      patterns[60225] = 25'b11101011_00111111_00101010_1;
      patterns[60226] = 25'b11101011_01000000_00101011_1;
      patterns[60227] = 25'b11101011_01000001_00101100_1;
      patterns[60228] = 25'b11101011_01000010_00101101_1;
      patterns[60229] = 25'b11101011_01000011_00101110_1;
      patterns[60230] = 25'b11101011_01000100_00101111_1;
      patterns[60231] = 25'b11101011_01000101_00110000_1;
      patterns[60232] = 25'b11101011_01000110_00110001_1;
      patterns[60233] = 25'b11101011_01000111_00110010_1;
      patterns[60234] = 25'b11101011_01001000_00110011_1;
      patterns[60235] = 25'b11101011_01001001_00110100_1;
      patterns[60236] = 25'b11101011_01001010_00110101_1;
      patterns[60237] = 25'b11101011_01001011_00110110_1;
      patterns[60238] = 25'b11101011_01001100_00110111_1;
      patterns[60239] = 25'b11101011_01001101_00111000_1;
      patterns[60240] = 25'b11101011_01001110_00111001_1;
      patterns[60241] = 25'b11101011_01001111_00111010_1;
      patterns[60242] = 25'b11101011_01010000_00111011_1;
      patterns[60243] = 25'b11101011_01010001_00111100_1;
      patterns[60244] = 25'b11101011_01010010_00111101_1;
      patterns[60245] = 25'b11101011_01010011_00111110_1;
      patterns[60246] = 25'b11101011_01010100_00111111_1;
      patterns[60247] = 25'b11101011_01010101_01000000_1;
      patterns[60248] = 25'b11101011_01010110_01000001_1;
      patterns[60249] = 25'b11101011_01010111_01000010_1;
      patterns[60250] = 25'b11101011_01011000_01000011_1;
      patterns[60251] = 25'b11101011_01011001_01000100_1;
      patterns[60252] = 25'b11101011_01011010_01000101_1;
      patterns[60253] = 25'b11101011_01011011_01000110_1;
      patterns[60254] = 25'b11101011_01011100_01000111_1;
      patterns[60255] = 25'b11101011_01011101_01001000_1;
      patterns[60256] = 25'b11101011_01011110_01001001_1;
      patterns[60257] = 25'b11101011_01011111_01001010_1;
      patterns[60258] = 25'b11101011_01100000_01001011_1;
      patterns[60259] = 25'b11101011_01100001_01001100_1;
      patterns[60260] = 25'b11101011_01100010_01001101_1;
      patterns[60261] = 25'b11101011_01100011_01001110_1;
      patterns[60262] = 25'b11101011_01100100_01001111_1;
      patterns[60263] = 25'b11101011_01100101_01010000_1;
      patterns[60264] = 25'b11101011_01100110_01010001_1;
      patterns[60265] = 25'b11101011_01100111_01010010_1;
      patterns[60266] = 25'b11101011_01101000_01010011_1;
      patterns[60267] = 25'b11101011_01101001_01010100_1;
      patterns[60268] = 25'b11101011_01101010_01010101_1;
      patterns[60269] = 25'b11101011_01101011_01010110_1;
      patterns[60270] = 25'b11101011_01101100_01010111_1;
      patterns[60271] = 25'b11101011_01101101_01011000_1;
      patterns[60272] = 25'b11101011_01101110_01011001_1;
      patterns[60273] = 25'b11101011_01101111_01011010_1;
      patterns[60274] = 25'b11101011_01110000_01011011_1;
      patterns[60275] = 25'b11101011_01110001_01011100_1;
      patterns[60276] = 25'b11101011_01110010_01011101_1;
      patterns[60277] = 25'b11101011_01110011_01011110_1;
      patterns[60278] = 25'b11101011_01110100_01011111_1;
      patterns[60279] = 25'b11101011_01110101_01100000_1;
      patterns[60280] = 25'b11101011_01110110_01100001_1;
      patterns[60281] = 25'b11101011_01110111_01100010_1;
      patterns[60282] = 25'b11101011_01111000_01100011_1;
      patterns[60283] = 25'b11101011_01111001_01100100_1;
      patterns[60284] = 25'b11101011_01111010_01100101_1;
      patterns[60285] = 25'b11101011_01111011_01100110_1;
      patterns[60286] = 25'b11101011_01111100_01100111_1;
      patterns[60287] = 25'b11101011_01111101_01101000_1;
      patterns[60288] = 25'b11101011_01111110_01101001_1;
      patterns[60289] = 25'b11101011_01111111_01101010_1;
      patterns[60290] = 25'b11101011_10000000_01101011_1;
      patterns[60291] = 25'b11101011_10000001_01101100_1;
      patterns[60292] = 25'b11101011_10000010_01101101_1;
      patterns[60293] = 25'b11101011_10000011_01101110_1;
      patterns[60294] = 25'b11101011_10000100_01101111_1;
      patterns[60295] = 25'b11101011_10000101_01110000_1;
      patterns[60296] = 25'b11101011_10000110_01110001_1;
      patterns[60297] = 25'b11101011_10000111_01110010_1;
      patterns[60298] = 25'b11101011_10001000_01110011_1;
      patterns[60299] = 25'b11101011_10001001_01110100_1;
      patterns[60300] = 25'b11101011_10001010_01110101_1;
      patterns[60301] = 25'b11101011_10001011_01110110_1;
      patterns[60302] = 25'b11101011_10001100_01110111_1;
      patterns[60303] = 25'b11101011_10001101_01111000_1;
      patterns[60304] = 25'b11101011_10001110_01111001_1;
      patterns[60305] = 25'b11101011_10001111_01111010_1;
      patterns[60306] = 25'b11101011_10010000_01111011_1;
      patterns[60307] = 25'b11101011_10010001_01111100_1;
      patterns[60308] = 25'b11101011_10010010_01111101_1;
      patterns[60309] = 25'b11101011_10010011_01111110_1;
      patterns[60310] = 25'b11101011_10010100_01111111_1;
      patterns[60311] = 25'b11101011_10010101_10000000_1;
      patterns[60312] = 25'b11101011_10010110_10000001_1;
      patterns[60313] = 25'b11101011_10010111_10000010_1;
      patterns[60314] = 25'b11101011_10011000_10000011_1;
      patterns[60315] = 25'b11101011_10011001_10000100_1;
      patterns[60316] = 25'b11101011_10011010_10000101_1;
      patterns[60317] = 25'b11101011_10011011_10000110_1;
      patterns[60318] = 25'b11101011_10011100_10000111_1;
      patterns[60319] = 25'b11101011_10011101_10001000_1;
      patterns[60320] = 25'b11101011_10011110_10001001_1;
      patterns[60321] = 25'b11101011_10011111_10001010_1;
      patterns[60322] = 25'b11101011_10100000_10001011_1;
      patterns[60323] = 25'b11101011_10100001_10001100_1;
      patterns[60324] = 25'b11101011_10100010_10001101_1;
      patterns[60325] = 25'b11101011_10100011_10001110_1;
      patterns[60326] = 25'b11101011_10100100_10001111_1;
      patterns[60327] = 25'b11101011_10100101_10010000_1;
      patterns[60328] = 25'b11101011_10100110_10010001_1;
      patterns[60329] = 25'b11101011_10100111_10010010_1;
      patterns[60330] = 25'b11101011_10101000_10010011_1;
      patterns[60331] = 25'b11101011_10101001_10010100_1;
      patterns[60332] = 25'b11101011_10101010_10010101_1;
      patterns[60333] = 25'b11101011_10101011_10010110_1;
      patterns[60334] = 25'b11101011_10101100_10010111_1;
      patterns[60335] = 25'b11101011_10101101_10011000_1;
      patterns[60336] = 25'b11101011_10101110_10011001_1;
      patterns[60337] = 25'b11101011_10101111_10011010_1;
      patterns[60338] = 25'b11101011_10110000_10011011_1;
      patterns[60339] = 25'b11101011_10110001_10011100_1;
      patterns[60340] = 25'b11101011_10110010_10011101_1;
      patterns[60341] = 25'b11101011_10110011_10011110_1;
      patterns[60342] = 25'b11101011_10110100_10011111_1;
      patterns[60343] = 25'b11101011_10110101_10100000_1;
      patterns[60344] = 25'b11101011_10110110_10100001_1;
      patterns[60345] = 25'b11101011_10110111_10100010_1;
      patterns[60346] = 25'b11101011_10111000_10100011_1;
      patterns[60347] = 25'b11101011_10111001_10100100_1;
      patterns[60348] = 25'b11101011_10111010_10100101_1;
      patterns[60349] = 25'b11101011_10111011_10100110_1;
      patterns[60350] = 25'b11101011_10111100_10100111_1;
      patterns[60351] = 25'b11101011_10111101_10101000_1;
      patterns[60352] = 25'b11101011_10111110_10101001_1;
      patterns[60353] = 25'b11101011_10111111_10101010_1;
      patterns[60354] = 25'b11101011_11000000_10101011_1;
      patterns[60355] = 25'b11101011_11000001_10101100_1;
      patterns[60356] = 25'b11101011_11000010_10101101_1;
      patterns[60357] = 25'b11101011_11000011_10101110_1;
      patterns[60358] = 25'b11101011_11000100_10101111_1;
      patterns[60359] = 25'b11101011_11000101_10110000_1;
      patterns[60360] = 25'b11101011_11000110_10110001_1;
      patterns[60361] = 25'b11101011_11000111_10110010_1;
      patterns[60362] = 25'b11101011_11001000_10110011_1;
      patterns[60363] = 25'b11101011_11001001_10110100_1;
      patterns[60364] = 25'b11101011_11001010_10110101_1;
      patterns[60365] = 25'b11101011_11001011_10110110_1;
      patterns[60366] = 25'b11101011_11001100_10110111_1;
      patterns[60367] = 25'b11101011_11001101_10111000_1;
      patterns[60368] = 25'b11101011_11001110_10111001_1;
      patterns[60369] = 25'b11101011_11001111_10111010_1;
      patterns[60370] = 25'b11101011_11010000_10111011_1;
      patterns[60371] = 25'b11101011_11010001_10111100_1;
      patterns[60372] = 25'b11101011_11010010_10111101_1;
      patterns[60373] = 25'b11101011_11010011_10111110_1;
      patterns[60374] = 25'b11101011_11010100_10111111_1;
      patterns[60375] = 25'b11101011_11010101_11000000_1;
      patterns[60376] = 25'b11101011_11010110_11000001_1;
      patterns[60377] = 25'b11101011_11010111_11000010_1;
      patterns[60378] = 25'b11101011_11011000_11000011_1;
      patterns[60379] = 25'b11101011_11011001_11000100_1;
      patterns[60380] = 25'b11101011_11011010_11000101_1;
      patterns[60381] = 25'b11101011_11011011_11000110_1;
      patterns[60382] = 25'b11101011_11011100_11000111_1;
      patterns[60383] = 25'b11101011_11011101_11001000_1;
      patterns[60384] = 25'b11101011_11011110_11001001_1;
      patterns[60385] = 25'b11101011_11011111_11001010_1;
      patterns[60386] = 25'b11101011_11100000_11001011_1;
      patterns[60387] = 25'b11101011_11100001_11001100_1;
      patterns[60388] = 25'b11101011_11100010_11001101_1;
      patterns[60389] = 25'b11101011_11100011_11001110_1;
      patterns[60390] = 25'b11101011_11100100_11001111_1;
      patterns[60391] = 25'b11101011_11100101_11010000_1;
      patterns[60392] = 25'b11101011_11100110_11010001_1;
      patterns[60393] = 25'b11101011_11100111_11010010_1;
      patterns[60394] = 25'b11101011_11101000_11010011_1;
      patterns[60395] = 25'b11101011_11101001_11010100_1;
      patterns[60396] = 25'b11101011_11101010_11010101_1;
      patterns[60397] = 25'b11101011_11101011_11010110_1;
      patterns[60398] = 25'b11101011_11101100_11010111_1;
      patterns[60399] = 25'b11101011_11101101_11011000_1;
      patterns[60400] = 25'b11101011_11101110_11011001_1;
      patterns[60401] = 25'b11101011_11101111_11011010_1;
      patterns[60402] = 25'b11101011_11110000_11011011_1;
      patterns[60403] = 25'b11101011_11110001_11011100_1;
      patterns[60404] = 25'b11101011_11110010_11011101_1;
      patterns[60405] = 25'b11101011_11110011_11011110_1;
      patterns[60406] = 25'b11101011_11110100_11011111_1;
      patterns[60407] = 25'b11101011_11110101_11100000_1;
      patterns[60408] = 25'b11101011_11110110_11100001_1;
      patterns[60409] = 25'b11101011_11110111_11100010_1;
      patterns[60410] = 25'b11101011_11111000_11100011_1;
      patterns[60411] = 25'b11101011_11111001_11100100_1;
      patterns[60412] = 25'b11101011_11111010_11100101_1;
      patterns[60413] = 25'b11101011_11111011_11100110_1;
      patterns[60414] = 25'b11101011_11111100_11100111_1;
      patterns[60415] = 25'b11101011_11111101_11101000_1;
      patterns[60416] = 25'b11101011_11111110_11101001_1;
      patterns[60417] = 25'b11101011_11111111_11101010_1;
      patterns[60418] = 25'b11101100_00000000_11101100_0;
      patterns[60419] = 25'b11101100_00000001_11101101_0;
      patterns[60420] = 25'b11101100_00000010_11101110_0;
      patterns[60421] = 25'b11101100_00000011_11101111_0;
      patterns[60422] = 25'b11101100_00000100_11110000_0;
      patterns[60423] = 25'b11101100_00000101_11110001_0;
      patterns[60424] = 25'b11101100_00000110_11110010_0;
      patterns[60425] = 25'b11101100_00000111_11110011_0;
      patterns[60426] = 25'b11101100_00001000_11110100_0;
      patterns[60427] = 25'b11101100_00001001_11110101_0;
      patterns[60428] = 25'b11101100_00001010_11110110_0;
      patterns[60429] = 25'b11101100_00001011_11110111_0;
      patterns[60430] = 25'b11101100_00001100_11111000_0;
      patterns[60431] = 25'b11101100_00001101_11111001_0;
      patterns[60432] = 25'b11101100_00001110_11111010_0;
      patterns[60433] = 25'b11101100_00001111_11111011_0;
      patterns[60434] = 25'b11101100_00010000_11111100_0;
      patterns[60435] = 25'b11101100_00010001_11111101_0;
      patterns[60436] = 25'b11101100_00010010_11111110_0;
      patterns[60437] = 25'b11101100_00010011_11111111_0;
      patterns[60438] = 25'b11101100_00010100_00000000_1;
      patterns[60439] = 25'b11101100_00010101_00000001_1;
      patterns[60440] = 25'b11101100_00010110_00000010_1;
      patterns[60441] = 25'b11101100_00010111_00000011_1;
      patterns[60442] = 25'b11101100_00011000_00000100_1;
      patterns[60443] = 25'b11101100_00011001_00000101_1;
      patterns[60444] = 25'b11101100_00011010_00000110_1;
      patterns[60445] = 25'b11101100_00011011_00000111_1;
      patterns[60446] = 25'b11101100_00011100_00001000_1;
      patterns[60447] = 25'b11101100_00011101_00001001_1;
      patterns[60448] = 25'b11101100_00011110_00001010_1;
      patterns[60449] = 25'b11101100_00011111_00001011_1;
      patterns[60450] = 25'b11101100_00100000_00001100_1;
      patterns[60451] = 25'b11101100_00100001_00001101_1;
      patterns[60452] = 25'b11101100_00100010_00001110_1;
      patterns[60453] = 25'b11101100_00100011_00001111_1;
      patterns[60454] = 25'b11101100_00100100_00010000_1;
      patterns[60455] = 25'b11101100_00100101_00010001_1;
      patterns[60456] = 25'b11101100_00100110_00010010_1;
      patterns[60457] = 25'b11101100_00100111_00010011_1;
      patterns[60458] = 25'b11101100_00101000_00010100_1;
      patterns[60459] = 25'b11101100_00101001_00010101_1;
      patterns[60460] = 25'b11101100_00101010_00010110_1;
      patterns[60461] = 25'b11101100_00101011_00010111_1;
      patterns[60462] = 25'b11101100_00101100_00011000_1;
      patterns[60463] = 25'b11101100_00101101_00011001_1;
      patterns[60464] = 25'b11101100_00101110_00011010_1;
      patterns[60465] = 25'b11101100_00101111_00011011_1;
      patterns[60466] = 25'b11101100_00110000_00011100_1;
      patterns[60467] = 25'b11101100_00110001_00011101_1;
      patterns[60468] = 25'b11101100_00110010_00011110_1;
      patterns[60469] = 25'b11101100_00110011_00011111_1;
      patterns[60470] = 25'b11101100_00110100_00100000_1;
      patterns[60471] = 25'b11101100_00110101_00100001_1;
      patterns[60472] = 25'b11101100_00110110_00100010_1;
      patterns[60473] = 25'b11101100_00110111_00100011_1;
      patterns[60474] = 25'b11101100_00111000_00100100_1;
      patterns[60475] = 25'b11101100_00111001_00100101_1;
      patterns[60476] = 25'b11101100_00111010_00100110_1;
      patterns[60477] = 25'b11101100_00111011_00100111_1;
      patterns[60478] = 25'b11101100_00111100_00101000_1;
      patterns[60479] = 25'b11101100_00111101_00101001_1;
      patterns[60480] = 25'b11101100_00111110_00101010_1;
      patterns[60481] = 25'b11101100_00111111_00101011_1;
      patterns[60482] = 25'b11101100_01000000_00101100_1;
      patterns[60483] = 25'b11101100_01000001_00101101_1;
      patterns[60484] = 25'b11101100_01000010_00101110_1;
      patterns[60485] = 25'b11101100_01000011_00101111_1;
      patterns[60486] = 25'b11101100_01000100_00110000_1;
      patterns[60487] = 25'b11101100_01000101_00110001_1;
      patterns[60488] = 25'b11101100_01000110_00110010_1;
      patterns[60489] = 25'b11101100_01000111_00110011_1;
      patterns[60490] = 25'b11101100_01001000_00110100_1;
      patterns[60491] = 25'b11101100_01001001_00110101_1;
      patterns[60492] = 25'b11101100_01001010_00110110_1;
      patterns[60493] = 25'b11101100_01001011_00110111_1;
      patterns[60494] = 25'b11101100_01001100_00111000_1;
      patterns[60495] = 25'b11101100_01001101_00111001_1;
      patterns[60496] = 25'b11101100_01001110_00111010_1;
      patterns[60497] = 25'b11101100_01001111_00111011_1;
      patterns[60498] = 25'b11101100_01010000_00111100_1;
      patterns[60499] = 25'b11101100_01010001_00111101_1;
      patterns[60500] = 25'b11101100_01010010_00111110_1;
      patterns[60501] = 25'b11101100_01010011_00111111_1;
      patterns[60502] = 25'b11101100_01010100_01000000_1;
      patterns[60503] = 25'b11101100_01010101_01000001_1;
      patterns[60504] = 25'b11101100_01010110_01000010_1;
      patterns[60505] = 25'b11101100_01010111_01000011_1;
      patterns[60506] = 25'b11101100_01011000_01000100_1;
      patterns[60507] = 25'b11101100_01011001_01000101_1;
      patterns[60508] = 25'b11101100_01011010_01000110_1;
      patterns[60509] = 25'b11101100_01011011_01000111_1;
      patterns[60510] = 25'b11101100_01011100_01001000_1;
      patterns[60511] = 25'b11101100_01011101_01001001_1;
      patterns[60512] = 25'b11101100_01011110_01001010_1;
      patterns[60513] = 25'b11101100_01011111_01001011_1;
      patterns[60514] = 25'b11101100_01100000_01001100_1;
      patterns[60515] = 25'b11101100_01100001_01001101_1;
      patterns[60516] = 25'b11101100_01100010_01001110_1;
      patterns[60517] = 25'b11101100_01100011_01001111_1;
      patterns[60518] = 25'b11101100_01100100_01010000_1;
      patterns[60519] = 25'b11101100_01100101_01010001_1;
      patterns[60520] = 25'b11101100_01100110_01010010_1;
      patterns[60521] = 25'b11101100_01100111_01010011_1;
      patterns[60522] = 25'b11101100_01101000_01010100_1;
      patterns[60523] = 25'b11101100_01101001_01010101_1;
      patterns[60524] = 25'b11101100_01101010_01010110_1;
      patterns[60525] = 25'b11101100_01101011_01010111_1;
      patterns[60526] = 25'b11101100_01101100_01011000_1;
      patterns[60527] = 25'b11101100_01101101_01011001_1;
      patterns[60528] = 25'b11101100_01101110_01011010_1;
      patterns[60529] = 25'b11101100_01101111_01011011_1;
      patterns[60530] = 25'b11101100_01110000_01011100_1;
      patterns[60531] = 25'b11101100_01110001_01011101_1;
      patterns[60532] = 25'b11101100_01110010_01011110_1;
      patterns[60533] = 25'b11101100_01110011_01011111_1;
      patterns[60534] = 25'b11101100_01110100_01100000_1;
      patterns[60535] = 25'b11101100_01110101_01100001_1;
      patterns[60536] = 25'b11101100_01110110_01100010_1;
      patterns[60537] = 25'b11101100_01110111_01100011_1;
      patterns[60538] = 25'b11101100_01111000_01100100_1;
      patterns[60539] = 25'b11101100_01111001_01100101_1;
      patterns[60540] = 25'b11101100_01111010_01100110_1;
      patterns[60541] = 25'b11101100_01111011_01100111_1;
      patterns[60542] = 25'b11101100_01111100_01101000_1;
      patterns[60543] = 25'b11101100_01111101_01101001_1;
      patterns[60544] = 25'b11101100_01111110_01101010_1;
      patterns[60545] = 25'b11101100_01111111_01101011_1;
      patterns[60546] = 25'b11101100_10000000_01101100_1;
      patterns[60547] = 25'b11101100_10000001_01101101_1;
      patterns[60548] = 25'b11101100_10000010_01101110_1;
      patterns[60549] = 25'b11101100_10000011_01101111_1;
      patterns[60550] = 25'b11101100_10000100_01110000_1;
      patterns[60551] = 25'b11101100_10000101_01110001_1;
      patterns[60552] = 25'b11101100_10000110_01110010_1;
      patterns[60553] = 25'b11101100_10000111_01110011_1;
      patterns[60554] = 25'b11101100_10001000_01110100_1;
      patterns[60555] = 25'b11101100_10001001_01110101_1;
      patterns[60556] = 25'b11101100_10001010_01110110_1;
      patterns[60557] = 25'b11101100_10001011_01110111_1;
      patterns[60558] = 25'b11101100_10001100_01111000_1;
      patterns[60559] = 25'b11101100_10001101_01111001_1;
      patterns[60560] = 25'b11101100_10001110_01111010_1;
      patterns[60561] = 25'b11101100_10001111_01111011_1;
      patterns[60562] = 25'b11101100_10010000_01111100_1;
      patterns[60563] = 25'b11101100_10010001_01111101_1;
      patterns[60564] = 25'b11101100_10010010_01111110_1;
      patterns[60565] = 25'b11101100_10010011_01111111_1;
      patterns[60566] = 25'b11101100_10010100_10000000_1;
      patterns[60567] = 25'b11101100_10010101_10000001_1;
      patterns[60568] = 25'b11101100_10010110_10000010_1;
      patterns[60569] = 25'b11101100_10010111_10000011_1;
      patterns[60570] = 25'b11101100_10011000_10000100_1;
      patterns[60571] = 25'b11101100_10011001_10000101_1;
      patterns[60572] = 25'b11101100_10011010_10000110_1;
      patterns[60573] = 25'b11101100_10011011_10000111_1;
      patterns[60574] = 25'b11101100_10011100_10001000_1;
      patterns[60575] = 25'b11101100_10011101_10001001_1;
      patterns[60576] = 25'b11101100_10011110_10001010_1;
      patterns[60577] = 25'b11101100_10011111_10001011_1;
      patterns[60578] = 25'b11101100_10100000_10001100_1;
      patterns[60579] = 25'b11101100_10100001_10001101_1;
      patterns[60580] = 25'b11101100_10100010_10001110_1;
      patterns[60581] = 25'b11101100_10100011_10001111_1;
      patterns[60582] = 25'b11101100_10100100_10010000_1;
      patterns[60583] = 25'b11101100_10100101_10010001_1;
      patterns[60584] = 25'b11101100_10100110_10010010_1;
      patterns[60585] = 25'b11101100_10100111_10010011_1;
      patterns[60586] = 25'b11101100_10101000_10010100_1;
      patterns[60587] = 25'b11101100_10101001_10010101_1;
      patterns[60588] = 25'b11101100_10101010_10010110_1;
      patterns[60589] = 25'b11101100_10101011_10010111_1;
      patterns[60590] = 25'b11101100_10101100_10011000_1;
      patterns[60591] = 25'b11101100_10101101_10011001_1;
      patterns[60592] = 25'b11101100_10101110_10011010_1;
      patterns[60593] = 25'b11101100_10101111_10011011_1;
      patterns[60594] = 25'b11101100_10110000_10011100_1;
      patterns[60595] = 25'b11101100_10110001_10011101_1;
      patterns[60596] = 25'b11101100_10110010_10011110_1;
      patterns[60597] = 25'b11101100_10110011_10011111_1;
      patterns[60598] = 25'b11101100_10110100_10100000_1;
      patterns[60599] = 25'b11101100_10110101_10100001_1;
      patterns[60600] = 25'b11101100_10110110_10100010_1;
      patterns[60601] = 25'b11101100_10110111_10100011_1;
      patterns[60602] = 25'b11101100_10111000_10100100_1;
      patterns[60603] = 25'b11101100_10111001_10100101_1;
      patterns[60604] = 25'b11101100_10111010_10100110_1;
      patterns[60605] = 25'b11101100_10111011_10100111_1;
      patterns[60606] = 25'b11101100_10111100_10101000_1;
      patterns[60607] = 25'b11101100_10111101_10101001_1;
      patterns[60608] = 25'b11101100_10111110_10101010_1;
      patterns[60609] = 25'b11101100_10111111_10101011_1;
      patterns[60610] = 25'b11101100_11000000_10101100_1;
      patterns[60611] = 25'b11101100_11000001_10101101_1;
      patterns[60612] = 25'b11101100_11000010_10101110_1;
      patterns[60613] = 25'b11101100_11000011_10101111_1;
      patterns[60614] = 25'b11101100_11000100_10110000_1;
      patterns[60615] = 25'b11101100_11000101_10110001_1;
      patterns[60616] = 25'b11101100_11000110_10110010_1;
      patterns[60617] = 25'b11101100_11000111_10110011_1;
      patterns[60618] = 25'b11101100_11001000_10110100_1;
      patterns[60619] = 25'b11101100_11001001_10110101_1;
      patterns[60620] = 25'b11101100_11001010_10110110_1;
      patterns[60621] = 25'b11101100_11001011_10110111_1;
      patterns[60622] = 25'b11101100_11001100_10111000_1;
      patterns[60623] = 25'b11101100_11001101_10111001_1;
      patterns[60624] = 25'b11101100_11001110_10111010_1;
      patterns[60625] = 25'b11101100_11001111_10111011_1;
      patterns[60626] = 25'b11101100_11010000_10111100_1;
      patterns[60627] = 25'b11101100_11010001_10111101_1;
      patterns[60628] = 25'b11101100_11010010_10111110_1;
      patterns[60629] = 25'b11101100_11010011_10111111_1;
      patterns[60630] = 25'b11101100_11010100_11000000_1;
      patterns[60631] = 25'b11101100_11010101_11000001_1;
      patterns[60632] = 25'b11101100_11010110_11000010_1;
      patterns[60633] = 25'b11101100_11010111_11000011_1;
      patterns[60634] = 25'b11101100_11011000_11000100_1;
      patterns[60635] = 25'b11101100_11011001_11000101_1;
      patterns[60636] = 25'b11101100_11011010_11000110_1;
      patterns[60637] = 25'b11101100_11011011_11000111_1;
      patterns[60638] = 25'b11101100_11011100_11001000_1;
      patterns[60639] = 25'b11101100_11011101_11001001_1;
      patterns[60640] = 25'b11101100_11011110_11001010_1;
      patterns[60641] = 25'b11101100_11011111_11001011_1;
      patterns[60642] = 25'b11101100_11100000_11001100_1;
      patterns[60643] = 25'b11101100_11100001_11001101_1;
      patterns[60644] = 25'b11101100_11100010_11001110_1;
      patterns[60645] = 25'b11101100_11100011_11001111_1;
      patterns[60646] = 25'b11101100_11100100_11010000_1;
      patterns[60647] = 25'b11101100_11100101_11010001_1;
      patterns[60648] = 25'b11101100_11100110_11010010_1;
      patterns[60649] = 25'b11101100_11100111_11010011_1;
      patterns[60650] = 25'b11101100_11101000_11010100_1;
      patterns[60651] = 25'b11101100_11101001_11010101_1;
      patterns[60652] = 25'b11101100_11101010_11010110_1;
      patterns[60653] = 25'b11101100_11101011_11010111_1;
      patterns[60654] = 25'b11101100_11101100_11011000_1;
      patterns[60655] = 25'b11101100_11101101_11011001_1;
      patterns[60656] = 25'b11101100_11101110_11011010_1;
      patterns[60657] = 25'b11101100_11101111_11011011_1;
      patterns[60658] = 25'b11101100_11110000_11011100_1;
      patterns[60659] = 25'b11101100_11110001_11011101_1;
      patterns[60660] = 25'b11101100_11110010_11011110_1;
      patterns[60661] = 25'b11101100_11110011_11011111_1;
      patterns[60662] = 25'b11101100_11110100_11100000_1;
      patterns[60663] = 25'b11101100_11110101_11100001_1;
      patterns[60664] = 25'b11101100_11110110_11100010_1;
      patterns[60665] = 25'b11101100_11110111_11100011_1;
      patterns[60666] = 25'b11101100_11111000_11100100_1;
      patterns[60667] = 25'b11101100_11111001_11100101_1;
      patterns[60668] = 25'b11101100_11111010_11100110_1;
      patterns[60669] = 25'b11101100_11111011_11100111_1;
      patterns[60670] = 25'b11101100_11111100_11101000_1;
      patterns[60671] = 25'b11101100_11111101_11101001_1;
      patterns[60672] = 25'b11101100_11111110_11101010_1;
      patterns[60673] = 25'b11101100_11111111_11101011_1;
      patterns[60674] = 25'b11101101_00000000_11101101_0;
      patterns[60675] = 25'b11101101_00000001_11101110_0;
      patterns[60676] = 25'b11101101_00000010_11101111_0;
      patterns[60677] = 25'b11101101_00000011_11110000_0;
      patterns[60678] = 25'b11101101_00000100_11110001_0;
      patterns[60679] = 25'b11101101_00000101_11110010_0;
      patterns[60680] = 25'b11101101_00000110_11110011_0;
      patterns[60681] = 25'b11101101_00000111_11110100_0;
      patterns[60682] = 25'b11101101_00001000_11110101_0;
      patterns[60683] = 25'b11101101_00001001_11110110_0;
      patterns[60684] = 25'b11101101_00001010_11110111_0;
      patterns[60685] = 25'b11101101_00001011_11111000_0;
      patterns[60686] = 25'b11101101_00001100_11111001_0;
      patterns[60687] = 25'b11101101_00001101_11111010_0;
      patterns[60688] = 25'b11101101_00001110_11111011_0;
      patterns[60689] = 25'b11101101_00001111_11111100_0;
      patterns[60690] = 25'b11101101_00010000_11111101_0;
      patterns[60691] = 25'b11101101_00010001_11111110_0;
      patterns[60692] = 25'b11101101_00010010_11111111_0;
      patterns[60693] = 25'b11101101_00010011_00000000_1;
      patterns[60694] = 25'b11101101_00010100_00000001_1;
      patterns[60695] = 25'b11101101_00010101_00000010_1;
      patterns[60696] = 25'b11101101_00010110_00000011_1;
      patterns[60697] = 25'b11101101_00010111_00000100_1;
      patterns[60698] = 25'b11101101_00011000_00000101_1;
      patterns[60699] = 25'b11101101_00011001_00000110_1;
      patterns[60700] = 25'b11101101_00011010_00000111_1;
      patterns[60701] = 25'b11101101_00011011_00001000_1;
      patterns[60702] = 25'b11101101_00011100_00001001_1;
      patterns[60703] = 25'b11101101_00011101_00001010_1;
      patterns[60704] = 25'b11101101_00011110_00001011_1;
      patterns[60705] = 25'b11101101_00011111_00001100_1;
      patterns[60706] = 25'b11101101_00100000_00001101_1;
      patterns[60707] = 25'b11101101_00100001_00001110_1;
      patterns[60708] = 25'b11101101_00100010_00001111_1;
      patterns[60709] = 25'b11101101_00100011_00010000_1;
      patterns[60710] = 25'b11101101_00100100_00010001_1;
      patterns[60711] = 25'b11101101_00100101_00010010_1;
      patterns[60712] = 25'b11101101_00100110_00010011_1;
      patterns[60713] = 25'b11101101_00100111_00010100_1;
      patterns[60714] = 25'b11101101_00101000_00010101_1;
      patterns[60715] = 25'b11101101_00101001_00010110_1;
      patterns[60716] = 25'b11101101_00101010_00010111_1;
      patterns[60717] = 25'b11101101_00101011_00011000_1;
      patterns[60718] = 25'b11101101_00101100_00011001_1;
      patterns[60719] = 25'b11101101_00101101_00011010_1;
      patterns[60720] = 25'b11101101_00101110_00011011_1;
      patterns[60721] = 25'b11101101_00101111_00011100_1;
      patterns[60722] = 25'b11101101_00110000_00011101_1;
      patterns[60723] = 25'b11101101_00110001_00011110_1;
      patterns[60724] = 25'b11101101_00110010_00011111_1;
      patterns[60725] = 25'b11101101_00110011_00100000_1;
      patterns[60726] = 25'b11101101_00110100_00100001_1;
      patterns[60727] = 25'b11101101_00110101_00100010_1;
      patterns[60728] = 25'b11101101_00110110_00100011_1;
      patterns[60729] = 25'b11101101_00110111_00100100_1;
      patterns[60730] = 25'b11101101_00111000_00100101_1;
      patterns[60731] = 25'b11101101_00111001_00100110_1;
      patterns[60732] = 25'b11101101_00111010_00100111_1;
      patterns[60733] = 25'b11101101_00111011_00101000_1;
      patterns[60734] = 25'b11101101_00111100_00101001_1;
      patterns[60735] = 25'b11101101_00111101_00101010_1;
      patterns[60736] = 25'b11101101_00111110_00101011_1;
      patterns[60737] = 25'b11101101_00111111_00101100_1;
      patterns[60738] = 25'b11101101_01000000_00101101_1;
      patterns[60739] = 25'b11101101_01000001_00101110_1;
      patterns[60740] = 25'b11101101_01000010_00101111_1;
      patterns[60741] = 25'b11101101_01000011_00110000_1;
      patterns[60742] = 25'b11101101_01000100_00110001_1;
      patterns[60743] = 25'b11101101_01000101_00110010_1;
      patterns[60744] = 25'b11101101_01000110_00110011_1;
      patterns[60745] = 25'b11101101_01000111_00110100_1;
      patterns[60746] = 25'b11101101_01001000_00110101_1;
      patterns[60747] = 25'b11101101_01001001_00110110_1;
      patterns[60748] = 25'b11101101_01001010_00110111_1;
      patterns[60749] = 25'b11101101_01001011_00111000_1;
      patterns[60750] = 25'b11101101_01001100_00111001_1;
      patterns[60751] = 25'b11101101_01001101_00111010_1;
      patterns[60752] = 25'b11101101_01001110_00111011_1;
      patterns[60753] = 25'b11101101_01001111_00111100_1;
      patterns[60754] = 25'b11101101_01010000_00111101_1;
      patterns[60755] = 25'b11101101_01010001_00111110_1;
      patterns[60756] = 25'b11101101_01010010_00111111_1;
      patterns[60757] = 25'b11101101_01010011_01000000_1;
      patterns[60758] = 25'b11101101_01010100_01000001_1;
      patterns[60759] = 25'b11101101_01010101_01000010_1;
      patterns[60760] = 25'b11101101_01010110_01000011_1;
      patterns[60761] = 25'b11101101_01010111_01000100_1;
      patterns[60762] = 25'b11101101_01011000_01000101_1;
      patterns[60763] = 25'b11101101_01011001_01000110_1;
      patterns[60764] = 25'b11101101_01011010_01000111_1;
      patterns[60765] = 25'b11101101_01011011_01001000_1;
      patterns[60766] = 25'b11101101_01011100_01001001_1;
      patterns[60767] = 25'b11101101_01011101_01001010_1;
      patterns[60768] = 25'b11101101_01011110_01001011_1;
      patterns[60769] = 25'b11101101_01011111_01001100_1;
      patterns[60770] = 25'b11101101_01100000_01001101_1;
      patterns[60771] = 25'b11101101_01100001_01001110_1;
      patterns[60772] = 25'b11101101_01100010_01001111_1;
      patterns[60773] = 25'b11101101_01100011_01010000_1;
      patterns[60774] = 25'b11101101_01100100_01010001_1;
      patterns[60775] = 25'b11101101_01100101_01010010_1;
      patterns[60776] = 25'b11101101_01100110_01010011_1;
      patterns[60777] = 25'b11101101_01100111_01010100_1;
      patterns[60778] = 25'b11101101_01101000_01010101_1;
      patterns[60779] = 25'b11101101_01101001_01010110_1;
      patterns[60780] = 25'b11101101_01101010_01010111_1;
      patterns[60781] = 25'b11101101_01101011_01011000_1;
      patterns[60782] = 25'b11101101_01101100_01011001_1;
      patterns[60783] = 25'b11101101_01101101_01011010_1;
      patterns[60784] = 25'b11101101_01101110_01011011_1;
      patterns[60785] = 25'b11101101_01101111_01011100_1;
      patterns[60786] = 25'b11101101_01110000_01011101_1;
      patterns[60787] = 25'b11101101_01110001_01011110_1;
      patterns[60788] = 25'b11101101_01110010_01011111_1;
      patterns[60789] = 25'b11101101_01110011_01100000_1;
      patterns[60790] = 25'b11101101_01110100_01100001_1;
      patterns[60791] = 25'b11101101_01110101_01100010_1;
      patterns[60792] = 25'b11101101_01110110_01100011_1;
      patterns[60793] = 25'b11101101_01110111_01100100_1;
      patterns[60794] = 25'b11101101_01111000_01100101_1;
      patterns[60795] = 25'b11101101_01111001_01100110_1;
      patterns[60796] = 25'b11101101_01111010_01100111_1;
      patterns[60797] = 25'b11101101_01111011_01101000_1;
      patterns[60798] = 25'b11101101_01111100_01101001_1;
      patterns[60799] = 25'b11101101_01111101_01101010_1;
      patterns[60800] = 25'b11101101_01111110_01101011_1;
      patterns[60801] = 25'b11101101_01111111_01101100_1;
      patterns[60802] = 25'b11101101_10000000_01101101_1;
      patterns[60803] = 25'b11101101_10000001_01101110_1;
      patterns[60804] = 25'b11101101_10000010_01101111_1;
      patterns[60805] = 25'b11101101_10000011_01110000_1;
      patterns[60806] = 25'b11101101_10000100_01110001_1;
      patterns[60807] = 25'b11101101_10000101_01110010_1;
      patterns[60808] = 25'b11101101_10000110_01110011_1;
      patterns[60809] = 25'b11101101_10000111_01110100_1;
      patterns[60810] = 25'b11101101_10001000_01110101_1;
      patterns[60811] = 25'b11101101_10001001_01110110_1;
      patterns[60812] = 25'b11101101_10001010_01110111_1;
      patterns[60813] = 25'b11101101_10001011_01111000_1;
      patterns[60814] = 25'b11101101_10001100_01111001_1;
      patterns[60815] = 25'b11101101_10001101_01111010_1;
      patterns[60816] = 25'b11101101_10001110_01111011_1;
      patterns[60817] = 25'b11101101_10001111_01111100_1;
      patterns[60818] = 25'b11101101_10010000_01111101_1;
      patterns[60819] = 25'b11101101_10010001_01111110_1;
      patterns[60820] = 25'b11101101_10010010_01111111_1;
      patterns[60821] = 25'b11101101_10010011_10000000_1;
      patterns[60822] = 25'b11101101_10010100_10000001_1;
      patterns[60823] = 25'b11101101_10010101_10000010_1;
      patterns[60824] = 25'b11101101_10010110_10000011_1;
      patterns[60825] = 25'b11101101_10010111_10000100_1;
      patterns[60826] = 25'b11101101_10011000_10000101_1;
      patterns[60827] = 25'b11101101_10011001_10000110_1;
      patterns[60828] = 25'b11101101_10011010_10000111_1;
      patterns[60829] = 25'b11101101_10011011_10001000_1;
      patterns[60830] = 25'b11101101_10011100_10001001_1;
      patterns[60831] = 25'b11101101_10011101_10001010_1;
      patterns[60832] = 25'b11101101_10011110_10001011_1;
      patterns[60833] = 25'b11101101_10011111_10001100_1;
      patterns[60834] = 25'b11101101_10100000_10001101_1;
      patterns[60835] = 25'b11101101_10100001_10001110_1;
      patterns[60836] = 25'b11101101_10100010_10001111_1;
      patterns[60837] = 25'b11101101_10100011_10010000_1;
      patterns[60838] = 25'b11101101_10100100_10010001_1;
      patterns[60839] = 25'b11101101_10100101_10010010_1;
      patterns[60840] = 25'b11101101_10100110_10010011_1;
      patterns[60841] = 25'b11101101_10100111_10010100_1;
      patterns[60842] = 25'b11101101_10101000_10010101_1;
      patterns[60843] = 25'b11101101_10101001_10010110_1;
      patterns[60844] = 25'b11101101_10101010_10010111_1;
      patterns[60845] = 25'b11101101_10101011_10011000_1;
      patterns[60846] = 25'b11101101_10101100_10011001_1;
      patterns[60847] = 25'b11101101_10101101_10011010_1;
      patterns[60848] = 25'b11101101_10101110_10011011_1;
      patterns[60849] = 25'b11101101_10101111_10011100_1;
      patterns[60850] = 25'b11101101_10110000_10011101_1;
      patterns[60851] = 25'b11101101_10110001_10011110_1;
      patterns[60852] = 25'b11101101_10110010_10011111_1;
      patterns[60853] = 25'b11101101_10110011_10100000_1;
      patterns[60854] = 25'b11101101_10110100_10100001_1;
      patterns[60855] = 25'b11101101_10110101_10100010_1;
      patterns[60856] = 25'b11101101_10110110_10100011_1;
      patterns[60857] = 25'b11101101_10110111_10100100_1;
      patterns[60858] = 25'b11101101_10111000_10100101_1;
      patterns[60859] = 25'b11101101_10111001_10100110_1;
      patterns[60860] = 25'b11101101_10111010_10100111_1;
      patterns[60861] = 25'b11101101_10111011_10101000_1;
      patterns[60862] = 25'b11101101_10111100_10101001_1;
      patterns[60863] = 25'b11101101_10111101_10101010_1;
      patterns[60864] = 25'b11101101_10111110_10101011_1;
      patterns[60865] = 25'b11101101_10111111_10101100_1;
      patterns[60866] = 25'b11101101_11000000_10101101_1;
      patterns[60867] = 25'b11101101_11000001_10101110_1;
      patterns[60868] = 25'b11101101_11000010_10101111_1;
      patterns[60869] = 25'b11101101_11000011_10110000_1;
      patterns[60870] = 25'b11101101_11000100_10110001_1;
      patterns[60871] = 25'b11101101_11000101_10110010_1;
      patterns[60872] = 25'b11101101_11000110_10110011_1;
      patterns[60873] = 25'b11101101_11000111_10110100_1;
      patterns[60874] = 25'b11101101_11001000_10110101_1;
      patterns[60875] = 25'b11101101_11001001_10110110_1;
      patterns[60876] = 25'b11101101_11001010_10110111_1;
      patterns[60877] = 25'b11101101_11001011_10111000_1;
      patterns[60878] = 25'b11101101_11001100_10111001_1;
      patterns[60879] = 25'b11101101_11001101_10111010_1;
      patterns[60880] = 25'b11101101_11001110_10111011_1;
      patterns[60881] = 25'b11101101_11001111_10111100_1;
      patterns[60882] = 25'b11101101_11010000_10111101_1;
      patterns[60883] = 25'b11101101_11010001_10111110_1;
      patterns[60884] = 25'b11101101_11010010_10111111_1;
      patterns[60885] = 25'b11101101_11010011_11000000_1;
      patterns[60886] = 25'b11101101_11010100_11000001_1;
      patterns[60887] = 25'b11101101_11010101_11000010_1;
      patterns[60888] = 25'b11101101_11010110_11000011_1;
      patterns[60889] = 25'b11101101_11010111_11000100_1;
      patterns[60890] = 25'b11101101_11011000_11000101_1;
      patterns[60891] = 25'b11101101_11011001_11000110_1;
      patterns[60892] = 25'b11101101_11011010_11000111_1;
      patterns[60893] = 25'b11101101_11011011_11001000_1;
      patterns[60894] = 25'b11101101_11011100_11001001_1;
      patterns[60895] = 25'b11101101_11011101_11001010_1;
      patterns[60896] = 25'b11101101_11011110_11001011_1;
      patterns[60897] = 25'b11101101_11011111_11001100_1;
      patterns[60898] = 25'b11101101_11100000_11001101_1;
      patterns[60899] = 25'b11101101_11100001_11001110_1;
      patterns[60900] = 25'b11101101_11100010_11001111_1;
      patterns[60901] = 25'b11101101_11100011_11010000_1;
      patterns[60902] = 25'b11101101_11100100_11010001_1;
      patterns[60903] = 25'b11101101_11100101_11010010_1;
      patterns[60904] = 25'b11101101_11100110_11010011_1;
      patterns[60905] = 25'b11101101_11100111_11010100_1;
      patterns[60906] = 25'b11101101_11101000_11010101_1;
      patterns[60907] = 25'b11101101_11101001_11010110_1;
      patterns[60908] = 25'b11101101_11101010_11010111_1;
      patterns[60909] = 25'b11101101_11101011_11011000_1;
      patterns[60910] = 25'b11101101_11101100_11011001_1;
      patterns[60911] = 25'b11101101_11101101_11011010_1;
      patterns[60912] = 25'b11101101_11101110_11011011_1;
      patterns[60913] = 25'b11101101_11101111_11011100_1;
      patterns[60914] = 25'b11101101_11110000_11011101_1;
      patterns[60915] = 25'b11101101_11110001_11011110_1;
      patterns[60916] = 25'b11101101_11110010_11011111_1;
      patterns[60917] = 25'b11101101_11110011_11100000_1;
      patterns[60918] = 25'b11101101_11110100_11100001_1;
      patterns[60919] = 25'b11101101_11110101_11100010_1;
      patterns[60920] = 25'b11101101_11110110_11100011_1;
      patterns[60921] = 25'b11101101_11110111_11100100_1;
      patterns[60922] = 25'b11101101_11111000_11100101_1;
      patterns[60923] = 25'b11101101_11111001_11100110_1;
      patterns[60924] = 25'b11101101_11111010_11100111_1;
      patterns[60925] = 25'b11101101_11111011_11101000_1;
      patterns[60926] = 25'b11101101_11111100_11101001_1;
      patterns[60927] = 25'b11101101_11111101_11101010_1;
      patterns[60928] = 25'b11101101_11111110_11101011_1;
      patterns[60929] = 25'b11101101_11111111_11101100_1;
      patterns[60930] = 25'b11101110_00000000_11101110_0;
      patterns[60931] = 25'b11101110_00000001_11101111_0;
      patterns[60932] = 25'b11101110_00000010_11110000_0;
      patterns[60933] = 25'b11101110_00000011_11110001_0;
      patterns[60934] = 25'b11101110_00000100_11110010_0;
      patterns[60935] = 25'b11101110_00000101_11110011_0;
      patterns[60936] = 25'b11101110_00000110_11110100_0;
      patterns[60937] = 25'b11101110_00000111_11110101_0;
      patterns[60938] = 25'b11101110_00001000_11110110_0;
      patterns[60939] = 25'b11101110_00001001_11110111_0;
      patterns[60940] = 25'b11101110_00001010_11111000_0;
      patterns[60941] = 25'b11101110_00001011_11111001_0;
      patterns[60942] = 25'b11101110_00001100_11111010_0;
      patterns[60943] = 25'b11101110_00001101_11111011_0;
      patterns[60944] = 25'b11101110_00001110_11111100_0;
      patterns[60945] = 25'b11101110_00001111_11111101_0;
      patterns[60946] = 25'b11101110_00010000_11111110_0;
      patterns[60947] = 25'b11101110_00010001_11111111_0;
      patterns[60948] = 25'b11101110_00010010_00000000_1;
      patterns[60949] = 25'b11101110_00010011_00000001_1;
      patterns[60950] = 25'b11101110_00010100_00000010_1;
      patterns[60951] = 25'b11101110_00010101_00000011_1;
      patterns[60952] = 25'b11101110_00010110_00000100_1;
      patterns[60953] = 25'b11101110_00010111_00000101_1;
      patterns[60954] = 25'b11101110_00011000_00000110_1;
      patterns[60955] = 25'b11101110_00011001_00000111_1;
      patterns[60956] = 25'b11101110_00011010_00001000_1;
      patterns[60957] = 25'b11101110_00011011_00001001_1;
      patterns[60958] = 25'b11101110_00011100_00001010_1;
      patterns[60959] = 25'b11101110_00011101_00001011_1;
      patterns[60960] = 25'b11101110_00011110_00001100_1;
      patterns[60961] = 25'b11101110_00011111_00001101_1;
      patterns[60962] = 25'b11101110_00100000_00001110_1;
      patterns[60963] = 25'b11101110_00100001_00001111_1;
      patterns[60964] = 25'b11101110_00100010_00010000_1;
      patterns[60965] = 25'b11101110_00100011_00010001_1;
      patterns[60966] = 25'b11101110_00100100_00010010_1;
      patterns[60967] = 25'b11101110_00100101_00010011_1;
      patterns[60968] = 25'b11101110_00100110_00010100_1;
      patterns[60969] = 25'b11101110_00100111_00010101_1;
      patterns[60970] = 25'b11101110_00101000_00010110_1;
      patterns[60971] = 25'b11101110_00101001_00010111_1;
      patterns[60972] = 25'b11101110_00101010_00011000_1;
      patterns[60973] = 25'b11101110_00101011_00011001_1;
      patterns[60974] = 25'b11101110_00101100_00011010_1;
      patterns[60975] = 25'b11101110_00101101_00011011_1;
      patterns[60976] = 25'b11101110_00101110_00011100_1;
      patterns[60977] = 25'b11101110_00101111_00011101_1;
      patterns[60978] = 25'b11101110_00110000_00011110_1;
      patterns[60979] = 25'b11101110_00110001_00011111_1;
      patterns[60980] = 25'b11101110_00110010_00100000_1;
      patterns[60981] = 25'b11101110_00110011_00100001_1;
      patterns[60982] = 25'b11101110_00110100_00100010_1;
      patterns[60983] = 25'b11101110_00110101_00100011_1;
      patterns[60984] = 25'b11101110_00110110_00100100_1;
      patterns[60985] = 25'b11101110_00110111_00100101_1;
      patterns[60986] = 25'b11101110_00111000_00100110_1;
      patterns[60987] = 25'b11101110_00111001_00100111_1;
      patterns[60988] = 25'b11101110_00111010_00101000_1;
      patterns[60989] = 25'b11101110_00111011_00101001_1;
      patterns[60990] = 25'b11101110_00111100_00101010_1;
      patterns[60991] = 25'b11101110_00111101_00101011_1;
      patterns[60992] = 25'b11101110_00111110_00101100_1;
      patterns[60993] = 25'b11101110_00111111_00101101_1;
      patterns[60994] = 25'b11101110_01000000_00101110_1;
      patterns[60995] = 25'b11101110_01000001_00101111_1;
      patterns[60996] = 25'b11101110_01000010_00110000_1;
      patterns[60997] = 25'b11101110_01000011_00110001_1;
      patterns[60998] = 25'b11101110_01000100_00110010_1;
      patterns[60999] = 25'b11101110_01000101_00110011_1;
      patterns[61000] = 25'b11101110_01000110_00110100_1;
      patterns[61001] = 25'b11101110_01000111_00110101_1;
      patterns[61002] = 25'b11101110_01001000_00110110_1;
      patterns[61003] = 25'b11101110_01001001_00110111_1;
      patterns[61004] = 25'b11101110_01001010_00111000_1;
      patterns[61005] = 25'b11101110_01001011_00111001_1;
      patterns[61006] = 25'b11101110_01001100_00111010_1;
      patterns[61007] = 25'b11101110_01001101_00111011_1;
      patterns[61008] = 25'b11101110_01001110_00111100_1;
      patterns[61009] = 25'b11101110_01001111_00111101_1;
      patterns[61010] = 25'b11101110_01010000_00111110_1;
      patterns[61011] = 25'b11101110_01010001_00111111_1;
      patterns[61012] = 25'b11101110_01010010_01000000_1;
      patterns[61013] = 25'b11101110_01010011_01000001_1;
      patterns[61014] = 25'b11101110_01010100_01000010_1;
      patterns[61015] = 25'b11101110_01010101_01000011_1;
      patterns[61016] = 25'b11101110_01010110_01000100_1;
      patterns[61017] = 25'b11101110_01010111_01000101_1;
      patterns[61018] = 25'b11101110_01011000_01000110_1;
      patterns[61019] = 25'b11101110_01011001_01000111_1;
      patterns[61020] = 25'b11101110_01011010_01001000_1;
      patterns[61021] = 25'b11101110_01011011_01001001_1;
      patterns[61022] = 25'b11101110_01011100_01001010_1;
      patterns[61023] = 25'b11101110_01011101_01001011_1;
      patterns[61024] = 25'b11101110_01011110_01001100_1;
      patterns[61025] = 25'b11101110_01011111_01001101_1;
      patterns[61026] = 25'b11101110_01100000_01001110_1;
      patterns[61027] = 25'b11101110_01100001_01001111_1;
      patterns[61028] = 25'b11101110_01100010_01010000_1;
      patterns[61029] = 25'b11101110_01100011_01010001_1;
      patterns[61030] = 25'b11101110_01100100_01010010_1;
      patterns[61031] = 25'b11101110_01100101_01010011_1;
      patterns[61032] = 25'b11101110_01100110_01010100_1;
      patterns[61033] = 25'b11101110_01100111_01010101_1;
      patterns[61034] = 25'b11101110_01101000_01010110_1;
      patterns[61035] = 25'b11101110_01101001_01010111_1;
      patterns[61036] = 25'b11101110_01101010_01011000_1;
      patterns[61037] = 25'b11101110_01101011_01011001_1;
      patterns[61038] = 25'b11101110_01101100_01011010_1;
      patterns[61039] = 25'b11101110_01101101_01011011_1;
      patterns[61040] = 25'b11101110_01101110_01011100_1;
      patterns[61041] = 25'b11101110_01101111_01011101_1;
      patterns[61042] = 25'b11101110_01110000_01011110_1;
      patterns[61043] = 25'b11101110_01110001_01011111_1;
      patterns[61044] = 25'b11101110_01110010_01100000_1;
      patterns[61045] = 25'b11101110_01110011_01100001_1;
      patterns[61046] = 25'b11101110_01110100_01100010_1;
      patterns[61047] = 25'b11101110_01110101_01100011_1;
      patterns[61048] = 25'b11101110_01110110_01100100_1;
      patterns[61049] = 25'b11101110_01110111_01100101_1;
      patterns[61050] = 25'b11101110_01111000_01100110_1;
      patterns[61051] = 25'b11101110_01111001_01100111_1;
      patterns[61052] = 25'b11101110_01111010_01101000_1;
      patterns[61053] = 25'b11101110_01111011_01101001_1;
      patterns[61054] = 25'b11101110_01111100_01101010_1;
      patterns[61055] = 25'b11101110_01111101_01101011_1;
      patterns[61056] = 25'b11101110_01111110_01101100_1;
      patterns[61057] = 25'b11101110_01111111_01101101_1;
      patterns[61058] = 25'b11101110_10000000_01101110_1;
      patterns[61059] = 25'b11101110_10000001_01101111_1;
      patterns[61060] = 25'b11101110_10000010_01110000_1;
      patterns[61061] = 25'b11101110_10000011_01110001_1;
      patterns[61062] = 25'b11101110_10000100_01110010_1;
      patterns[61063] = 25'b11101110_10000101_01110011_1;
      patterns[61064] = 25'b11101110_10000110_01110100_1;
      patterns[61065] = 25'b11101110_10000111_01110101_1;
      patterns[61066] = 25'b11101110_10001000_01110110_1;
      patterns[61067] = 25'b11101110_10001001_01110111_1;
      patterns[61068] = 25'b11101110_10001010_01111000_1;
      patterns[61069] = 25'b11101110_10001011_01111001_1;
      patterns[61070] = 25'b11101110_10001100_01111010_1;
      patterns[61071] = 25'b11101110_10001101_01111011_1;
      patterns[61072] = 25'b11101110_10001110_01111100_1;
      patterns[61073] = 25'b11101110_10001111_01111101_1;
      patterns[61074] = 25'b11101110_10010000_01111110_1;
      patterns[61075] = 25'b11101110_10010001_01111111_1;
      patterns[61076] = 25'b11101110_10010010_10000000_1;
      patterns[61077] = 25'b11101110_10010011_10000001_1;
      patterns[61078] = 25'b11101110_10010100_10000010_1;
      patterns[61079] = 25'b11101110_10010101_10000011_1;
      patterns[61080] = 25'b11101110_10010110_10000100_1;
      patterns[61081] = 25'b11101110_10010111_10000101_1;
      patterns[61082] = 25'b11101110_10011000_10000110_1;
      patterns[61083] = 25'b11101110_10011001_10000111_1;
      patterns[61084] = 25'b11101110_10011010_10001000_1;
      patterns[61085] = 25'b11101110_10011011_10001001_1;
      patterns[61086] = 25'b11101110_10011100_10001010_1;
      patterns[61087] = 25'b11101110_10011101_10001011_1;
      patterns[61088] = 25'b11101110_10011110_10001100_1;
      patterns[61089] = 25'b11101110_10011111_10001101_1;
      patterns[61090] = 25'b11101110_10100000_10001110_1;
      patterns[61091] = 25'b11101110_10100001_10001111_1;
      patterns[61092] = 25'b11101110_10100010_10010000_1;
      patterns[61093] = 25'b11101110_10100011_10010001_1;
      patterns[61094] = 25'b11101110_10100100_10010010_1;
      patterns[61095] = 25'b11101110_10100101_10010011_1;
      patterns[61096] = 25'b11101110_10100110_10010100_1;
      patterns[61097] = 25'b11101110_10100111_10010101_1;
      patterns[61098] = 25'b11101110_10101000_10010110_1;
      patterns[61099] = 25'b11101110_10101001_10010111_1;
      patterns[61100] = 25'b11101110_10101010_10011000_1;
      patterns[61101] = 25'b11101110_10101011_10011001_1;
      patterns[61102] = 25'b11101110_10101100_10011010_1;
      patterns[61103] = 25'b11101110_10101101_10011011_1;
      patterns[61104] = 25'b11101110_10101110_10011100_1;
      patterns[61105] = 25'b11101110_10101111_10011101_1;
      patterns[61106] = 25'b11101110_10110000_10011110_1;
      patterns[61107] = 25'b11101110_10110001_10011111_1;
      patterns[61108] = 25'b11101110_10110010_10100000_1;
      patterns[61109] = 25'b11101110_10110011_10100001_1;
      patterns[61110] = 25'b11101110_10110100_10100010_1;
      patterns[61111] = 25'b11101110_10110101_10100011_1;
      patterns[61112] = 25'b11101110_10110110_10100100_1;
      patterns[61113] = 25'b11101110_10110111_10100101_1;
      patterns[61114] = 25'b11101110_10111000_10100110_1;
      patterns[61115] = 25'b11101110_10111001_10100111_1;
      patterns[61116] = 25'b11101110_10111010_10101000_1;
      patterns[61117] = 25'b11101110_10111011_10101001_1;
      patterns[61118] = 25'b11101110_10111100_10101010_1;
      patterns[61119] = 25'b11101110_10111101_10101011_1;
      patterns[61120] = 25'b11101110_10111110_10101100_1;
      patterns[61121] = 25'b11101110_10111111_10101101_1;
      patterns[61122] = 25'b11101110_11000000_10101110_1;
      patterns[61123] = 25'b11101110_11000001_10101111_1;
      patterns[61124] = 25'b11101110_11000010_10110000_1;
      patterns[61125] = 25'b11101110_11000011_10110001_1;
      patterns[61126] = 25'b11101110_11000100_10110010_1;
      patterns[61127] = 25'b11101110_11000101_10110011_1;
      patterns[61128] = 25'b11101110_11000110_10110100_1;
      patterns[61129] = 25'b11101110_11000111_10110101_1;
      patterns[61130] = 25'b11101110_11001000_10110110_1;
      patterns[61131] = 25'b11101110_11001001_10110111_1;
      patterns[61132] = 25'b11101110_11001010_10111000_1;
      patterns[61133] = 25'b11101110_11001011_10111001_1;
      patterns[61134] = 25'b11101110_11001100_10111010_1;
      patterns[61135] = 25'b11101110_11001101_10111011_1;
      patterns[61136] = 25'b11101110_11001110_10111100_1;
      patterns[61137] = 25'b11101110_11001111_10111101_1;
      patterns[61138] = 25'b11101110_11010000_10111110_1;
      patterns[61139] = 25'b11101110_11010001_10111111_1;
      patterns[61140] = 25'b11101110_11010010_11000000_1;
      patterns[61141] = 25'b11101110_11010011_11000001_1;
      patterns[61142] = 25'b11101110_11010100_11000010_1;
      patterns[61143] = 25'b11101110_11010101_11000011_1;
      patterns[61144] = 25'b11101110_11010110_11000100_1;
      patterns[61145] = 25'b11101110_11010111_11000101_1;
      patterns[61146] = 25'b11101110_11011000_11000110_1;
      patterns[61147] = 25'b11101110_11011001_11000111_1;
      patterns[61148] = 25'b11101110_11011010_11001000_1;
      patterns[61149] = 25'b11101110_11011011_11001001_1;
      patterns[61150] = 25'b11101110_11011100_11001010_1;
      patterns[61151] = 25'b11101110_11011101_11001011_1;
      patterns[61152] = 25'b11101110_11011110_11001100_1;
      patterns[61153] = 25'b11101110_11011111_11001101_1;
      patterns[61154] = 25'b11101110_11100000_11001110_1;
      patterns[61155] = 25'b11101110_11100001_11001111_1;
      patterns[61156] = 25'b11101110_11100010_11010000_1;
      patterns[61157] = 25'b11101110_11100011_11010001_1;
      patterns[61158] = 25'b11101110_11100100_11010010_1;
      patterns[61159] = 25'b11101110_11100101_11010011_1;
      patterns[61160] = 25'b11101110_11100110_11010100_1;
      patterns[61161] = 25'b11101110_11100111_11010101_1;
      patterns[61162] = 25'b11101110_11101000_11010110_1;
      patterns[61163] = 25'b11101110_11101001_11010111_1;
      patterns[61164] = 25'b11101110_11101010_11011000_1;
      patterns[61165] = 25'b11101110_11101011_11011001_1;
      patterns[61166] = 25'b11101110_11101100_11011010_1;
      patterns[61167] = 25'b11101110_11101101_11011011_1;
      patterns[61168] = 25'b11101110_11101110_11011100_1;
      patterns[61169] = 25'b11101110_11101111_11011101_1;
      patterns[61170] = 25'b11101110_11110000_11011110_1;
      patterns[61171] = 25'b11101110_11110001_11011111_1;
      patterns[61172] = 25'b11101110_11110010_11100000_1;
      patterns[61173] = 25'b11101110_11110011_11100001_1;
      patterns[61174] = 25'b11101110_11110100_11100010_1;
      patterns[61175] = 25'b11101110_11110101_11100011_1;
      patterns[61176] = 25'b11101110_11110110_11100100_1;
      patterns[61177] = 25'b11101110_11110111_11100101_1;
      patterns[61178] = 25'b11101110_11111000_11100110_1;
      patterns[61179] = 25'b11101110_11111001_11100111_1;
      patterns[61180] = 25'b11101110_11111010_11101000_1;
      patterns[61181] = 25'b11101110_11111011_11101001_1;
      patterns[61182] = 25'b11101110_11111100_11101010_1;
      patterns[61183] = 25'b11101110_11111101_11101011_1;
      patterns[61184] = 25'b11101110_11111110_11101100_1;
      patterns[61185] = 25'b11101110_11111111_11101101_1;
      patterns[61186] = 25'b11101111_00000000_11101111_0;
      patterns[61187] = 25'b11101111_00000001_11110000_0;
      patterns[61188] = 25'b11101111_00000010_11110001_0;
      patterns[61189] = 25'b11101111_00000011_11110010_0;
      patterns[61190] = 25'b11101111_00000100_11110011_0;
      patterns[61191] = 25'b11101111_00000101_11110100_0;
      patterns[61192] = 25'b11101111_00000110_11110101_0;
      patterns[61193] = 25'b11101111_00000111_11110110_0;
      patterns[61194] = 25'b11101111_00001000_11110111_0;
      patterns[61195] = 25'b11101111_00001001_11111000_0;
      patterns[61196] = 25'b11101111_00001010_11111001_0;
      patterns[61197] = 25'b11101111_00001011_11111010_0;
      patterns[61198] = 25'b11101111_00001100_11111011_0;
      patterns[61199] = 25'b11101111_00001101_11111100_0;
      patterns[61200] = 25'b11101111_00001110_11111101_0;
      patterns[61201] = 25'b11101111_00001111_11111110_0;
      patterns[61202] = 25'b11101111_00010000_11111111_0;
      patterns[61203] = 25'b11101111_00010001_00000000_1;
      patterns[61204] = 25'b11101111_00010010_00000001_1;
      patterns[61205] = 25'b11101111_00010011_00000010_1;
      patterns[61206] = 25'b11101111_00010100_00000011_1;
      patterns[61207] = 25'b11101111_00010101_00000100_1;
      patterns[61208] = 25'b11101111_00010110_00000101_1;
      patterns[61209] = 25'b11101111_00010111_00000110_1;
      patterns[61210] = 25'b11101111_00011000_00000111_1;
      patterns[61211] = 25'b11101111_00011001_00001000_1;
      patterns[61212] = 25'b11101111_00011010_00001001_1;
      patterns[61213] = 25'b11101111_00011011_00001010_1;
      patterns[61214] = 25'b11101111_00011100_00001011_1;
      patterns[61215] = 25'b11101111_00011101_00001100_1;
      patterns[61216] = 25'b11101111_00011110_00001101_1;
      patterns[61217] = 25'b11101111_00011111_00001110_1;
      patterns[61218] = 25'b11101111_00100000_00001111_1;
      patterns[61219] = 25'b11101111_00100001_00010000_1;
      patterns[61220] = 25'b11101111_00100010_00010001_1;
      patterns[61221] = 25'b11101111_00100011_00010010_1;
      patterns[61222] = 25'b11101111_00100100_00010011_1;
      patterns[61223] = 25'b11101111_00100101_00010100_1;
      patterns[61224] = 25'b11101111_00100110_00010101_1;
      patterns[61225] = 25'b11101111_00100111_00010110_1;
      patterns[61226] = 25'b11101111_00101000_00010111_1;
      patterns[61227] = 25'b11101111_00101001_00011000_1;
      patterns[61228] = 25'b11101111_00101010_00011001_1;
      patterns[61229] = 25'b11101111_00101011_00011010_1;
      patterns[61230] = 25'b11101111_00101100_00011011_1;
      patterns[61231] = 25'b11101111_00101101_00011100_1;
      patterns[61232] = 25'b11101111_00101110_00011101_1;
      patterns[61233] = 25'b11101111_00101111_00011110_1;
      patterns[61234] = 25'b11101111_00110000_00011111_1;
      patterns[61235] = 25'b11101111_00110001_00100000_1;
      patterns[61236] = 25'b11101111_00110010_00100001_1;
      patterns[61237] = 25'b11101111_00110011_00100010_1;
      patterns[61238] = 25'b11101111_00110100_00100011_1;
      patterns[61239] = 25'b11101111_00110101_00100100_1;
      patterns[61240] = 25'b11101111_00110110_00100101_1;
      patterns[61241] = 25'b11101111_00110111_00100110_1;
      patterns[61242] = 25'b11101111_00111000_00100111_1;
      patterns[61243] = 25'b11101111_00111001_00101000_1;
      patterns[61244] = 25'b11101111_00111010_00101001_1;
      patterns[61245] = 25'b11101111_00111011_00101010_1;
      patterns[61246] = 25'b11101111_00111100_00101011_1;
      patterns[61247] = 25'b11101111_00111101_00101100_1;
      patterns[61248] = 25'b11101111_00111110_00101101_1;
      patterns[61249] = 25'b11101111_00111111_00101110_1;
      patterns[61250] = 25'b11101111_01000000_00101111_1;
      patterns[61251] = 25'b11101111_01000001_00110000_1;
      patterns[61252] = 25'b11101111_01000010_00110001_1;
      patterns[61253] = 25'b11101111_01000011_00110010_1;
      patterns[61254] = 25'b11101111_01000100_00110011_1;
      patterns[61255] = 25'b11101111_01000101_00110100_1;
      patterns[61256] = 25'b11101111_01000110_00110101_1;
      patterns[61257] = 25'b11101111_01000111_00110110_1;
      patterns[61258] = 25'b11101111_01001000_00110111_1;
      patterns[61259] = 25'b11101111_01001001_00111000_1;
      patterns[61260] = 25'b11101111_01001010_00111001_1;
      patterns[61261] = 25'b11101111_01001011_00111010_1;
      patterns[61262] = 25'b11101111_01001100_00111011_1;
      patterns[61263] = 25'b11101111_01001101_00111100_1;
      patterns[61264] = 25'b11101111_01001110_00111101_1;
      patterns[61265] = 25'b11101111_01001111_00111110_1;
      patterns[61266] = 25'b11101111_01010000_00111111_1;
      patterns[61267] = 25'b11101111_01010001_01000000_1;
      patterns[61268] = 25'b11101111_01010010_01000001_1;
      patterns[61269] = 25'b11101111_01010011_01000010_1;
      patterns[61270] = 25'b11101111_01010100_01000011_1;
      patterns[61271] = 25'b11101111_01010101_01000100_1;
      patterns[61272] = 25'b11101111_01010110_01000101_1;
      patterns[61273] = 25'b11101111_01010111_01000110_1;
      patterns[61274] = 25'b11101111_01011000_01000111_1;
      patterns[61275] = 25'b11101111_01011001_01001000_1;
      patterns[61276] = 25'b11101111_01011010_01001001_1;
      patterns[61277] = 25'b11101111_01011011_01001010_1;
      patterns[61278] = 25'b11101111_01011100_01001011_1;
      patterns[61279] = 25'b11101111_01011101_01001100_1;
      patterns[61280] = 25'b11101111_01011110_01001101_1;
      patterns[61281] = 25'b11101111_01011111_01001110_1;
      patterns[61282] = 25'b11101111_01100000_01001111_1;
      patterns[61283] = 25'b11101111_01100001_01010000_1;
      patterns[61284] = 25'b11101111_01100010_01010001_1;
      patterns[61285] = 25'b11101111_01100011_01010010_1;
      patterns[61286] = 25'b11101111_01100100_01010011_1;
      patterns[61287] = 25'b11101111_01100101_01010100_1;
      patterns[61288] = 25'b11101111_01100110_01010101_1;
      patterns[61289] = 25'b11101111_01100111_01010110_1;
      patterns[61290] = 25'b11101111_01101000_01010111_1;
      patterns[61291] = 25'b11101111_01101001_01011000_1;
      patterns[61292] = 25'b11101111_01101010_01011001_1;
      patterns[61293] = 25'b11101111_01101011_01011010_1;
      patterns[61294] = 25'b11101111_01101100_01011011_1;
      patterns[61295] = 25'b11101111_01101101_01011100_1;
      patterns[61296] = 25'b11101111_01101110_01011101_1;
      patterns[61297] = 25'b11101111_01101111_01011110_1;
      patterns[61298] = 25'b11101111_01110000_01011111_1;
      patterns[61299] = 25'b11101111_01110001_01100000_1;
      patterns[61300] = 25'b11101111_01110010_01100001_1;
      patterns[61301] = 25'b11101111_01110011_01100010_1;
      patterns[61302] = 25'b11101111_01110100_01100011_1;
      patterns[61303] = 25'b11101111_01110101_01100100_1;
      patterns[61304] = 25'b11101111_01110110_01100101_1;
      patterns[61305] = 25'b11101111_01110111_01100110_1;
      patterns[61306] = 25'b11101111_01111000_01100111_1;
      patterns[61307] = 25'b11101111_01111001_01101000_1;
      patterns[61308] = 25'b11101111_01111010_01101001_1;
      patterns[61309] = 25'b11101111_01111011_01101010_1;
      patterns[61310] = 25'b11101111_01111100_01101011_1;
      patterns[61311] = 25'b11101111_01111101_01101100_1;
      patterns[61312] = 25'b11101111_01111110_01101101_1;
      patterns[61313] = 25'b11101111_01111111_01101110_1;
      patterns[61314] = 25'b11101111_10000000_01101111_1;
      patterns[61315] = 25'b11101111_10000001_01110000_1;
      patterns[61316] = 25'b11101111_10000010_01110001_1;
      patterns[61317] = 25'b11101111_10000011_01110010_1;
      patterns[61318] = 25'b11101111_10000100_01110011_1;
      patterns[61319] = 25'b11101111_10000101_01110100_1;
      patterns[61320] = 25'b11101111_10000110_01110101_1;
      patterns[61321] = 25'b11101111_10000111_01110110_1;
      patterns[61322] = 25'b11101111_10001000_01110111_1;
      patterns[61323] = 25'b11101111_10001001_01111000_1;
      patterns[61324] = 25'b11101111_10001010_01111001_1;
      patterns[61325] = 25'b11101111_10001011_01111010_1;
      patterns[61326] = 25'b11101111_10001100_01111011_1;
      patterns[61327] = 25'b11101111_10001101_01111100_1;
      patterns[61328] = 25'b11101111_10001110_01111101_1;
      patterns[61329] = 25'b11101111_10001111_01111110_1;
      patterns[61330] = 25'b11101111_10010000_01111111_1;
      patterns[61331] = 25'b11101111_10010001_10000000_1;
      patterns[61332] = 25'b11101111_10010010_10000001_1;
      patterns[61333] = 25'b11101111_10010011_10000010_1;
      patterns[61334] = 25'b11101111_10010100_10000011_1;
      patterns[61335] = 25'b11101111_10010101_10000100_1;
      patterns[61336] = 25'b11101111_10010110_10000101_1;
      patterns[61337] = 25'b11101111_10010111_10000110_1;
      patterns[61338] = 25'b11101111_10011000_10000111_1;
      patterns[61339] = 25'b11101111_10011001_10001000_1;
      patterns[61340] = 25'b11101111_10011010_10001001_1;
      patterns[61341] = 25'b11101111_10011011_10001010_1;
      patterns[61342] = 25'b11101111_10011100_10001011_1;
      patterns[61343] = 25'b11101111_10011101_10001100_1;
      patterns[61344] = 25'b11101111_10011110_10001101_1;
      patterns[61345] = 25'b11101111_10011111_10001110_1;
      patterns[61346] = 25'b11101111_10100000_10001111_1;
      patterns[61347] = 25'b11101111_10100001_10010000_1;
      patterns[61348] = 25'b11101111_10100010_10010001_1;
      patterns[61349] = 25'b11101111_10100011_10010010_1;
      patterns[61350] = 25'b11101111_10100100_10010011_1;
      patterns[61351] = 25'b11101111_10100101_10010100_1;
      patterns[61352] = 25'b11101111_10100110_10010101_1;
      patterns[61353] = 25'b11101111_10100111_10010110_1;
      patterns[61354] = 25'b11101111_10101000_10010111_1;
      patterns[61355] = 25'b11101111_10101001_10011000_1;
      patterns[61356] = 25'b11101111_10101010_10011001_1;
      patterns[61357] = 25'b11101111_10101011_10011010_1;
      patterns[61358] = 25'b11101111_10101100_10011011_1;
      patterns[61359] = 25'b11101111_10101101_10011100_1;
      patterns[61360] = 25'b11101111_10101110_10011101_1;
      patterns[61361] = 25'b11101111_10101111_10011110_1;
      patterns[61362] = 25'b11101111_10110000_10011111_1;
      patterns[61363] = 25'b11101111_10110001_10100000_1;
      patterns[61364] = 25'b11101111_10110010_10100001_1;
      patterns[61365] = 25'b11101111_10110011_10100010_1;
      patterns[61366] = 25'b11101111_10110100_10100011_1;
      patterns[61367] = 25'b11101111_10110101_10100100_1;
      patterns[61368] = 25'b11101111_10110110_10100101_1;
      patterns[61369] = 25'b11101111_10110111_10100110_1;
      patterns[61370] = 25'b11101111_10111000_10100111_1;
      patterns[61371] = 25'b11101111_10111001_10101000_1;
      patterns[61372] = 25'b11101111_10111010_10101001_1;
      patterns[61373] = 25'b11101111_10111011_10101010_1;
      patterns[61374] = 25'b11101111_10111100_10101011_1;
      patterns[61375] = 25'b11101111_10111101_10101100_1;
      patterns[61376] = 25'b11101111_10111110_10101101_1;
      patterns[61377] = 25'b11101111_10111111_10101110_1;
      patterns[61378] = 25'b11101111_11000000_10101111_1;
      patterns[61379] = 25'b11101111_11000001_10110000_1;
      patterns[61380] = 25'b11101111_11000010_10110001_1;
      patterns[61381] = 25'b11101111_11000011_10110010_1;
      patterns[61382] = 25'b11101111_11000100_10110011_1;
      patterns[61383] = 25'b11101111_11000101_10110100_1;
      patterns[61384] = 25'b11101111_11000110_10110101_1;
      patterns[61385] = 25'b11101111_11000111_10110110_1;
      patterns[61386] = 25'b11101111_11001000_10110111_1;
      patterns[61387] = 25'b11101111_11001001_10111000_1;
      patterns[61388] = 25'b11101111_11001010_10111001_1;
      patterns[61389] = 25'b11101111_11001011_10111010_1;
      patterns[61390] = 25'b11101111_11001100_10111011_1;
      patterns[61391] = 25'b11101111_11001101_10111100_1;
      patterns[61392] = 25'b11101111_11001110_10111101_1;
      patterns[61393] = 25'b11101111_11001111_10111110_1;
      patterns[61394] = 25'b11101111_11010000_10111111_1;
      patterns[61395] = 25'b11101111_11010001_11000000_1;
      patterns[61396] = 25'b11101111_11010010_11000001_1;
      patterns[61397] = 25'b11101111_11010011_11000010_1;
      patterns[61398] = 25'b11101111_11010100_11000011_1;
      patterns[61399] = 25'b11101111_11010101_11000100_1;
      patterns[61400] = 25'b11101111_11010110_11000101_1;
      patterns[61401] = 25'b11101111_11010111_11000110_1;
      patterns[61402] = 25'b11101111_11011000_11000111_1;
      patterns[61403] = 25'b11101111_11011001_11001000_1;
      patterns[61404] = 25'b11101111_11011010_11001001_1;
      patterns[61405] = 25'b11101111_11011011_11001010_1;
      patterns[61406] = 25'b11101111_11011100_11001011_1;
      patterns[61407] = 25'b11101111_11011101_11001100_1;
      patterns[61408] = 25'b11101111_11011110_11001101_1;
      patterns[61409] = 25'b11101111_11011111_11001110_1;
      patterns[61410] = 25'b11101111_11100000_11001111_1;
      patterns[61411] = 25'b11101111_11100001_11010000_1;
      patterns[61412] = 25'b11101111_11100010_11010001_1;
      patterns[61413] = 25'b11101111_11100011_11010010_1;
      patterns[61414] = 25'b11101111_11100100_11010011_1;
      patterns[61415] = 25'b11101111_11100101_11010100_1;
      patterns[61416] = 25'b11101111_11100110_11010101_1;
      patterns[61417] = 25'b11101111_11100111_11010110_1;
      patterns[61418] = 25'b11101111_11101000_11010111_1;
      patterns[61419] = 25'b11101111_11101001_11011000_1;
      patterns[61420] = 25'b11101111_11101010_11011001_1;
      patterns[61421] = 25'b11101111_11101011_11011010_1;
      patterns[61422] = 25'b11101111_11101100_11011011_1;
      patterns[61423] = 25'b11101111_11101101_11011100_1;
      patterns[61424] = 25'b11101111_11101110_11011101_1;
      patterns[61425] = 25'b11101111_11101111_11011110_1;
      patterns[61426] = 25'b11101111_11110000_11011111_1;
      patterns[61427] = 25'b11101111_11110001_11100000_1;
      patterns[61428] = 25'b11101111_11110010_11100001_1;
      patterns[61429] = 25'b11101111_11110011_11100010_1;
      patterns[61430] = 25'b11101111_11110100_11100011_1;
      patterns[61431] = 25'b11101111_11110101_11100100_1;
      patterns[61432] = 25'b11101111_11110110_11100101_1;
      patterns[61433] = 25'b11101111_11110111_11100110_1;
      patterns[61434] = 25'b11101111_11111000_11100111_1;
      patterns[61435] = 25'b11101111_11111001_11101000_1;
      patterns[61436] = 25'b11101111_11111010_11101001_1;
      patterns[61437] = 25'b11101111_11111011_11101010_1;
      patterns[61438] = 25'b11101111_11111100_11101011_1;
      patterns[61439] = 25'b11101111_11111101_11101100_1;
      patterns[61440] = 25'b11101111_11111110_11101101_1;
      patterns[61441] = 25'b11101111_11111111_11101110_1;
      patterns[61442] = 25'b11110000_00000000_11110000_0;
      patterns[61443] = 25'b11110000_00000001_11110001_0;
      patterns[61444] = 25'b11110000_00000010_11110010_0;
      patterns[61445] = 25'b11110000_00000011_11110011_0;
      patterns[61446] = 25'b11110000_00000100_11110100_0;
      patterns[61447] = 25'b11110000_00000101_11110101_0;
      patterns[61448] = 25'b11110000_00000110_11110110_0;
      patterns[61449] = 25'b11110000_00000111_11110111_0;
      patterns[61450] = 25'b11110000_00001000_11111000_0;
      patterns[61451] = 25'b11110000_00001001_11111001_0;
      patterns[61452] = 25'b11110000_00001010_11111010_0;
      patterns[61453] = 25'b11110000_00001011_11111011_0;
      patterns[61454] = 25'b11110000_00001100_11111100_0;
      patterns[61455] = 25'b11110000_00001101_11111101_0;
      patterns[61456] = 25'b11110000_00001110_11111110_0;
      patterns[61457] = 25'b11110000_00001111_11111111_0;
      patterns[61458] = 25'b11110000_00010000_00000000_1;
      patterns[61459] = 25'b11110000_00010001_00000001_1;
      patterns[61460] = 25'b11110000_00010010_00000010_1;
      patterns[61461] = 25'b11110000_00010011_00000011_1;
      patterns[61462] = 25'b11110000_00010100_00000100_1;
      patterns[61463] = 25'b11110000_00010101_00000101_1;
      patterns[61464] = 25'b11110000_00010110_00000110_1;
      patterns[61465] = 25'b11110000_00010111_00000111_1;
      patterns[61466] = 25'b11110000_00011000_00001000_1;
      patterns[61467] = 25'b11110000_00011001_00001001_1;
      patterns[61468] = 25'b11110000_00011010_00001010_1;
      patterns[61469] = 25'b11110000_00011011_00001011_1;
      patterns[61470] = 25'b11110000_00011100_00001100_1;
      patterns[61471] = 25'b11110000_00011101_00001101_1;
      patterns[61472] = 25'b11110000_00011110_00001110_1;
      patterns[61473] = 25'b11110000_00011111_00001111_1;
      patterns[61474] = 25'b11110000_00100000_00010000_1;
      patterns[61475] = 25'b11110000_00100001_00010001_1;
      patterns[61476] = 25'b11110000_00100010_00010010_1;
      patterns[61477] = 25'b11110000_00100011_00010011_1;
      patterns[61478] = 25'b11110000_00100100_00010100_1;
      patterns[61479] = 25'b11110000_00100101_00010101_1;
      patterns[61480] = 25'b11110000_00100110_00010110_1;
      patterns[61481] = 25'b11110000_00100111_00010111_1;
      patterns[61482] = 25'b11110000_00101000_00011000_1;
      patterns[61483] = 25'b11110000_00101001_00011001_1;
      patterns[61484] = 25'b11110000_00101010_00011010_1;
      patterns[61485] = 25'b11110000_00101011_00011011_1;
      patterns[61486] = 25'b11110000_00101100_00011100_1;
      patterns[61487] = 25'b11110000_00101101_00011101_1;
      patterns[61488] = 25'b11110000_00101110_00011110_1;
      patterns[61489] = 25'b11110000_00101111_00011111_1;
      patterns[61490] = 25'b11110000_00110000_00100000_1;
      patterns[61491] = 25'b11110000_00110001_00100001_1;
      patterns[61492] = 25'b11110000_00110010_00100010_1;
      patterns[61493] = 25'b11110000_00110011_00100011_1;
      patterns[61494] = 25'b11110000_00110100_00100100_1;
      patterns[61495] = 25'b11110000_00110101_00100101_1;
      patterns[61496] = 25'b11110000_00110110_00100110_1;
      patterns[61497] = 25'b11110000_00110111_00100111_1;
      patterns[61498] = 25'b11110000_00111000_00101000_1;
      patterns[61499] = 25'b11110000_00111001_00101001_1;
      patterns[61500] = 25'b11110000_00111010_00101010_1;
      patterns[61501] = 25'b11110000_00111011_00101011_1;
      patterns[61502] = 25'b11110000_00111100_00101100_1;
      patterns[61503] = 25'b11110000_00111101_00101101_1;
      patterns[61504] = 25'b11110000_00111110_00101110_1;
      patterns[61505] = 25'b11110000_00111111_00101111_1;
      patterns[61506] = 25'b11110000_01000000_00110000_1;
      patterns[61507] = 25'b11110000_01000001_00110001_1;
      patterns[61508] = 25'b11110000_01000010_00110010_1;
      patterns[61509] = 25'b11110000_01000011_00110011_1;
      patterns[61510] = 25'b11110000_01000100_00110100_1;
      patterns[61511] = 25'b11110000_01000101_00110101_1;
      patterns[61512] = 25'b11110000_01000110_00110110_1;
      patterns[61513] = 25'b11110000_01000111_00110111_1;
      patterns[61514] = 25'b11110000_01001000_00111000_1;
      patterns[61515] = 25'b11110000_01001001_00111001_1;
      patterns[61516] = 25'b11110000_01001010_00111010_1;
      patterns[61517] = 25'b11110000_01001011_00111011_1;
      patterns[61518] = 25'b11110000_01001100_00111100_1;
      patterns[61519] = 25'b11110000_01001101_00111101_1;
      patterns[61520] = 25'b11110000_01001110_00111110_1;
      patterns[61521] = 25'b11110000_01001111_00111111_1;
      patterns[61522] = 25'b11110000_01010000_01000000_1;
      patterns[61523] = 25'b11110000_01010001_01000001_1;
      patterns[61524] = 25'b11110000_01010010_01000010_1;
      patterns[61525] = 25'b11110000_01010011_01000011_1;
      patterns[61526] = 25'b11110000_01010100_01000100_1;
      patterns[61527] = 25'b11110000_01010101_01000101_1;
      patterns[61528] = 25'b11110000_01010110_01000110_1;
      patterns[61529] = 25'b11110000_01010111_01000111_1;
      patterns[61530] = 25'b11110000_01011000_01001000_1;
      patterns[61531] = 25'b11110000_01011001_01001001_1;
      patterns[61532] = 25'b11110000_01011010_01001010_1;
      patterns[61533] = 25'b11110000_01011011_01001011_1;
      patterns[61534] = 25'b11110000_01011100_01001100_1;
      patterns[61535] = 25'b11110000_01011101_01001101_1;
      patterns[61536] = 25'b11110000_01011110_01001110_1;
      patterns[61537] = 25'b11110000_01011111_01001111_1;
      patterns[61538] = 25'b11110000_01100000_01010000_1;
      patterns[61539] = 25'b11110000_01100001_01010001_1;
      patterns[61540] = 25'b11110000_01100010_01010010_1;
      patterns[61541] = 25'b11110000_01100011_01010011_1;
      patterns[61542] = 25'b11110000_01100100_01010100_1;
      patterns[61543] = 25'b11110000_01100101_01010101_1;
      patterns[61544] = 25'b11110000_01100110_01010110_1;
      patterns[61545] = 25'b11110000_01100111_01010111_1;
      patterns[61546] = 25'b11110000_01101000_01011000_1;
      patterns[61547] = 25'b11110000_01101001_01011001_1;
      patterns[61548] = 25'b11110000_01101010_01011010_1;
      patterns[61549] = 25'b11110000_01101011_01011011_1;
      patterns[61550] = 25'b11110000_01101100_01011100_1;
      patterns[61551] = 25'b11110000_01101101_01011101_1;
      patterns[61552] = 25'b11110000_01101110_01011110_1;
      patterns[61553] = 25'b11110000_01101111_01011111_1;
      patterns[61554] = 25'b11110000_01110000_01100000_1;
      patterns[61555] = 25'b11110000_01110001_01100001_1;
      patterns[61556] = 25'b11110000_01110010_01100010_1;
      patterns[61557] = 25'b11110000_01110011_01100011_1;
      patterns[61558] = 25'b11110000_01110100_01100100_1;
      patterns[61559] = 25'b11110000_01110101_01100101_1;
      patterns[61560] = 25'b11110000_01110110_01100110_1;
      patterns[61561] = 25'b11110000_01110111_01100111_1;
      patterns[61562] = 25'b11110000_01111000_01101000_1;
      patterns[61563] = 25'b11110000_01111001_01101001_1;
      patterns[61564] = 25'b11110000_01111010_01101010_1;
      patterns[61565] = 25'b11110000_01111011_01101011_1;
      patterns[61566] = 25'b11110000_01111100_01101100_1;
      patterns[61567] = 25'b11110000_01111101_01101101_1;
      patterns[61568] = 25'b11110000_01111110_01101110_1;
      patterns[61569] = 25'b11110000_01111111_01101111_1;
      patterns[61570] = 25'b11110000_10000000_01110000_1;
      patterns[61571] = 25'b11110000_10000001_01110001_1;
      patterns[61572] = 25'b11110000_10000010_01110010_1;
      patterns[61573] = 25'b11110000_10000011_01110011_1;
      patterns[61574] = 25'b11110000_10000100_01110100_1;
      patterns[61575] = 25'b11110000_10000101_01110101_1;
      patterns[61576] = 25'b11110000_10000110_01110110_1;
      patterns[61577] = 25'b11110000_10000111_01110111_1;
      patterns[61578] = 25'b11110000_10001000_01111000_1;
      patterns[61579] = 25'b11110000_10001001_01111001_1;
      patterns[61580] = 25'b11110000_10001010_01111010_1;
      patterns[61581] = 25'b11110000_10001011_01111011_1;
      patterns[61582] = 25'b11110000_10001100_01111100_1;
      patterns[61583] = 25'b11110000_10001101_01111101_1;
      patterns[61584] = 25'b11110000_10001110_01111110_1;
      patterns[61585] = 25'b11110000_10001111_01111111_1;
      patterns[61586] = 25'b11110000_10010000_10000000_1;
      patterns[61587] = 25'b11110000_10010001_10000001_1;
      patterns[61588] = 25'b11110000_10010010_10000010_1;
      patterns[61589] = 25'b11110000_10010011_10000011_1;
      patterns[61590] = 25'b11110000_10010100_10000100_1;
      patterns[61591] = 25'b11110000_10010101_10000101_1;
      patterns[61592] = 25'b11110000_10010110_10000110_1;
      patterns[61593] = 25'b11110000_10010111_10000111_1;
      patterns[61594] = 25'b11110000_10011000_10001000_1;
      patterns[61595] = 25'b11110000_10011001_10001001_1;
      patterns[61596] = 25'b11110000_10011010_10001010_1;
      patterns[61597] = 25'b11110000_10011011_10001011_1;
      patterns[61598] = 25'b11110000_10011100_10001100_1;
      patterns[61599] = 25'b11110000_10011101_10001101_1;
      patterns[61600] = 25'b11110000_10011110_10001110_1;
      patterns[61601] = 25'b11110000_10011111_10001111_1;
      patterns[61602] = 25'b11110000_10100000_10010000_1;
      patterns[61603] = 25'b11110000_10100001_10010001_1;
      patterns[61604] = 25'b11110000_10100010_10010010_1;
      patterns[61605] = 25'b11110000_10100011_10010011_1;
      patterns[61606] = 25'b11110000_10100100_10010100_1;
      patterns[61607] = 25'b11110000_10100101_10010101_1;
      patterns[61608] = 25'b11110000_10100110_10010110_1;
      patterns[61609] = 25'b11110000_10100111_10010111_1;
      patterns[61610] = 25'b11110000_10101000_10011000_1;
      patterns[61611] = 25'b11110000_10101001_10011001_1;
      patterns[61612] = 25'b11110000_10101010_10011010_1;
      patterns[61613] = 25'b11110000_10101011_10011011_1;
      patterns[61614] = 25'b11110000_10101100_10011100_1;
      patterns[61615] = 25'b11110000_10101101_10011101_1;
      patterns[61616] = 25'b11110000_10101110_10011110_1;
      patterns[61617] = 25'b11110000_10101111_10011111_1;
      patterns[61618] = 25'b11110000_10110000_10100000_1;
      patterns[61619] = 25'b11110000_10110001_10100001_1;
      patterns[61620] = 25'b11110000_10110010_10100010_1;
      patterns[61621] = 25'b11110000_10110011_10100011_1;
      patterns[61622] = 25'b11110000_10110100_10100100_1;
      patterns[61623] = 25'b11110000_10110101_10100101_1;
      patterns[61624] = 25'b11110000_10110110_10100110_1;
      patterns[61625] = 25'b11110000_10110111_10100111_1;
      patterns[61626] = 25'b11110000_10111000_10101000_1;
      patterns[61627] = 25'b11110000_10111001_10101001_1;
      patterns[61628] = 25'b11110000_10111010_10101010_1;
      patterns[61629] = 25'b11110000_10111011_10101011_1;
      patterns[61630] = 25'b11110000_10111100_10101100_1;
      patterns[61631] = 25'b11110000_10111101_10101101_1;
      patterns[61632] = 25'b11110000_10111110_10101110_1;
      patterns[61633] = 25'b11110000_10111111_10101111_1;
      patterns[61634] = 25'b11110000_11000000_10110000_1;
      patterns[61635] = 25'b11110000_11000001_10110001_1;
      patterns[61636] = 25'b11110000_11000010_10110010_1;
      patterns[61637] = 25'b11110000_11000011_10110011_1;
      patterns[61638] = 25'b11110000_11000100_10110100_1;
      patterns[61639] = 25'b11110000_11000101_10110101_1;
      patterns[61640] = 25'b11110000_11000110_10110110_1;
      patterns[61641] = 25'b11110000_11000111_10110111_1;
      patterns[61642] = 25'b11110000_11001000_10111000_1;
      patterns[61643] = 25'b11110000_11001001_10111001_1;
      patterns[61644] = 25'b11110000_11001010_10111010_1;
      patterns[61645] = 25'b11110000_11001011_10111011_1;
      patterns[61646] = 25'b11110000_11001100_10111100_1;
      patterns[61647] = 25'b11110000_11001101_10111101_1;
      patterns[61648] = 25'b11110000_11001110_10111110_1;
      patterns[61649] = 25'b11110000_11001111_10111111_1;
      patterns[61650] = 25'b11110000_11010000_11000000_1;
      patterns[61651] = 25'b11110000_11010001_11000001_1;
      patterns[61652] = 25'b11110000_11010010_11000010_1;
      patterns[61653] = 25'b11110000_11010011_11000011_1;
      patterns[61654] = 25'b11110000_11010100_11000100_1;
      patterns[61655] = 25'b11110000_11010101_11000101_1;
      patterns[61656] = 25'b11110000_11010110_11000110_1;
      patterns[61657] = 25'b11110000_11010111_11000111_1;
      patterns[61658] = 25'b11110000_11011000_11001000_1;
      patterns[61659] = 25'b11110000_11011001_11001001_1;
      patterns[61660] = 25'b11110000_11011010_11001010_1;
      patterns[61661] = 25'b11110000_11011011_11001011_1;
      patterns[61662] = 25'b11110000_11011100_11001100_1;
      patterns[61663] = 25'b11110000_11011101_11001101_1;
      patterns[61664] = 25'b11110000_11011110_11001110_1;
      patterns[61665] = 25'b11110000_11011111_11001111_1;
      patterns[61666] = 25'b11110000_11100000_11010000_1;
      patterns[61667] = 25'b11110000_11100001_11010001_1;
      patterns[61668] = 25'b11110000_11100010_11010010_1;
      patterns[61669] = 25'b11110000_11100011_11010011_1;
      patterns[61670] = 25'b11110000_11100100_11010100_1;
      patterns[61671] = 25'b11110000_11100101_11010101_1;
      patterns[61672] = 25'b11110000_11100110_11010110_1;
      patterns[61673] = 25'b11110000_11100111_11010111_1;
      patterns[61674] = 25'b11110000_11101000_11011000_1;
      patterns[61675] = 25'b11110000_11101001_11011001_1;
      patterns[61676] = 25'b11110000_11101010_11011010_1;
      patterns[61677] = 25'b11110000_11101011_11011011_1;
      patterns[61678] = 25'b11110000_11101100_11011100_1;
      patterns[61679] = 25'b11110000_11101101_11011101_1;
      patterns[61680] = 25'b11110000_11101110_11011110_1;
      patterns[61681] = 25'b11110000_11101111_11011111_1;
      patterns[61682] = 25'b11110000_11110000_11100000_1;
      patterns[61683] = 25'b11110000_11110001_11100001_1;
      patterns[61684] = 25'b11110000_11110010_11100010_1;
      patterns[61685] = 25'b11110000_11110011_11100011_1;
      patterns[61686] = 25'b11110000_11110100_11100100_1;
      patterns[61687] = 25'b11110000_11110101_11100101_1;
      patterns[61688] = 25'b11110000_11110110_11100110_1;
      patterns[61689] = 25'b11110000_11110111_11100111_1;
      patterns[61690] = 25'b11110000_11111000_11101000_1;
      patterns[61691] = 25'b11110000_11111001_11101001_1;
      patterns[61692] = 25'b11110000_11111010_11101010_1;
      patterns[61693] = 25'b11110000_11111011_11101011_1;
      patterns[61694] = 25'b11110000_11111100_11101100_1;
      patterns[61695] = 25'b11110000_11111101_11101101_1;
      patterns[61696] = 25'b11110000_11111110_11101110_1;
      patterns[61697] = 25'b11110000_11111111_11101111_1;
      patterns[61698] = 25'b11110001_00000000_11110001_0;
      patterns[61699] = 25'b11110001_00000001_11110010_0;
      patterns[61700] = 25'b11110001_00000010_11110011_0;
      patterns[61701] = 25'b11110001_00000011_11110100_0;
      patterns[61702] = 25'b11110001_00000100_11110101_0;
      patterns[61703] = 25'b11110001_00000101_11110110_0;
      patterns[61704] = 25'b11110001_00000110_11110111_0;
      patterns[61705] = 25'b11110001_00000111_11111000_0;
      patterns[61706] = 25'b11110001_00001000_11111001_0;
      patterns[61707] = 25'b11110001_00001001_11111010_0;
      patterns[61708] = 25'b11110001_00001010_11111011_0;
      patterns[61709] = 25'b11110001_00001011_11111100_0;
      patterns[61710] = 25'b11110001_00001100_11111101_0;
      patterns[61711] = 25'b11110001_00001101_11111110_0;
      patterns[61712] = 25'b11110001_00001110_11111111_0;
      patterns[61713] = 25'b11110001_00001111_00000000_1;
      patterns[61714] = 25'b11110001_00010000_00000001_1;
      patterns[61715] = 25'b11110001_00010001_00000010_1;
      patterns[61716] = 25'b11110001_00010010_00000011_1;
      patterns[61717] = 25'b11110001_00010011_00000100_1;
      patterns[61718] = 25'b11110001_00010100_00000101_1;
      patterns[61719] = 25'b11110001_00010101_00000110_1;
      patterns[61720] = 25'b11110001_00010110_00000111_1;
      patterns[61721] = 25'b11110001_00010111_00001000_1;
      patterns[61722] = 25'b11110001_00011000_00001001_1;
      patterns[61723] = 25'b11110001_00011001_00001010_1;
      patterns[61724] = 25'b11110001_00011010_00001011_1;
      patterns[61725] = 25'b11110001_00011011_00001100_1;
      patterns[61726] = 25'b11110001_00011100_00001101_1;
      patterns[61727] = 25'b11110001_00011101_00001110_1;
      patterns[61728] = 25'b11110001_00011110_00001111_1;
      patterns[61729] = 25'b11110001_00011111_00010000_1;
      patterns[61730] = 25'b11110001_00100000_00010001_1;
      patterns[61731] = 25'b11110001_00100001_00010010_1;
      patterns[61732] = 25'b11110001_00100010_00010011_1;
      patterns[61733] = 25'b11110001_00100011_00010100_1;
      patterns[61734] = 25'b11110001_00100100_00010101_1;
      patterns[61735] = 25'b11110001_00100101_00010110_1;
      patterns[61736] = 25'b11110001_00100110_00010111_1;
      patterns[61737] = 25'b11110001_00100111_00011000_1;
      patterns[61738] = 25'b11110001_00101000_00011001_1;
      patterns[61739] = 25'b11110001_00101001_00011010_1;
      patterns[61740] = 25'b11110001_00101010_00011011_1;
      patterns[61741] = 25'b11110001_00101011_00011100_1;
      patterns[61742] = 25'b11110001_00101100_00011101_1;
      patterns[61743] = 25'b11110001_00101101_00011110_1;
      patterns[61744] = 25'b11110001_00101110_00011111_1;
      patterns[61745] = 25'b11110001_00101111_00100000_1;
      patterns[61746] = 25'b11110001_00110000_00100001_1;
      patterns[61747] = 25'b11110001_00110001_00100010_1;
      patterns[61748] = 25'b11110001_00110010_00100011_1;
      patterns[61749] = 25'b11110001_00110011_00100100_1;
      patterns[61750] = 25'b11110001_00110100_00100101_1;
      patterns[61751] = 25'b11110001_00110101_00100110_1;
      patterns[61752] = 25'b11110001_00110110_00100111_1;
      patterns[61753] = 25'b11110001_00110111_00101000_1;
      patterns[61754] = 25'b11110001_00111000_00101001_1;
      patterns[61755] = 25'b11110001_00111001_00101010_1;
      patterns[61756] = 25'b11110001_00111010_00101011_1;
      patterns[61757] = 25'b11110001_00111011_00101100_1;
      patterns[61758] = 25'b11110001_00111100_00101101_1;
      patterns[61759] = 25'b11110001_00111101_00101110_1;
      patterns[61760] = 25'b11110001_00111110_00101111_1;
      patterns[61761] = 25'b11110001_00111111_00110000_1;
      patterns[61762] = 25'b11110001_01000000_00110001_1;
      patterns[61763] = 25'b11110001_01000001_00110010_1;
      patterns[61764] = 25'b11110001_01000010_00110011_1;
      patterns[61765] = 25'b11110001_01000011_00110100_1;
      patterns[61766] = 25'b11110001_01000100_00110101_1;
      patterns[61767] = 25'b11110001_01000101_00110110_1;
      patterns[61768] = 25'b11110001_01000110_00110111_1;
      patterns[61769] = 25'b11110001_01000111_00111000_1;
      patterns[61770] = 25'b11110001_01001000_00111001_1;
      patterns[61771] = 25'b11110001_01001001_00111010_1;
      patterns[61772] = 25'b11110001_01001010_00111011_1;
      patterns[61773] = 25'b11110001_01001011_00111100_1;
      patterns[61774] = 25'b11110001_01001100_00111101_1;
      patterns[61775] = 25'b11110001_01001101_00111110_1;
      patterns[61776] = 25'b11110001_01001110_00111111_1;
      patterns[61777] = 25'b11110001_01001111_01000000_1;
      patterns[61778] = 25'b11110001_01010000_01000001_1;
      patterns[61779] = 25'b11110001_01010001_01000010_1;
      patterns[61780] = 25'b11110001_01010010_01000011_1;
      patterns[61781] = 25'b11110001_01010011_01000100_1;
      patterns[61782] = 25'b11110001_01010100_01000101_1;
      patterns[61783] = 25'b11110001_01010101_01000110_1;
      patterns[61784] = 25'b11110001_01010110_01000111_1;
      patterns[61785] = 25'b11110001_01010111_01001000_1;
      patterns[61786] = 25'b11110001_01011000_01001001_1;
      patterns[61787] = 25'b11110001_01011001_01001010_1;
      patterns[61788] = 25'b11110001_01011010_01001011_1;
      patterns[61789] = 25'b11110001_01011011_01001100_1;
      patterns[61790] = 25'b11110001_01011100_01001101_1;
      patterns[61791] = 25'b11110001_01011101_01001110_1;
      patterns[61792] = 25'b11110001_01011110_01001111_1;
      patterns[61793] = 25'b11110001_01011111_01010000_1;
      patterns[61794] = 25'b11110001_01100000_01010001_1;
      patterns[61795] = 25'b11110001_01100001_01010010_1;
      patterns[61796] = 25'b11110001_01100010_01010011_1;
      patterns[61797] = 25'b11110001_01100011_01010100_1;
      patterns[61798] = 25'b11110001_01100100_01010101_1;
      patterns[61799] = 25'b11110001_01100101_01010110_1;
      patterns[61800] = 25'b11110001_01100110_01010111_1;
      patterns[61801] = 25'b11110001_01100111_01011000_1;
      patterns[61802] = 25'b11110001_01101000_01011001_1;
      patterns[61803] = 25'b11110001_01101001_01011010_1;
      patterns[61804] = 25'b11110001_01101010_01011011_1;
      patterns[61805] = 25'b11110001_01101011_01011100_1;
      patterns[61806] = 25'b11110001_01101100_01011101_1;
      patterns[61807] = 25'b11110001_01101101_01011110_1;
      patterns[61808] = 25'b11110001_01101110_01011111_1;
      patterns[61809] = 25'b11110001_01101111_01100000_1;
      patterns[61810] = 25'b11110001_01110000_01100001_1;
      patterns[61811] = 25'b11110001_01110001_01100010_1;
      patterns[61812] = 25'b11110001_01110010_01100011_1;
      patterns[61813] = 25'b11110001_01110011_01100100_1;
      patterns[61814] = 25'b11110001_01110100_01100101_1;
      patterns[61815] = 25'b11110001_01110101_01100110_1;
      patterns[61816] = 25'b11110001_01110110_01100111_1;
      patterns[61817] = 25'b11110001_01110111_01101000_1;
      patterns[61818] = 25'b11110001_01111000_01101001_1;
      patterns[61819] = 25'b11110001_01111001_01101010_1;
      patterns[61820] = 25'b11110001_01111010_01101011_1;
      patterns[61821] = 25'b11110001_01111011_01101100_1;
      patterns[61822] = 25'b11110001_01111100_01101101_1;
      patterns[61823] = 25'b11110001_01111101_01101110_1;
      patterns[61824] = 25'b11110001_01111110_01101111_1;
      patterns[61825] = 25'b11110001_01111111_01110000_1;
      patterns[61826] = 25'b11110001_10000000_01110001_1;
      patterns[61827] = 25'b11110001_10000001_01110010_1;
      patterns[61828] = 25'b11110001_10000010_01110011_1;
      patterns[61829] = 25'b11110001_10000011_01110100_1;
      patterns[61830] = 25'b11110001_10000100_01110101_1;
      patterns[61831] = 25'b11110001_10000101_01110110_1;
      patterns[61832] = 25'b11110001_10000110_01110111_1;
      patterns[61833] = 25'b11110001_10000111_01111000_1;
      patterns[61834] = 25'b11110001_10001000_01111001_1;
      patterns[61835] = 25'b11110001_10001001_01111010_1;
      patterns[61836] = 25'b11110001_10001010_01111011_1;
      patterns[61837] = 25'b11110001_10001011_01111100_1;
      patterns[61838] = 25'b11110001_10001100_01111101_1;
      patterns[61839] = 25'b11110001_10001101_01111110_1;
      patterns[61840] = 25'b11110001_10001110_01111111_1;
      patterns[61841] = 25'b11110001_10001111_10000000_1;
      patterns[61842] = 25'b11110001_10010000_10000001_1;
      patterns[61843] = 25'b11110001_10010001_10000010_1;
      patterns[61844] = 25'b11110001_10010010_10000011_1;
      patterns[61845] = 25'b11110001_10010011_10000100_1;
      patterns[61846] = 25'b11110001_10010100_10000101_1;
      patterns[61847] = 25'b11110001_10010101_10000110_1;
      patterns[61848] = 25'b11110001_10010110_10000111_1;
      patterns[61849] = 25'b11110001_10010111_10001000_1;
      patterns[61850] = 25'b11110001_10011000_10001001_1;
      patterns[61851] = 25'b11110001_10011001_10001010_1;
      patterns[61852] = 25'b11110001_10011010_10001011_1;
      patterns[61853] = 25'b11110001_10011011_10001100_1;
      patterns[61854] = 25'b11110001_10011100_10001101_1;
      patterns[61855] = 25'b11110001_10011101_10001110_1;
      patterns[61856] = 25'b11110001_10011110_10001111_1;
      patterns[61857] = 25'b11110001_10011111_10010000_1;
      patterns[61858] = 25'b11110001_10100000_10010001_1;
      patterns[61859] = 25'b11110001_10100001_10010010_1;
      patterns[61860] = 25'b11110001_10100010_10010011_1;
      patterns[61861] = 25'b11110001_10100011_10010100_1;
      patterns[61862] = 25'b11110001_10100100_10010101_1;
      patterns[61863] = 25'b11110001_10100101_10010110_1;
      patterns[61864] = 25'b11110001_10100110_10010111_1;
      patterns[61865] = 25'b11110001_10100111_10011000_1;
      patterns[61866] = 25'b11110001_10101000_10011001_1;
      patterns[61867] = 25'b11110001_10101001_10011010_1;
      patterns[61868] = 25'b11110001_10101010_10011011_1;
      patterns[61869] = 25'b11110001_10101011_10011100_1;
      patterns[61870] = 25'b11110001_10101100_10011101_1;
      patterns[61871] = 25'b11110001_10101101_10011110_1;
      patterns[61872] = 25'b11110001_10101110_10011111_1;
      patterns[61873] = 25'b11110001_10101111_10100000_1;
      patterns[61874] = 25'b11110001_10110000_10100001_1;
      patterns[61875] = 25'b11110001_10110001_10100010_1;
      patterns[61876] = 25'b11110001_10110010_10100011_1;
      patterns[61877] = 25'b11110001_10110011_10100100_1;
      patterns[61878] = 25'b11110001_10110100_10100101_1;
      patterns[61879] = 25'b11110001_10110101_10100110_1;
      patterns[61880] = 25'b11110001_10110110_10100111_1;
      patterns[61881] = 25'b11110001_10110111_10101000_1;
      patterns[61882] = 25'b11110001_10111000_10101001_1;
      patterns[61883] = 25'b11110001_10111001_10101010_1;
      patterns[61884] = 25'b11110001_10111010_10101011_1;
      patterns[61885] = 25'b11110001_10111011_10101100_1;
      patterns[61886] = 25'b11110001_10111100_10101101_1;
      patterns[61887] = 25'b11110001_10111101_10101110_1;
      patterns[61888] = 25'b11110001_10111110_10101111_1;
      patterns[61889] = 25'b11110001_10111111_10110000_1;
      patterns[61890] = 25'b11110001_11000000_10110001_1;
      patterns[61891] = 25'b11110001_11000001_10110010_1;
      patterns[61892] = 25'b11110001_11000010_10110011_1;
      patterns[61893] = 25'b11110001_11000011_10110100_1;
      patterns[61894] = 25'b11110001_11000100_10110101_1;
      patterns[61895] = 25'b11110001_11000101_10110110_1;
      patterns[61896] = 25'b11110001_11000110_10110111_1;
      patterns[61897] = 25'b11110001_11000111_10111000_1;
      patterns[61898] = 25'b11110001_11001000_10111001_1;
      patterns[61899] = 25'b11110001_11001001_10111010_1;
      patterns[61900] = 25'b11110001_11001010_10111011_1;
      patterns[61901] = 25'b11110001_11001011_10111100_1;
      patterns[61902] = 25'b11110001_11001100_10111101_1;
      patterns[61903] = 25'b11110001_11001101_10111110_1;
      patterns[61904] = 25'b11110001_11001110_10111111_1;
      patterns[61905] = 25'b11110001_11001111_11000000_1;
      patterns[61906] = 25'b11110001_11010000_11000001_1;
      patterns[61907] = 25'b11110001_11010001_11000010_1;
      patterns[61908] = 25'b11110001_11010010_11000011_1;
      patterns[61909] = 25'b11110001_11010011_11000100_1;
      patterns[61910] = 25'b11110001_11010100_11000101_1;
      patterns[61911] = 25'b11110001_11010101_11000110_1;
      patterns[61912] = 25'b11110001_11010110_11000111_1;
      patterns[61913] = 25'b11110001_11010111_11001000_1;
      patterns[61914] = 25'b11110001_11011000_11001001_1;
      patterns[61915] = 25'b11110001_11011001_11001010_1;
      patterns[61916] = 25'b11110001_11011010_11001011_1;
      patterns[61917] = 25'b11110001_11011011_11001100_1;
      patterns[61918] = 25'b11110001_11011100_11001101_1;
      patterns[61919] = 25'b11110001_11011101_11001110_1;
      patterns[61920] = 25'b11110001_11011110_11001111_1;
      patterns[61921] = 25'b11110001_11011111_11010000_1;
      patterns[61922] = 25'b11110001_11100000_11010001_1;
      patterns[61923] = 25'b11110001_11100001_11010010_1;
      patterns[61924] = 25'b11110001_11100010_11010011_1;
      patterns[61925] = 25'b11110001_11100011_11010100_1;
      patterns[61926] = 25'b11110001_11100100_11010101_1;
      patterns[61927] = 25'b11110001_11100101_11010110_1;
      patterns[61928] = 25'b11110001_11100110_11010111_1;
      patterns[61929] = 25'b11110001_11100111_11011000_1;
      patterns[61930] = 25'b11110001_11101000_11011001_1;
      patterns[61931] = 25'b11110001_11101001_11011010_1;
      patterns[61932] = 25'b11110001_11101010_11011011_1;
      patterns[61933] = 25'b11110001_11101011_11011100_1;
      patterns[61934] = 25'b11110001_11101100_11011101_1;
      patterns[61935] = 25'b11110001_11101101_11011110_1;
      patterns[61936] = 25'b11110001_11101110_11011111_1;
      patterns[61937] = 25'b11110001_11101111_11100000_1;
      patterns[61938] = 25'b11110001_11110000_11100001_1;
      patterns[61939] = 25'b11110001_11110001_11100010_1;
      patterns[61940] = 25'b11110001_11110010_11100011_1;
      patterns[61941] = 25'b11110001_11110011_11100100_1;
      patterns[61942] = 25'b11110001_11110100_11100101_1;
      patterns[61943] = 25'b11110001_11110101_11100110_1;
      patterns[61944] = 25'b11110001_11110110_11100111_1;
      patterns[61945] = 25'b11110001_11110111_11101000_1;
      patterns[61946] = 25'b11110001_11111000_11101001_1;
      patterns[61947] = 25'b11110001_11111001_11101010_1;
      patterns[61948] = 25'b11110001_11111010_11101011_1;
      patterns[61949] = 25'b11110001_11111011_11101100_1;
      patterns[61950] = 25'b11110001_11111100_11101101_1;
      patterns[61951] = 25'b11110001_11111101_11101110_1;
      patterns[61952] = 25'b11110001_11111110_11101111_1;
      patterns[61953] = 25'b11110001_11111111_11110000_1;
      patterns[61954] = 25'b11110010_00000000_11110010_0;
      patterns[61955] = 25'b11110010_00000001_11110011_0;
      patterns[61956] = 25'b11110010_00000010_11110100_0;
      patterns[61957] = 25'b11110010_00000011_11110101_0;
      patterns[61958] = 25'b11110010_00000100_11110110_0;
      patterns[61959] = 25'b11110010_00000101_11110111_0;
      patterns[61960] = 25'b11110010_00000110_11111000_0;
      patterns[61961] = 25'b11110010_00000111_11111001_0;
      patterns[61962] = 25'b11110010_00001000_11111010_0;
      patterns[61963] = 25'b11110010_00001001_11111011_0;
      patterns[61964] = 25'b11110010_00001010_11111100_0;
      patterns[61965] = 25'b11110010_00001011_11111101_0;
      patterns[61966] = 25'b11110010_00001100_11111110_0;
      patterns[61967] = 25'b11110010_00001101_11111111_0;
      patterns[61968] = 25'b11110010_00001110_00000000_1;
      patterns[61969] = 25'b11110010_00001111_00000001_1;
      patterns[61970] = 25'b11110010_00010000_00000010_1;
      patterns[61971] = 25'b11110010_00010001_00000011_1;
      patterns[61972] = 25'b11110010_00010010_00000100_1;
      patterns[61973] = 25'b11110010_00010011_00000101_1;
      patterns[61974] = 25'b11110010_00010100_00000110_1;
      patterns[61975] = 25'b11110010_00010101_00000111_1;
      patterns[61976] = 25'b11110010_00010110_00001000_1;
      patterns[61977] = 25'b11110010_00010111_00001001_1;
      patterns[61978] = 25'b11110010_00011000_00001010_1;
      patterns[61979] = 25'b11110010_00011001_00001011_1;
      patterns[61980] = 25'b11110010_00011010_00001100_1;
      patterns[61981] = 25'b11110010_00011011_00001101_1;
      patterns[61982] = 25'b11110010_00011100_00001110_1;
      patterns[61983] = 25'b11110010_00011101_00001111_1;
      patterns[61984] = 25'b11110010_00011110_00010000_1;
      patterns[61985] = 25'b11110010_00011111_00010001_1;
      patterns[61986] = 25'b11110010_00100000_00010010_1;
      patterns[61987] = 25'b11110010_00100001_00010011_1;
      patterns[61988] = 25'b11110010_00100010_00010100_1;
      patterns[61989] = 25'b11110010_00100011_00010101_1;
      patterns[61990] = 25'b11110010_00100100_00010110_1;
      patterns[61991] = 25'b11110010_00100101_00010111_1;
      patterns[61992] = 25'b11110010_00100110_00011000_1;
      patterns[61993] = 25'b11110010_00100111_00011001_1;
      patterns[61994] = 25'b11110010_00101000_00011010_1;
      patterns[61995] = 25'b11110010_00101001_00011011_1;
      patterns[61996] = 25'b11110010_00101010_00011100_1;
      patterns[61997] = 25'b11110010_00101011_00011101_1;
      patterns[61998] = 25'b11110010_00101100_00011110_1;
      patterns[61999] = 25'b11110010_00101101_00011111_1;
      patterns[62000] = 25'b11110010_00101110_00100000_1;
      patterns[62001] = 25'b11110010_00101111_00100001_1;
      patterns[62002] = 25'b11110010_00110000_00100010_1;
      patterns[62003] = 25'b11110010_00110001_00100011_1;
      patterns[62004] = 25'b11110010_00110010_00100100_1;
      patterns[62005] = 25'b11110010_00110011_00100101_1;
      patterns[62006] = 25'b11110010_00110100_00100110_1;
      patterns[62007] = 25'b11110010_00110101_00100111_1;
      patterns[62008] = 25'b11110010_00110110_00101000_1;
      patterns[62009] = 25'b11110010_00110111_00101001_1;
      patterns[62010] = 25'b11110010_00111000_00101010_1;
      patterns[62011] = 25'b11110010_00111001_00101011_1;
      patterns[62012] = 25'b11110010_00111010_00101100_1;
      patterns[62013] = 25'b11110010_00111011_00101101_1;
      patterns[62014] = 25'b11110010_00111100_00101110_1;
      patterns[62015] = 25'b11110010_00111101_00101111_1;
      patterns[62016] = 25'b11110010_00111110_00110000_1;
      patterns[62017] = 25'b11110010_00111111_00110001_1;
      patterns[62018] = 25'b11110010_01000000_00110010_1;
      patterns[62019] = 25'b11110010_01000001_00110011_1;
      patterns[62020] = 25'b11110010_01000010_00110100_1;
      patterns[62021] = 25'b11110010_01000011_00110101_1;
      patterns[62022] = 25'b11110010_01000100_00110110_1;
      patterns[62023] = 25'b11110010_01000101_00110111_1;
      patterns[62024] = 25'b11110010_01000110_00111000_1;
      patterns[62025] = 25'b11110010_01000111_00111001_1;
      patterns[62026] = 25'b11110010_01001000_00111010_1;
      patterns[62027] = 25'b11110010_01001001_00111011_1;
      patterns[62028] = 25'b11110010_01001010_00111100_1;
      patterns[62029] = 25'b11110010_01001011_00111101_1;
      patterns[62030] = 25'b11110010_01001100_00111110_1;
      patterns[62031] = 25'b11110010_01001101_00111111_1;
      patterns[62032] = 25'b11110010_01001110_01000000_1;
      patterns[62033] = 25'b11110010_01001111_01000001_1;
      patterns[62034] = 25'b11110010_01010000_01000010_1;
      patterns[62035] = 25'b11110010_01010001_01000011_1;
      patterns[62036] = 25'b11110010_01010010_01000100_1;
      patterns[62037] = 25'b11110010_01010011_01000101_1;
      patterns[62038] = 25'b11110010_01010100_01000110_1;
      patterns[62039] = 25'b11110010_01010101_01000111_1;
      patterns[62040] = 25'b11110010_01010110_01001000_1;
      patterns[62041] = 25'b11110010_01010111_01001001_1;
      patterns[62042] = 25'b11110010_01011000_01001010_1;
      patterns[62043] = 25'b11110010_01011001_01001011_1;
      patterns[62044] = 25'b11110010_01011010_01001100_1;
      patterns[62045] = 25'b11110010_01011011_01001101_1;
      patterns[62046] = 25'b11110010_01011100_01001110_1;
      patterns[62047] = 25'b11110010_01011101_01001111_1;
      patterns[62048] = 25'b11110010_01011110_01010000_1;
      patterns[62049] = 25'b11110010_01011111_01010001_1;
      patterns[62050] = 25'b11110010_01100000_01010010_1;
      patterns[62051] = 25'b11110010_01100001_01010011_1;
      patterns[62052] = 25'b11110010_01100010_01010100_1;
      patterns[62053] = 25'b11110010_01100011_01010101_1;
      patterns[62054] = 25'b11110010_01100100_01010110_1;
      patterns[62055] = 25'b11110010_01100101_01010111_1;
      patterns[62056] = 25'b11110010_01100110_01011000_1;
      patterns[62057] = 25'b11110010_01100111_01011001_1;
      patterns[62058] = 25'b11110010_01101000_01011010_1;
      patterns[62059] = 25'b11110010_01101001_01011011_1;
      patterns[62060] = 25'b11110010_01101010_01011100_1;
      patterns[62061] = 25'b11110010_01101011_01011101_1;
      patterns[62062] = 25'b11110010_01101100_01011110_1;
      patterns[62063] = 25'b11110010_01101101_01011111_1;
      patterns[62064] = 25'b11110010_01101110_01100000_1;
      patterns[62065] = 25'b11110010_01101111_01100001_1;
      patterns[62066] = 25'b11110010_01110000_01100010_1;
      patterns[62067] = 25'b11110010_01110001_01100011_1;
      patterns[62068] = 25'b11110010_01110010_01100100_1;
      patterns[62069] = 25'b11110010_01110011_01100101_1;
      patterns[62070] = 25'b11110010_01110100_01100110_1;
      patterns[62071] = 25'b11110010_01110101_01100111_1;
      patterns[62072] = 25'b11110010_01110110_01101000_1;
      patterns[62073] = 25'b11110010_01110111_01101001_1;
      patterns[62074] = 25'b11110010_01111000_01101010_1;
      patterns[62075] = 25'b11110010_01111001_01101011_1;
      patterns[62076] = 25'b11110010_01111010_01101100_1;
      patterns[62077] = 25'b11110010_01111011_01101101_1;
      patterns[62078] = 25'b11110010_01111100_01101110_1;
      patterns[62079] = 25'b11110010_01111101_01101111_1;
      patterns[62080] = 25'b11110010_01111110_01110000_1;
      patterns[62081] = 25'b11110010_01111111_01110001_1;
      patterns[62082] = 25'b11110010_10000000_01110010_1;
      patterns[62083] = 25'b11110010_10000001_01110011_1;
      patterns[62084] = 25'b11110010_10000010_01110100_1;
      patterns[62085] = 25'b11110010_10000011_01110101_1;
      patterns[62086] = 25'b11110010_10000100_01110110_1;
      patterns[62087] = 25'b11110010_10000101_01110111_1;
      patterns[62088] = 25'b11110010_10000110_01111000_1;
      patterns[62089] = 25'b11110010_10000111_01111001_1;
      patterns[62090] = 25'b11110010_10001000_01111010_1;
      patterns[62091] = 25'b11110010_10001001_01111011_1;
      patterns[62092] = 25'b11110010_10001010_01111100_1;
      patterns[62093] = 25'b11110010_10001011_01111101_1;
      patterns[62094] = 25'b11110010_10001100_01111110_1;
      patterns[62095] = 25'b11110010_10001101_01111111_1;
      patterns[62096] = 25'b11110010_10001110_10000000_1;
      patterns[62097] = 25'b11110010_10001111_10000001_1;
      patterns[62098] = 25'b11110010_10010000_10000010_1;
      patterns[62099] = 25'b11110010_10010001_10000011_1;
      patterns[62100] = 25'b11110010_10010010_10000100_1;
      patterns[62101] = 25'b11110010_10010011_10000101_1;
      patterns[62102] = 25'b11110010_10010100_10000110_1;
      patterns[62103] = 25'b11110010_10010101_10000111_1;
      patterns[62104] = 25'b11110010_10010110_10001000_1;
      patterns[62105] = 25'b11110010_10010111_10001001_1;
      patterns[62106] = 25'b11110010_10011000_10001010_1;
      patterns[62107] = 25'b11110010_10011001_10001011_1;
      patterns[62108] = 25'b11110010_10011010_10001100_1;
      patterns[62109] = 25'b11110010_10011011_10001101_1;
      patterns[62110] = 25'b11110010_10011100_10001110_1;
      patterns[62111] = 25'b11110010_10011101_10001111_1;
      patterns[62112] = 25'b11110010_10011110_10010000_1;
      patterns[62113] = 25'b11110010_10011111_10010001_1;
      patterns[62114] = 25'b11110010_10100000_10010010_1;
      patterns[62115] = 25'b11110010_10100001_10010011_1;
      patterns[62116] = 25'b11110010_10100010_10010100_1;
      patterns[62117] = 25'b11110010_10100011_10010101_1;
      patterns[62118] = 25'b11110010_10100100_10010110_1;
      patterns[62119] = 25'b11110010_10100101_10010111_1;
      patterns[62120] = 25'b11110010_10100110_10011000_1;
      patterns[62121] = 25'b11110010_10100111_10011001_1;
      patterns[62122] = 25'b11110010_10101000_10011010_1;
      patterns[62123] = 25'b11110010_10101001_10011011_1;
      patterns[62124] = 25'b11110010_10101010_10011100_1;
      patterns[62125] = 25'b11110010_10101011_10011101_1;
      patterns[62126] = 25'b11110010_10101100_10011110_1;
      patterns[62127] = 25'b11110010_10101101_10011111_1;
      patterns[62128] = 25'b11110010_10101110_10100000_1;
      patterns[62129] = 25'b11110010_10101111_10100001_1;
      patterns[62130] = 25'b11110010_10110000_10100010_1;
      patterns[62131] = 25'b11110010_10110001_10100011_1;
      patterns[62132] = 25'b11110010_10110010_10100100_1;
      patterns[62133] = 25'b11110010_10110011_10100101_1;
      patterns[62134] = 25'b11110010_10110100_10100110_1;
      patterns[62135] = 25'b11110010_10110101_10100111_1;
      patterns[62136] = 25'b11110010_10110110_10101000_1;
      patterns[62137] = 25'b11110010_10110111_10101001_1;
      patterns[62138] = 25'b11110010_10111000_10101010_1;
      patterns[62139] = 25'b11110010_10111001_10101011_1;
      patterns[62140] = 25'b11110010_10111010_10101100_1;
      patterns[62141] = 25'b11110010_10111011_10101101_1;
      patterns[62142] = 25'b11110010_10111100_10101110_1;
      patterns[62143] = 25'b11110010_10111101_10101111_1;
      patterns[62144] = 25'b11110010_10111110_10110000_1;
      patterns[62145] = 25'b11110010_10111111_10110001_1;
      patterns[62146] = 25'b11110010_11000000_10110010_1;
      patterns[62147] = 25'b11110010_11000001_10110011_1;
      patterns[62148] = 25'b11110010_11000010_10110100_1;
      patterns[62149] = 25'b11110010_11000011_10110101_1;
      patterns[62150] = 25'b11110010_11000100_10110110_1;
      patterns[62151] = 25'b11110010_11000101_10110111_1;
      patterns[62152] = 25'b11110010_11000110_10111000_1;
      patterns[62153] = 25'b11110010_11000111_10111001_1;
      patterns[62154] = 25'b11110010_11001000_10111010_1;
      patterns[62155] = 25'b11110010_11001001_10111011_1;
      patterns[62156] = 25'b11110010_11001010_10111100_1;
      patterns[62157] = 25'b11110010_11001011_10111101_1;
      patterns[62158] = 25'b11110010_11001100_10111110_1;
      patterns[62159] = 25'b11110010_11001101_10111111_1;
      patterns[62160] = 25'b11110010_11001110_11000000_1;
      patterns[62161] = 25'b11110010_11001111_11000001_1;
      patterns[62162] = 25'b11110010_11010000_11000010_1;
      patterns[62163] = 25'b11110010_11010001_11000011_1;
      patterns[62164] = 25'b11110010_11010010_11000100_1;
      patterns[62165] = 25'b11110010_11010011_11000101_1;
      patterns[62166] = 25'b11110010_11010100_11000110_1;
      patterns[62167] = 25'b11110010_11010101_11000111_1;
      patterns[62168] = 25'b11110010_11010110_11001000_1;
      patterns[62169] = 25'b11110010_11010111_11001001_1;
      patterns[62170] = 25'b11110010_11011000_11001010_1;
      patterns[62171] = 25'b11110010_11011001_11001011_1;
      patterns[62172] = 25'b11110010_11011010_11001100_1;
      patterns[62173] = 25'b11110010_11011011_11001101_1;
      patterns[62174] = 25'b11110010_11011100_11001110_1;
      patterns[62175] = 25'b11110010_11011101_11001111_1;
      patterns[62176] = 25'b11110010_11011110_11010000_1;
      patterns[62177] = 25'b11110010_11011111_11010001_1;
      patterns[62178] = 25'b11110010_11100000_11010010_1;
      patterns[62179] = 25'b11110010_11100001_11010011_1;
      patterns[62180] = 25'b11110010_11100010_11010100_1;
      patterns[62181] = 25'b11110010_11100011_11010101_1;
      patterns[62182] = 25'b11110010_11100100_11010110_1;
      patterns[62183] = 25'b11110010_11100101_11010111_1;
      patterns[62184] = 25'b11110010_11100110_11011000_1;
      patterns[62185] = 25'b11110010_11100111_11011001_1;
      patterns[62186] = 25'b11110010_11101000_11011010_1;
      patterns[62187] = 25'b11110010_11101001_11011011_1;
      patterns[62188] = 25'b11110010_11101010_11011100_1;
      patterns[62189] = 25'b11110010_11101011_11011101_1;
      patterns[62190] = 25'b11110010_11101100_11011110_1;
      patterns[62191] = 25'b11110010_11101101_11011111_1;
      patterns[62192] = 25'b11110010_11101110_11100000_1;
      patterns[62193] = 25'b11110010_11101111_11100001_1;
      patterns[62194] = 25'b11110010_11110000_11100010_1;
      patterns[62195] = 25'b11110010_11110001_11100011_1;
      patterns[62196] = 25'b11110010_11110010_11100100_1;
      patterns[62197] = 25'b11110010_11110011_11100101_1;
      patterns[62198] = 25'b11110010_11110100_11100110_1;
      patterns[62199] = 25'b11110010_11110101_11100111_1;
      patterns[62200] = 25'b11110010_11110110_11101000_1;
      patterns[62201] = 25'b11110010_11110111_11101001_1;
      patterns[62202] = 25'b11110010_11111000_11101010_1;
      patterns[62203] = 25'b11110010_11111001_11101011_1;
      patterns[62204] = 25'b11110010_11111010_11101100_1;
      patterns[62205] = 25'b11110010_11111011_11101101_1;
      patterns[62206] = 25'b11110010_11111100_11101110_1;
      patterns[62207] = 25'b11110010_11111101_11101111_1;
      patterns[62208] = 25'b11110010_11111110_11110000_1;
      patterns[62209] = 25'b11110010_11111111_11110001_1;
      patterns[62210] = 25'b11110011_00000000_11110011_0;
      patterns[62211] = 25'b11110011_00000001_11110100_0;
      patterns[62212] = 25'b11110011_00000010_11110101_0;
      patterns[62213] = 25'b11110011_00000011_11110110_0;
      patterns[62214] = 25'b11110011_00000100_11110111_0;
      patterns[62215] = 25'b11110011_00000101_11111000_0;
      patterns[62216] = 25'b11110011_00000110_11111001_0;
      patterns[62217] = 25'b11110011_00000111_11111010_0;
      patterns[62218] = 25'b11110011_00001000_11111011_0;
      patterns[62219] = 25'b11110011_00001001_11111100_0;
      patterns[62220] = 25'b11110011_00001010_11111101_0;
      patterns[62221] = 25'b11110011_00001011_11111110_0;
      patterns[62222] = 25'b11110011_00001100_11111111_0;
      patterns[62223] = 25'b11110011_00001101_00000000_1;
      patterns[62224] = 25'b11110011_00001110_00000001_1;
      patterns[62225] = 25'b11110011_00001111_00000010_1;
      patterns[62226] = 25'b11110011_00010000_00000011_1;
      patterns[62227] = 25'b11110011_00010001_00000100_1;
      patterns[62228] = 25'b11110011_00010010_00000101_1;
      patterns[62229] = 25'b11110011_00010011_00000110_1;
      patterns[62230] = 25'b11110011_00010100_00000111_1;
      patterns[62231] = 25'b11110011_00010101_00001000_1;
      patterns[62232] = 25'b11110011_00010110_00001001_1;
      patterns[62233] = 25'b11110011_00010111_00001010_1;
      patterns[62234] = 25'b11110011_00011000_00001011_1;
      patterns[62235] = 25'b11110011_00011001_00001100_1;
      patterns[62236] = 25'b11110011_00011010_00001101_1;
      patterns[62237] = 25'b11110011_00011011_00001110_1;
      patterns[62238] = 25'b11110011_00011100_00001111_1;
      patterns[62239] = 25'b11110011_00011101_00010000_1;
      patterns[62240] = 25'b11110011_00011110_00010001_1;
      patterns[62241] = 25'b11110011_00011111_00010010_1;
      patterns[62242] = 25'b11110011_00100000_00010011_1;
      patterns[62243] = 25'b11110011_00100001_00010100_1;
      patterns[62244] = 25'b11110011_00100010_00010101_1;
      patterns[62245] = 25'b11110011_00100011_00010110_1;
      patterns[62246] = 25'b11110011_00100100_00010111_1;
      patterns[62247] = 25'b11110011_00100101_00011000_1;
      patterns[62248] = 25'b11110011_00100110_00011001_1;
      patterns[62249] = 25'b11110011_00100111_00011010_1;
      patterns[62250] = 25'b11110011_00101000_00011011_1;
      patterns[62251] = 25'b11110011_00101001_00011100_1;
      patterns[62252] = 25'b11110011_00101010_00011101_1;
      patterns[62253] = 25'b11110011_00101011_00011110_1;
      patterns[62254] = 25'b11110011_00101100_00011111_1;
      patterns[62255] = 25'b11110011_00101101_00100000_1;
      patterns[62256] = 25'b11110011_00101110_00100001_1;
      patterns[62257] = 25'b11110011_00101111_00100010_1;
      patterns[62258] = 25'b11110011_00110000_00100011_1;
      patterns[62259] = 25'b11110011_00110001_00100100_1;
      patterns[62260] = 25'b11110011_00110010_00100101_1;
      patterns[62261] = 25'b11110011_00110011_00100110_1;
      patterns[62262] = 25'b11110011_00110100_00100111_1;
      patterns[62263] = 25'b11110011_00110101_00101000_1;
      patterns[62264] = 25'b11110011_00110110_00101001_1;
      patterns[62265] = 25'b11110011_00110111_00101010_1;
      patterns[62266] = 25'b11110011_00111000_00101011_1;
      patterns[62267] = 25'b11110011_00111001_00101100_1;
      patterns[62268] = 25'b11110011_00111010_00101101_1;
      patterns[62269] = 25'b11110011_00111011_00101110_1;
      patterns[62270] = 25'b11110011_00111100_00101111_1;
      patterns[62271] = 25'b11110011_00111101_00110000_1;
      patterns[62272] = 25'b11110011_00111110_00110001_1;
      patterns[62273] = 25'b11110011_00111111_00110010_1;
      patterns[62274] = 25'b11110011_01000000_00110011_1;
      patterns[62275] = 25'b11110011_01000001_00110100_1;
      patterns[62276] = 25'b11110011_01000010_00110101_1;
      patterns[62277] = 25'b11110011_01000011_00110110_1;
      patterns[62278] = 25'b11110011_01000100_00110111_1;
      patterns[62279] = 25'b11110011_01000101_00111000_1;
      patterns[62280] = 25'b11110011_01000110_00111001_1;
      patterns[62281] = 25'b11110011_01000111_00111010_1;
      patterns[62282] = 25'b11110011_01001000_00111011_1;
      patterns[62283] = 25'b11110011_01001001_00111100_1;
      patterns[62284] = 25'b11110011_01001010_00111101_1;
      patterns[62285] = 25'b11110011_01001011_00111110_1;
      patterns[62286] = 25'b11110011_01001100_00111111_1;
      patterns[62287] = 25'b11110011_01001101_01000000_1;
      patterns[62288] = 25'b11110011_01001110_01000001_1;
      patterns[62289] = 25'b11110011_01001111_01000010_1;
      patterns[62290] = 25'b11110011_01010000_01000011_1;
      patterns[62291] = 25'b11110011_01010001_01000100_1;
      patterns[62292] = 25'b11110011_01010010_01000101_1;
      patterns[62293] = 25'b11110011_01010011_01000110_1;
      patterns[62294] = 25'b11110011_01010100_01000111_1;
      patterns[62295] = 25'b11110011_01010101_01001000_1;
      patterns[62296] = 25'b11110011_01010110_01001001_1;
      patterns[62297] = 25'b11110011_01010111_01001010_1;
      patterns[62298] = 25'b11110011_01011000_01001011_1;
      patterns[62299] = 25'b11110011_01011001_01001100_1;
      patterns[62300] = 25'b11110011_01011010_01001101_1;
      patterns[62301] = 25'b11110011_01011011_01001110_1;
      patterns[62302] = 25'b11110011_01011100_01001111_1;
      patterns[62303] = 25'b11110011_01011101_01010000_1;
      patterns[62304] = 25'b11110011_01011110_01010001_1;
      patterns[62305] = 25'b11110011_01011111_01010010_1;
      patterns[62306] = 25'b11110011_01100000_01010011_1;
      patterns[62307] = 25'b11110011_01100001_01010100_1;
      patterns[62308] = 25'b11110011_01100010_01010101_1;
      patterns[62309] = 25'b11110011_01100011_01010110_1;
      patterns[62310] = 25'b11110011_01100100_01010111_1;
      patterns[62311] = 25'b11110011_01100101_01011000_1;
      patterns[62312] = 25'b11110011_01100110_01011001_1;
      patterns[62313] = 25'b11110011_01100111_01011010_1;
      patterns[62314] = 25'b11110011_01101000_01011011_1;
      patterns[62315] = 25'b11110011_01101001_01011100_1;
      patterns[62316] = 25'b11110011_01101010_01011101_1;
      patterns[62317] = 25'b11110011_01101011_01011110_1;
      patterns[62318] = 25'b11110011_01101100_01011111_1;
      patterns[62319] = 25'b11110011_01101101_01100000_1;
      patterns[62320] = 25'b11110011_01101110_01100001_1;
      patterns[62321] = 25'b11110011_01101111_01100010_1;
      patterns[62322] = 25'b11110011_01110000_01100011_1;
      patterns[62323] = 25'b11110011_01110001_01100100_1;
      patterns[62324] = 25'b11110011_01110010_01100101_1;
      patterns[62325] = 25'b11110011_01110011_01100110_1;
      patterns[62326] = 25'b11110011_01110100_01100111_1;
      patterns[62327] = 25'b11110011_01110101_01101000_1;
      patterns[62328] = 25'b11110011_01110110_01101001_1;
      patterns[62329] = 25'b11110011_01110111_01101010_1;
      patterns[62330] = 25'b11110011_01111000_01101011_1;
      patterns[62331] = 25'b11110011_01111001_01101100_1;
      patterns[62332] = 25'b11110011_01111010_01101101_1;
      patterns[62333] = 25'b11110011_01111011_01101110_1;
      patterns[62334] = 25'b11110011_01111100_01101111_1;
      patterns[62335] = 25'b11110011_01111101_01110000_1;
      patterns[62336] = 25'b11110011_01111110_01110001_1;
      patterns[62337] = 25'b11110011_01111111_01110010_1;
      patterns[62338] = 25'b11110011_10000000_01110011_1;
      patterns[62339] = 25'b11110011_10000001_01110100_1;
      patterns[62340] = 25'b11110011_10000010_01110101_1;
      patterns[62341] = 25'b11110011_10000011_01110110_1;
      patterns[62342] = 25'b11110011_10000100_01110111_1;
      patterns[62343] = 25'b11110011_10000101_01111000_1;
      patterns[62344] = 25'b11110011_10000110_01111001_1;
      patterns[62345] = 25'b11110011_10000111_01111010_1;
      patterns[62346] = 25'b11110011_10001000_01111011_1;
      patterns[62347] = 25'b11110011_10001001_01111100_1;
      patterns[62348] = 25'b11110011_10001010_01111101_1;
      patterns[62349] = 25'b11110011_10001011_01111110_1;
      patterns[62350] = 25'b11110011_10001100_01111111_1;
      patterns[62351] = 25'b11110011_10001101_10000000_1;
      patterns[62352] = 25'b11110011_10001110_10000001_1;
      patterns[62353] = 25'b11110011_10001111_10000010_1;
      patterns[62354] = 25'b11110011_10010000_10000011_1;
      patterns[62355] = 25'b11110011_10010001_10000100_1;
      patterns[62356] = 25'b11110011_10010010_10000101_1;
      patterns[62357] = 25'b11110011_10010011_10000110_1;
      patterns[62358] = 25'b11110011_10010100_10000111_1;
      patterns[62359] = 25'b11110011_10010101_10001000_1;
      patterns[62360] = 25'b11110011_10010110_10001001_1;
      patterns[62361] = 25'b11110011_10010111_10001010_1;
      patterns[62362] = 25'b11110011_10011000_10001011_1;
      patterns[62363] = 25'b11110011_10011001_10001100_1;
      patterns[62364] = 25'b11110011_10011010_10001101_1;
      patterns[62365] = 25'b11110011_10011011_10001110_1;
      patterns[62366] = 25'b11110011_10011100_10001111_1;
      patterns[62367] = 25'b11110011_10011101_10010000_1;
      patterns[62368] = 25'b11110011_10011110_10010001_1;
      patterns[62369] = 25'b11110011_10011111_10010010_1;
      patterns[62370] = 25'b11110011_10100000_10010011_1;
      patterns[62371] = 25'b11110011_10100001_10010100_1;
      patterns[62372] = 25'b11110011_10100010_10010101_1;
      patterns[62373] = 25'b11110011_10100011_10010110_1;
      patterns[62374] = 25'b11110011_10100100_10010111_1;
      patterns[62375] = 25'b11110011_10100101_10011000_1;
      patterns[62376] = 25'b11110011_10100110_10011001_1;
      patterns[62377] = 25'b11110011_10100111_10011010_1;
      patterns[62378] = 25'b11110011_10101000_10011011_1;
      patterns[62379] = 25'b11110011_10101001_10011100_1;
      patterns[62380] = 25'b11110011_10101010_10011101_1;
      patterns[62381] = 25'b11110011_10101011_10011110_1;
      patterns[62382] = 25'b11110011_10101100_10011111_1;
      patterns[62383] = 25'b11110011_10101101_10100000_1;
      patterns[62384] = 25'b11110011_10101110_10100001_1;
      patterns[62385] = 25'b11110011_10101111_10100010_1;
      patterns[62386] = 25'b11110011_10110000_10100011_1;
      patterns[62387] = 25'b11110011_10110001_10100100_1;
      patterns[62388] = 25'b11110011_10110010_10100101_1;
      patterns[62389] = 25'b11110011_10110011_10100110_1;
      patterns[62390] = 25'b11110011_10110100_10100111_1;
      patterns[62391] = 25'b11110011_10110101_10101000_1;
      patterns[62392] = 25'b11110011_10110110_10101001_1;
      patterns[62393] = 25'b11110011_10110111_10101010_1;
      patterns[62394] = 25'b11110011_10111000_10101011_1;
      patterns[62395] = 25'b11110011_10111001_10101100_1;
      patterns[62396] = 25'b11110011_10111010_10101101_1;
      patterns[62397] = 25'b11110011_10111011_10101110_1;
      patterns[62398] = 25'b11110011_10111100_10101111_1;
      patterns[62399] = 25'b11110011_10111101_10110000_1;
      patterns[62400] = 25'b11110011_10111110_10110001_1;
      patterns[62401] = 25'b11110011_10111111_10110010_1;
      patterns[62402] = 25'b11110011_11000000_10110011_1;
      patterns[62403] = 25'b11110011_11000001_10110100_1;
      patterns[62404] = 25'b11110011_11000010_10110101_1;
      patterns[62405] = 25'b11110011_11000011_10110110_1;
      patterns[62406] = 25'b11110011_11000100_10110111_1;
      patterns[62407] = 25'b11110011_11000101_10111000_1;
      patterns[62408] = 25'b11110011_11000110_10111001_1;
      patterns[62409] = 25'b11110011_11000111_10111010_1;
      patterns[62410] = 25'b11110011_11001000_10111011_1;
      patterns[62411] = 25'b11110011_11001001_10111100_1;
      patterns[62412] = 25'b11110011_11001010_10111101_1;
      patterns[62413] = 25'b11110011_11001011_10111110_1;
      patterns[62414] = 25'b11110011_11001100_10111111_1;
      patterns[62415] = 25'b11110011_11001101_11000000_1;
      patterns[62416] = 25'b11110011_11001110_11000001_1;
      patterns[62417] = 25'b11110011_11001111_11000010_1;
      patterns[62418] = 25'b11110011_11010000_11000011_1;
      patterns[62419] = 25'b11110011_11010001_11000100_1;
      patterns[62420] = 25'b11110011_11010010_11000101_1;
      patterns[62421] = 25'b11110011_11010011_11000110_1;
      patterns[62422] = 25'b11110011_11010100_11000111_1;
      patterns[62423] = 25'b11110011_11010101_11001000_1;
      patterns[62424] = 25'b11110011_11010110_11001001_1;
      patterns[62425] = 25'b11110011_11010111_11001010_1;
      patterns[62426] = 25'b11110011_11011000_11001011_1;
      patterns[62427] = 25'b11110011_11011001_11001100_1;
      patterns[62428] = 25'b11110011_11011010_11001101_1;
      patterns[62429] = 25'b11110011_11011011_11001110_1;
      patterns[62430] = 25'b11110011_11011100_11001111_1;
      patterns[62431] = 25'b11110011_11011101_11010000_1;
      patterns[62432] = 25'b11110011_11011110_11010001_1;
      patterns[62433] = 25'b11110011_11011111_11010010_1;
      patterns[62434] = 25'b11110011_11100000_11010011_1;
      patterns[62435] = 25'b11110011_11100001_11010100_1;
      patterns[62436] = 25'b11110011_11100010_11010101_1;
      patterns[62437] = 25'b11110011_11100011_11010110_1;
      patterns[62438] = 25'b11110011_11100100_11010111_1;
      patterns[62439] = 25'b11110011_11100101_11011000_1;
      patterns[62440] = 25'b11110011_11100110_11011001_1;
      patterns[62441] = 25'b11110011_11100111_11011010_1;
      patterns[62442] = 25'b11110011_11101000_11011011_1;
      patterns[62443] = 25'b11110011_11101001_11011100_1;
      patterns[62444] = 25'b11110011_11101010_11011101_1;
      patterns[62445] = 25'b11110011_11101011_11011110_1;
      patterns[62446] = 25'b11110011_11101100_11011111_1;
      patterns[62447] = 25'b11110011_11101101_11100000_1;
      patterns[62448] = 25'b11110011_11101110_11100001_1;
      patterns[62449] = 25'b11110011_11101111_11100010_1;
      patterns[62450] = 25'b11110011_11110000_11100011_1;
      patterns[62451] = 25'b11110011_11110001_11100100_1;
      patterns[62452] = 25'b11110011_11110010_11100101_1;
      patterns[62453] = 25'b11110011_11110011_11100110_1;
      patterns[62454] = 25'b11110011_11110100_11100111_1;
      patterns[62455] = 25'b11110011_11110101_11101000_1;
      patterns[62456] = 25'b11110011_11110110_11101001_1;
      patterns[62457] = 25'b11110011_11110111_11101010_1;
      patterns[62458] = 25'b11110011_11111000_11101011_1;
      patterns[62459] = 25'b11110011_11111001_11101100_1;
      patterns[62460] = 25'b11110011_11111010_11101101_1;
      patterns[62461] = 25'b11110011_11111011_11101110_1;
      patterns[62462] = 25'b11110011_11111100_11101111_1;
      patterns[62463] = 25'b11110011_11111101_11110000_1;
      patterns[62464] = 25'b11110011_11111110_11110001_1;
      patterns[62465] = 25'b11110011_11111111_11110010_1;
      patterns[62466] = 25'b11110100_00000000_11110100_0;
      patterns[62467] = 25'b11110100_00000001_11110101_0;
      patterns[62468] = 25'b11110100_00000010_11110110_0;
      patterns[62469] = 25'b11110100_00000011_11110111_0;
      patterns[62470] = 25'b11110100_00000100_11111000_0;
      patterns[62471] = 25'b11110100_00000101_11111001_0;
      patterns[62472] = 25'b11110100_00000110_11111010_0;
      patterns[62473] = 25'b11110100_00000111_11111011_0;
      patterns[62474] = 25'b11110100_00001000_11111100_0;
      patterns[62475] = 25'b11110100_00001001_11111101_0;
      patterns[62476] = 25'b11110100_00001010_11111110_0;
      patterns[62477] = 25'b11110100_00001011_11111111_0;
      patterns[62478] = 25'b11110100_00001100_00000000_1;
      patterns[62479] = 25'b11110100_00001101_00000001_1;
      patterns[62480] = 25'b11110100_00001110_00000010_1;
      patterns[62481] = 25'b11110100_00001111_00000011_1;
      patterns[62482] = 25'b11110100_00010000_00000100_1;
      patterns[62483] = 25'b11110100_00010001_00000101_1;
      patterns[62484] = 25'b11110100_00010010_00000110_1;
      patterns[62485] = 25'b11110100_00010011_00000111_1;
      patterns[62486] = 25'b11110100_00010100_00001000_1;
      patterns[62487] = 25'b11110100_00010101_00001001_1;
      patterns[62488] = 25'b11110100_00010110_00001010_1;
      patterns[62489] = 25'b11110100_00010111_00001011_1;
      patterns[62490] = 25'b11110100_00011000_00001100_1;
      patterns[62491] = 25'b11110100_00011001_00001101_1;
      patterns[62492] = 25'b11110100_00011010_00001110_1;
      patterns[62493] = 25'b11110100_00011011_00001111_1;
      patterns[62494] = 25'b11110100_00011100_00010000_1;
      patterns[62495] = 25'b11110100_00011101_00010001_1;
      patterns[62496] = 25'b11110100_00011110_00010010_1;
      patterns[62497] = 25'b11110100_00011111_00010011_1;
      patterns[62498] = 25'b11110100_00100000_00010100_1;
      patterns[62499] = 25'b11110100_00100001_00010101_1;
      patterns[62500] = 25'b11110100_00100010_00010110_1;
      patterns[62501] = 25'b11110100_00100011_00010111_1;
      patterns[62502] = 25'b11110100_00100100_00011000_1;
      patterns[62503] = 25'b11110100_00100101_00011001_1;
      patterns[62504] = 25'b11110100_00100110_00011010_1;
      patterns[62505] = 25'b11110100_00100111_00011011_1;
      patterns[62506] = 25'b11110100_00101000_00011100_1;
      patterns[62507] = 25'b11110100_00101001_00011101_1;
      patterns[62508] = 25'b11110100_00101010_00011110_1;
      patterns[62509] = 25'b11110100_00101011_00011111_1;
      patterns[62510] = 25'b11110100_00101100_00100000_1;
      patterns[62511] = 25'b11110100_00101101_00100001_1;
      patterns[62512] = 25'b11110100_00101110_00100010_1;
      patterns[62513] = 25'b11110100_00101111_00100011_1;
      patterns[62514] = 25'b11110100_00110000_00100100_1;
      patterns[62515] = 25'b11110100_00110001_00100101_1;
      patterns[62516] = 25'b11110100_00110010_00100110_1;
      patterns[62517] = 25'b11110100_00110011_00100111_1;
      patterns[62518] = 25'b11110100_00110100_00101000_1;
      patterns[62519] = 25'b11110100_00110101_00101001_1;
      patterns[62520] = 25'b11110100_00110110_00101010_1;
      patterns[62521] = 25'b11110100_00110111_00101011_1;
      patterns[62522] = 25'b11110100_00111000_00101100_1;
      patterns[62523] = 25'b11110100_00111001_00101101_1;
      patterns[62524] = 25'b11110100_00111010_00101110_1;
      patterns[62525] = 25'b11110100_00111011_00101111_1;
      patterns[62526] = 25'b11110100_00111100_00110000_1;
      patterns[62527] = 25'b11110100_00111101_00110001_1;
      patterns[62528] = 25'b11110100_00111110_00110010_1;
      patterns[62529] = 25'b11110100_00111111_00110011_1;
      patterns[62530] = 25'b11110100_01000000_00110100_1;
      patterns[62531] = 25'b11110100_01000001_00110101_1;
      patterns[62532] = 25'b11110100_01000010_00110110_1;
      patterns[62533] = 25'b11110100_01000011_00110111_1;
      patterns[62534] = 25'b11110100_01000100_00111000_1;
      patterns[62535] = 25'b11110100_01000101_00111001_1;
      patterns[62536] = 25'b11110100_01000110_00111010_1;
      patterns[62537] = 25'b11110100_01000111_00111011_1;
      patterns[62538] = 25'b11110100_01001000_00111100_1;
      patterns[62539] = 25'b11110100_01001001_00111101_1;
      patterns[62540] = 25'b11110100_01001010_00111110_1;
      patterns[62541] = 25'b11110100_01001011_00111111_1;
      patterns[62542] = 25'b11110100_01001100_01000000_1;
      patterns[62543] = 25'b11110100_01001101_01000001_1;
      patterns[62544] = 25'b11110100_01001110_01000010_1;
      patterns[62545] = 25'b11110100_01001111_01000011_1;
      patterns[62546] = 25'b11110100_01010000_01000100_1;
      patterns[62547] = 25'b11110100_01010001_01000101_1;
      patterns[62548] = 25'b11110100_01010010_01000110_1;
      patterns[62549] = 25'b11110100_01010011_01000111_1;
      patterns[62550] = 25'b11110100_01010100_01001000_1;
      patterns[62551] = 25'b11110100_01010101_01001001_1;
      patterns[62552] = 25'b11110100_01010110_01001010_1;
      patterns[62553] = 25'b11110100_01010111_01001011_1;
      patterns[62554] = 25'b11110100_01011000_01001100_1;
      patterns[62555] = 25'b11110100_01011001_01001101_1;
      patterns[62556] = 25'b11110100_01011010_01001110_1;
      patterns[62557] = 25'b11110100_01011011_01001111_1;
      patterns[62558] = 25'b11110100_01011100_01010000_1;
      patterns[62559] = 25'b11110100_01011101_01010001_1;
      patterns[62560] = 25'b11110100_01011110_01010010_1;
      patterns[62561] = 25'b11110100_01011111_01010011_1;
      patterns[62562] = 25'b11110100_01100000_01010100_1;
      patterns[62563] = 25'b11110100_01100001_01010101_1;
      patterns[62564] = 25'b11110100_01100010_01010110_1;
      patterns[62565] = 25'b11110100_01100011_01010111_1;
      patterns[62566] = 25'b11110100_01100100_01011000_1;
      patterns[62567] = 25'b11110100_01100101_01011001_1;
      patterns[62568] = 25'b11110100_01100110_01011010_1;
      patterns[62569] = 25'b11110100_01100111_01011011_1;
      patterns[62570] = 25'b11110100_01101000_01011100_1;
      patterns[62571] = 25'b11110100_01101001_01011101_1;
      patterns[62572] = 25'b11110100_01101010_01011110_1;
      patterns[62573] = 25'b11110100_01101011_01011111_1;
      patterns[62574] = 25'b11110100_01101100_01100000_1;
      patterns[62575] = 25'b11110100_01101101_01100001_1;
      patterns[62576] = 25'b11110100_01101110_01100010_1;
      patterns[62577] = 25'b11110100_01101111_01100011_1;
      patterns[62578] = 25'b11110100_01110000_01100100_1;
      patterns[62579] = 25'b11110100_01110001_01100101_1;
      patterns[62580] = 25'b11110100_01110010_01100110_1;
      patterns[62581] = 25'b11110100_01110011_01100111_1;
      patterns[62582] = 25'b11110100_01110100_01101000_1;
      patterns[62583] = 25'b11110100_01110101_01101001_1;
      patterns[62584] = 25'b11110100_01110110_01101010_1;
      patterns[62585] = 25'b11110100_01110111_01101011_1;
      patterns[62586] = 25'b11110100_01111000_01101100_1;
      patterns[62587] = 25'b11110100_01111001_01101101_1;
      patterns[62588] = 25'b11110100_01111010_01101110_1;
      patterns[62589] = 25'b11110100_01111011_01101111_1;
      patterns[62590] = 25'b11110100_01111100_01110000_1;
      patterns[62591] = 25'b11110100_01111101_01110001_1;
      patterns[62592] = 25'b11110100_01111110_01110010_1;
      patterns[62593] = 25'b11110100_01111111_01110011_1;
      patterns[62594] = 25'b11110100_10000000_01110100_1;
      patterns[62595] = 25'b11110100_10000001_01110101_1;
      patterns[62596] = 25'b11110100_10000010_01110110_1;
      patterns[62597] = 25'b11110100_10000011_01110111_1;
      patterns[62598] = 25'b11110100_10000100_01111000_1;
      patterns[62599] = 25'b11110100_10000101_01111001_1;
      patterns[62600] = 25'b11110100_10000110_01111010_1;
      patterns[62601] = 25'b11110100_10000111_01111011_1;
      patterns[62602] = 25'b11110100_10001000_01111100_1;
      patterns[62603] = 25'b11110100_10001001_01111101_1;
      patterns[62604] = 25'b11110100_10001010_01111110_1;
      patterns[62605] = 25'b11110100_10001011_01111111_1;
      patterns[62606] = 25'b11110100_10001100_10000000_1;
      patterns[62607] = 25'b11110100_10001101_10000001_1;
      patterns[62608] = 25'b11110100_10001110_10000010_1;
      patterns[62609] = 25'b11110100_10001111_10000011_1;
      patterns[62610] = 25'b11110100_10010000_10000100_1;
      patterns[62611] = 25'b11110100_10010001_10000101_1;
      patterns[62612] = 25'b11110100_10010010_10000110_1;
      patterns[62613] = 25'b11110100_10010011_10000111_1;
      patterns[62614] = 25'b11110100_10010100_10001000_1;
      patterns[62615] = 25'b11110100_10010101_10001001_1;
      patterns[62616] = 25'b11110100_10010110_10001010_1;
      patterns[62617] = 25'b11110100_10010111_10001011_1;
      patterns[62618] = 25'b11110100_10011000_10001100_1;
      patterns[62619] = 25'b11110100_10011001_10001101_1;
      patterns[62620] = 25'b11110100_10011010_10001110_1;
      patterns[62621] = 25'b11110100_10011011_10001111_1;
      patterns[62622] = 25'b11110100_10011100_10010000_1;
      patterns[62623] = 25'b11110100_10011101_10010001_1;
      patterns[62624] = 25'b11110100_10011110_10010010_1;
      patterns[62625] = 25'b11110100_10011111_10010011_1;
      patterns[62626] = 25'b11110100_10100000_10010100_1;
      patterns[62627] = 25'b11110100_10100001_10010101_1;
      patterns[62628] = 25'b11110100_10100010_10010110_1;
      patterns[62629] = 25'b11110100_10100011_10010111_1;
      patterns[62630] = 25'b11110100_10100100_10011000_1;
      patterns[62631] = 25'b11110100_10100101_10011001_1;
      patterns[62632] = 25'b11110100_10100110_10011010_1;
      patterns[62633] = 25'b11110100_10100111_10011011_1;
      patterns[62634] = 25'b11110100_10101000_10011100_1;
      patterns[62635] = 25'b11110100_10101001_10011101_1;
      patterns[62636] = 25'b11110100_10101010_10011110_1;
      patterns[62637] = 25'b11110100_10101011_10011111_1;
      patterns[62638] = 25'b11110100_10101100_10100000_1;
      patterns[62639] = 25'b11110100_10101101_10100001_1;
      patterns[62640] = 25'b11110100_10101110_10100010_1;
      patterns[62641] = 25'b11110100_10101111_10100011_1;
      patterns[62642] = 25'b11110100_10110000_10100100_1;
      patterns[62643] = 25'b11110100_10110001_10100101_1;
      patterns[62644] = 25'b11110100_10110010_10100110_1;
      patterns[62645] = 25'b11110100_10110011_10100111_1;
      patterns[62646] = 25'b11110100_10110100_10101000_1;
      patterns[62647] = 25'b11110100_10110101_10101001_1;
      patterns[62648] = 25'b11110100_10110110_10101010_1;
      patterns[62649] = 25'b11110100_10110111_10101011_1;
      patterns[62650] = 25'b11110100_10111000_10101100_1;
      patterns[62651] = 25'b11110100_10111001_10101101_1;
      patterns[62652] = 25'b11110100_10111010_10101110_1;
      patterns[62653] = 25'b11110100_10111011_10101111_1;
      patterns[62654] = 25'b11110100_10111100_10110000_1;
      patterns[62655] = 25'b11110100_10111101_10110001_1;
      patterns[62656] = 25'b11110100_10111110_10110010_1;
      patterns[62657] = 25'b11110100_10111111_10110011_1;
      patterns[62658] = 25'b11110100_11000000_10110100_1;
      patterns[62659] = 25'b11110100_11000001_10110101_1;
      patterns[62660] = 25'b11110100_11000010_10110110_1;
      patterns[62661] = 25'b11110100_11000011_10110111_1;
      patterns[62662] = 25'b11110100_11000100_10111000_1;
      patterns[62663] = 25'b11110100_11000101_10111001_1;
      patterns[62664] = 25'b11110100_11000110_10111010_1;
      patterns[62665] = 25'b11110100_11000111_10111011_1;
      patterns[62666] = 25'b11110100_11001000_10111100_1;
      patterns[62667] = 25'b11110100_11001001_10111101_1;
      patterns[62668] = 25'b11110100_11001010_10111110_1;
      patterns[62669] = 25'b11110100_11001011_10111111_1;
      patterns[62670] = 25'b11110100_11001100_11000000_1;
      patterns[62671] = 25'b11110100_11001101_11000001_1;
      patterns[62672] = 25'b11110100_11001110_11000010_1;
      patterns[62673] = 25'b11110100_11001111_11000011_1;
      patterns[62674] = 25'b11110100_11010000_11000100_1;
      patterns[62675] = 25'b11110100_11010001_11000101_1;
      patterns[62676] = 25'b11110100_11010010_11000110_1;
      patterns[62677] = 25'b11110100_11010011_11000111_1;
      patterns[62678] = 25'b11110100_11010100_11001000_1;
      patterns[62679] = 25'b11110100_11010101_11001001_1;
      patterns[62680] = 25'b11110100_11010110_11001010_1;
      patterns[62681] = 25'b11110100_11010111_11001011_1;
      patterns[62682] = 25'b11110100_11011000_11001100_1;
      patterns[62683] = 25'b11110100_11011001_11001101_1;
      patterns[62684] = 25'b11110100_11011010_11001110_1;
      patterns[62685] = 25'b11110100_11011011_11001111_1;
      patterns[62686] = 25'b11110100_11011100_11010000_1;
      patterns[62687] = 25'b11110100_11011101_11010001_1;
      patterns[62688] = 25'b11110100_11011110_11010010_1;
      patterns[62689] = 25'b11110100_11011111_11010011_1;
      patterns[62690] = 25'b11110100_11100000_11010100_1;
      patterns[62691] = 25'b11110100_11100001_11010101_1;
      patterns[62692] = 25'b11110100_11100010_11010110_1;
      patterns[62693] = 25'b11110100_11100011_11010111_1;
      patterns[62694] = 25'b11110100_11100100_11011000_1;
      patterns[62695] = 25'b11110100_11100101_11011001_1;
      patterns[62696] = 25'b11110100_11100110_11011010_1;
      patterns[62697] = 25'b11110100_11100111_11011011_1;
      patterns[62698] = 25'b11110100_11101000_11011100_1;
      patterns[62699] = 25'b11110100_11101001_11011101_1;
      patterns[62700] = 25'b11110100_11101010_11011110_1;
      patterns[62701] = 25'b11110100_11101011_11011111_1;
      patterns[62702] = 25'b11110100_11101100_11100000_1;
      patterns[62703] = 25'b11110100_11101101_11100001_1;
      patterns[62704] = 25'b11110100_11101110_11100010_1;
      patterns[62705] = 25'b11110100_11101111_11100011_1;
      patterns[62706] = 25'b11110100_11110000_11100100_1;
      patterns[62707] = 25'b11110100_11110001_11100101_1;
      patterns[62708] = 25'b11110100_11110010_11100110_1;
      patterns[62709] = 25'b11110100_11110011_11100111_1;
      patterns[62710] = 25'b11110100_11110100_11101000_1;
      patterns[62711] = 25'b11110100_11110101_11101001_1;
      patterns[62712] = 25'b11110100_11110110_11101010_1;
      patterns[62713] = 25'b11110100_11110111_11101011_1;
      patterns[62714] = 25'b11110100_11111000_11101100_1;
      patterns[62715] = 25'b11110100_11111001_11101101_1;
      patterns[62716] = 25'b11110100_11111010_11101110_1;
      patterns[62717] = 25'b11110100_11111011_11101111_1;
      patterns[62718] = 25'b11110100_11111100_11110000_1;
      patterns[62719] = 25'b11110100_11111101_11110001_1;
      patterns[62720] = 25'b11110100_11111110_11110010_1;
      patterns[62721] = 25'b11110100_11111111_11110011_1;
      patterns[62722] = 25'b11110101_00000000_11110101_0;
      patterns[62723] = 25'b11110101_00000001_11110110_0;
      patterns[62724] = 25'b11110101_00000010_11110111_0;
      patterns[62725] = 25'b11110101_00000011_11111000_0;
      patterns[62726] = 25'b11110101_00000100_11111001_0;
      patterns[62727] = 25'b11110101_00000101_11111010_0;
      patterns[62728] = 25'b11110101_00000110_11111011_0;
      patterns[62729] = 25'b11110101_00000111_11111100_0;
      patterns[62730] = 25'b11110101_00001000_11111101_0;
      patterns[62731] = 25'b11110101_00001001_11111110_0;
      patterns[62732] = 25'b11110101_00001010_11111111_0;
      patterns[62733] = 25'b11110101_00001011_00000000_1;
      patterns[62734] = 25'b11110101_00001100_00000001_1;
      patterns[62735] = 25'b11110101_00001101_00000010_1;
      patterns[62736] = 25'b11110101_00001110_00000011_1;
      patterns[62737] = 25'b11110101_00001111_00000100_1;
      patterns[62738] = 25'b11110101_00010000_00000101_1;
      patterns[62739] = 25'b11110101_00010001_00000110_1;
      patterns[62740] = 25'b11110101_00010010_00000111_1;
      patterns[62741] = 25'b11110101_00010011_00001000_1;
      patterns[62742] = 25'b11110101_00010100_00001001_1;
      patterns[62743] = 25'b11110101_00010101_00001010_1;
      patterns[62744] = 25'b11110101_00010110_00001011_1;
      patterns[62745] = 25'b11110101_00010111_00001100_1;
      patterns[62746] = 25'b11110101_00011000_00001101_1;
      patterns[62747] = 25'b11110101_00011001_00001110_1;
      patterns[62748] = 25'b11110101_00011010_00001111_1;
      patterns[62749] = 25'b11110101_00011011_00010000_1;
      patterns[62750] = 25'b11110101_00011100_00010001_1;
      patterns[62751] = 25'b11110101_00011101_00010010_1;
      patterns[62752] = 25'b11110101_00011110_00010011_1;
      patterns[62753] = 25'b11110101_00011111_00010100_1;
      patterns[62754] = 25'b11110101_00100000_00010101_1;
      patterns[62755] = 25'b11110101_00100001_00010110_1;
      patterns[62756] = 25'b11110101_00100010_00010111_1;
      patterns[62757] = 25'b11110101_00100011_00011000_1;
      patterns[62758] = 25'b11110101_00100100_00011001_1;
      patterns[62759] = 25'b11110101_00100101_00011010_1;
      patterns[62760] = 25'b11110101_00100110_00011011_1;
      patterns[62761] = 25'b11110101_00100111_00011100_1;
      patterns[62762] = 25'b11110101_00101000_00011101_1;
      patterns[62763] = 25'b11110101_00101001_00011110_1;
      patterns[62764] = 25'b11110101_00101010_00011111_1;
      patterns[62765] = 25'b11110101_00101011_00100000_1;
      patterns[62766] = 25'b11110101_00101100_00100001_1;
      patterns[62767] = 25'b11110101_00101101_00100010_1;
      patterns[62768] = 25'b11110101_00101110_00100011_1;
      patterns[62769] = 25'b11110101_00101111_00100100_1;
      patterns[62770] = 25'b11110101_00110000_00100101_1;
      patterns[62771] = 25'b11110101_00110001_00100110_1;
      patterns[62772] = 25'b11110101_00110010_00100111_1;
      patterns[62773] = 25'b11110101_00110011_00101000_1;
      patterns[62774] = 25'b11110101_00110100_00101001_1;
      patterns[62775] = 25'b11110101_00110101_00101010_1;
      patterns[62776] = 25'b11110101_00110110_00101011_1;
      patterns[62777] = 25'b11110101_00110111_00101100_1;
      patterns[62778] = 25'b11110101_00111000_00101101_1;
      patterns[62779] = 25'b11110101_00111001_00101110_1;
      patterns[62780] = 25'b11110101_00111010_00101111_1;
      patterns[62781] = 25'b11110101_00111011_00110000_1;
      patterns[62782] = 25'b11110101_00111100_00110001_1;
      patterns[62783] = 25'b11110101_00111101_00110010_1;
      patterns[62784] = 25'b11110101_00111110_00110011_1;
      patterns[62785] = 25'b11110101_00111111_00110100_1;
      patterns[62786] = 25'b11110101_01000000_00110101_1;
      patterns[62787] = 25'b11110101_01000001_00110110_1;
      patterns[62788] = 25'b11110101_01000010_00110111_1;
      patterns[62789] = 25'b11110101_01000011_00111000_1;
      patterns[62790] = 25'b11110101_01000100_00111001_1;
      patterns[62791] = 25'b11110101_01000101_00111010_1;
      patterns[62792] = 25'b11110101_01000110_00111011_1;
      patterns[62793] = 25'b11110101_01000111_00111100_1;
      patterns[62794] = 25'b11110101_01001000_00111101_1;
      patterns[62795] = 25'b11110101_01001001_00111110_1;
      patterns[62796] = 25'b11110101_01001010_00111111_1;
      patterns[62797] = 25'b11110101_01001011_01000000_1;
      patterns[62798] = 25'b11110101_01001100_01000001_1;
      patterns[62799] = 25'b11110101_01001101_01000010_1;
      patterns[62800] = 25'b11110101_01001110_01000011_1;
      patterns[62801] = 25'b11110101_01001111_01000100_1;
      patterns[62802] = 25'b11110101_01010000_01000101_1;
      patterns[62803] = 25'b11110101_01010001_01000110_1;
      patterns[62804] = 25'b11110101_01010010_01000111_1;
      patterns[62805] = 25'b11110101_01010011_01001000_1;
      patterns[62806] = 25'b11110101_01010100_01001001_1;
      patterns[62807] = 25'b11110101_01010101_01001010_1;
      patterns[62808] = 25'b11110101_01010110_01001011_1;
      patterns[62809] = 25'b11110101_01010111_01001100_1;
      patterns[62810] = 25'b11110101_01011000_01001101_1;
      patterns[62811] = 25'b11110101_01011001_01001110_1;
      patterns[62812] = 25'b11110101_01011010_01001111_1;
      patterns[62813] = 25'b11110101_01011011_01010000_1;
      patterns[62814] = 25'b11110101_01011100_01010001_1;
      patterns[62815] = 25'b11110101_01011101_01010010_1;
      patterns[62816] = 25'b11110101_01011110_01010011_1;
      patterns[62817] = 25'b11110101_01011111_01010100_1;
      patterns[62818] = 25'b11110101_01100000_01010101_1;
      patterns[62819] = 25'b11110101_01100001_01010110_1;
      patterns[62820] = 25'b11110101_01100010_01010111_1;
      patterns[62821] = 25'b11110101_01100011_01011000_1;
      patterns[62822] = 25'b11110101_01100100_01011001_1;
      patterns[62823] = 25'b11110101_01100101_01011010_1;
      patterns[62824] = 25'b11110101_01100110_01011011_1;
      patterns[62825] = 25'b11110101_01100111_01011100_1;
      patterns[62826] = 25'b11110101_01101000_01011101_1;
      patterns[62827] = 25'b11110101_01101001_01011110_1;
      patterns[62828] = 25'b11110101_01101010_01011111_1;
      patterns[62829] = 25'b11110101_01101011_01100000_1;
      patterns[62830] = 25'b11110101_01101100_01100001_1;
      patterns[62831] = 25'b11110101_01101101_01100010_1;
      patterns[62832] = 25'b11110101_01101110_01100011_1;
      patterns[62833] = 25'b11110101_01101111_01100100_1;
      patterns[62834] = 25'b11110101_01110000_01100101_1;
      patterns[62835] = 25'b11110101_01110001_01100110_1;
      patterns[62836] = 25'b11110101_01110010_01100111_1;
      patterns[62837] = 25'b11110101_01110011_01101000_1;
      patterns[62838] = 25'b11110101_01110100_01101001_1;
      patterns[62839] = 25'b11110101_01110101_01101010_1;
      patterns[62840] = 25'b11110101_01110110_01101011_1;
      patterns[62841] = 25'b11110101_01110111_01101100_1;
      patterns[62842] = 25'b11110101_01111000_01101101_1;
      patterns[62843] = 25'b11110101_01111001_01101110_1;
      patterns[62844] = 25'b11110101_01111010_01101111_1;
      patterns[62845] = 25'b11110101_01111011_01110000_1;
      patterns[62846] = 25'b11110101_01111100_01110001_1;
      patterns[62847] = 25'b11110101_01111101_01110010_1;
      patterns[62848] = 25'b11110101_01111110_01110011_1;
      patterns[62849] = 25'b11110101_01111111_01110100_1;
      patterns[62850] = 25'b11110101_10000000_01110101_1;
      patterns[62851] = 25'b11110101_10000001_01110110_1;
      patterns[62852] = 25'b11110101_10000010_01110111_1;
      patterns[62853] = 25'b11110101_10000011_01111000_1;
      patterns[62854] = 25'b11110101_10000100_01111001_1;
      patterns[62855] = 25'b11110101_10000101_01111010_1;
      patterns[62856] = 25'b11110101_10000110_01111011_1;
      patterns[62857] = 25'b11110101_10000111_01111100_1;
      patterns[62858] = 25'b11110101_10001000_01111101_1;
      patterns[62859] = 25'b11110101_10001001_01111110_1;
      patterns[62860] = 25'b11110101_10001010_01111111_1;
      patterns[62861] = 25'b11110101_10001011_10000000_1;
      patterns[62862] = 25'b11110101_10001100_10000001_1;
      patterns[62863] = 25'b11110101_10001101_10000010_1;
      patterns[62864] = 25'b11110101_10001110_10000011_1;
      patterns[62865] = 25'b11110101_10001111_10000100_1;
      patterns[62866] = 25'b11110101_10010000_10000101_1;
      patterns[62867] = 25'b11110101_10010001_10000110_1;
      patterns[62868] = 25'b11110101_10010010_10000111_1;
      patterns[62869] = 25'b11110101_10010011_10001000_1;
      patterns[62870] = 25'b11110101_10010100_10001001_1;
      patterns[62871] = 25'b11110101_10010101_10001010_1;
      patterns[62872] = 25'b11110101_10010110_10001011_1;
      patterns[62873] = 25'b11110101_10010111_10001100_1;
      patterns[62874] = 25'b11110101_10011000_10001101_1;
      patterns[62875] = 25'b11110101_10011001_10001110_1;
      patterns[62876] = 25'b11110101_10011010_10001111_1;
      patterns[62877] = 25'b11110101_10011011_10010000_1;
      patterns[62878] = 25'b11110101_10011100_10010001_1;
      patterns[62879] = 25'b11110101_10011101_10010010_1;
      patterns[62880] = 25'b11110101_10011110_10010011_1;
      patterns[62881] = 25'b11110101_10011111_10010100_1;
      patterns[62882] = 25'b11110101_10100000_10010101_1;
      patterns[62883] = 25'b11110101_10100001_10010110_1;
      patterns[62884] = 25'b11110101_10100010_10010111_1;
      patterns[62885] = 25'b11110101_10100011_10011000_1;
      patterns[62886] = 25'b11110101_10100100_10011001_1;
      patterns[62887] = 25'b11110101_10100101_10011010_1;
      patterns[62888] = 25'b11110101_10100110_10011011_1;
      patterns[62889] = 25'b11110101_10100111_10011100_1;
      patterns[62890] = 25'b11110101_10101000_10011101_1;
      patterns[62891] = 25'b11110101_10101001_10011110_1;
      patterns[62892] = 25'b11110101_10101010_10011111_1;
      patterns[62893] = 25'b11110101_10101011_10100000_1;
      patterns[62894] = 25'b11110101_10101100_10100001_1;
      patterns[62895] = 25'b11110101_10101101_10100010_1;
      patterns[62896] = 25'b11110101_10101110_10100011_1;
      patterns[62897] = 25'b11110101_10101111_10100100_1;
      patterns[62898] = 25'b11110101_10110000_10100101_1;
      patterns[62899] = 25'b11110101_10110001_10100110_1;
      patterns[62900] = 25'b11110101_10110010_10100111_1;
      patterns[62901] = 25'b11110101_10110011_10101000_1;
      patterns[62902] = 25'b11110101_10110100_10101001_1;
      patterns[62903] = 25'b11110101_10110101_10101010_1;
      patterns[62904] = 25'b11110101_10110110_10101011_1;
      patterns[62905] = 25'b11110101_10110111_10101100_1;
      patterns[62906] = 25'b11110101_10111000_10101101_1;
      patterns[62907] = 25'b11110101_10111001_10101110_1;
      patterns[62908] = 25'b11110101_10111010_10101111_1;
      patterns[62909] = 25'b11110101_10111011_10110000_1;
      patterns[62910] = 25'b11110101_10111100_10110001_1;
      patterns[62911] = 25'b11110101_10111101_10110010_1;
      patterns[62912] = 25'b11110101_10111110_10110011_1;
      patterns[62913] = 25'b11110101_10111111_10110100_1;
      patterns[62914] = 25'b11110101_11000000_10110101_1;
      patterns[62915] = 25'b11110101_11000001_10110110_1;
      patterns[62916] = 25'b11110101_11000010_10110111_1;
      patterns[62917] = 25'b11110101_11000011_10111000_1;
      patterns[62918] = 25'b11110101_11000100_10111001_1;
      patterns[62919] = 25'b11110101_11000101_10111010_1;
      patterns[62920] = 25'b11110101_11000110_10111011_1;
      patterns[62921] = 25'b11110101_11000111_10111100_1;
      patterns[62922] = 25'b11110101_11001000_10111101_1;
      patterns[62923] = 25'b11110101_11001001_10111110_1;
      patterns[62924] = 25'b11110101_11001010_10111111_1;
      patterns[62925] = 25'b11110101_11001011_11000000_1;
      patterns[62926] = 25'b11110101_11001100_11000001_1;
      patterns[62927] = 25'b11110101_11001101_11000010_1;
      patterns[62928] = 25'b11110101_11001110_11000011_1;
      patterns[62929] = 25'b11110101_11001111_11000100_1;
      patterns[62930] = 25'b11110101_11010000_11000101_1;
      patterns[62931] = 25'b11110101_11010001_11000110_1;
      patterns[62932] = 25'b11110101_11010010_11000111_1;
      patterns[62933] = 25'b11110101_11010011_11001000_1;
      patterns[62934] = 25'b11110101_11010100_11001001_1;
      patterns[62935] = 25'b11110101_11010101_11001010_1;
      patterns[62936] = 25'b11110101_11010110_11001011_1;
      patterns[62937] = 25'b11110101_11010111_11001100_1;
      patterns[62938] = 25'b11110101_11011000_11001101_1;
      patterns[62939] = 25'b11110101_11011001_11001110_1;
      patterns[62940] = 25'b11110101_11011010_11001111_1;
      patterns[62941] = 25'b11110101_11011011_11010000_1;
      patterns[62942] = 25'b11110101_11011100_11010001_1;
      patterns[62943] = 25'b11110101_11011101_11010010_1;
      patterns[62944] = 25'b11110101_11011110_11010011_1;
      patterns[62945] = 25'b11110101_11011111_11010100_1;
      patterns[62946] = 25'b11110101_11100000_11010101_1;
      patterns[62947] = 25'b11110101_11100001_11010110_1;
      patterns[62948] = 25'b11110101_11100010_11010111_1;
      patterns[62949] = 25'b11110101_11100011_11011000_1;
      patterns[62950] = 25'b11110101_11100100_11011001_1;
      patterns[62951] = 25'b11110101_11100101_11011010_1;
      patterns[62952] = 25'b11110101_11100110_11011011_1;
      patterns[62953] = 25'b11110101_11100111_11011100_1;
      patterns[62954] = 25'b11110101_11101000_11011101_1;
      patterns[62955] = 25'b11110101_11101001_11011110_1;
      patterns[62956] = 25'b11110101_11101010_11011111_1;
      patterns[62957] = 25'b11110101_11101011_11100000_1;
      patterns[62958] = 25'b11110101_11101100_11100001_1;
      patterns[62959] = 25'b11110101_11101101_11100010_1;
      patterns[62960] = 25'b11110101_11101110_11100011_1;
      patterns[62961] = 25'b11110101_11101111_11100100_1;
      patterns[62962] = 25'b11110101_11110000_11100101_1;
      patterns[62963] = 25'b11110101_11110001_11100110_1;
      patterns[62964] = 25'b11110101_11110010_11100111_1;
      patterns[62965] = 25'b11110101_11110011_11101000_1;
      patterns[62966] = 25'b11110101_11110100_11101001_1;
      patterns[62967] = 25'b11110101_11110101_11101010_1;
      patterns[62968] = 25'b11110101_11110110_11101011_1;
      patterns[62969] = 25'b11110101_11110111_11101100_1;
      patterns[62970] = 25'b11110101_11111000_11101101_1;
      patterns[62971] = 25'b11110101_11111001_11101110_1;
      patterns[62972] = 25'b11110101_11111010_11101111_1;
      patterns[62973] = 25'b11110101_11111011_11110000_1;
      patterns[62974] = 25'b11110101_11111100_11110001_1;
      patterns[62975] = 25'b11110101_11111101_11110010_1;
      patterns[62976] = 25'b11110101_11111110_11110011_1;
      patterns[62977] = 25'b11110101_11111111_11110100_1;
      patterns[62978] = 25'b11110110_00000000_11110110_0;
      patterns[62979] = 25'b11110110_00000001_11110111_0;
      patterns[62980] = 25'b11110110_00000010_11111000_0;
      patterns[62981] = 25'b11110110_00000011_11111001_0;
      patterns[62982] = 25'b11110110_00000100_11111010_0;
      patterns[62983] = 25'b11110110_00000101_11111011_0;
      patterns[62984] = 25'b11110110_00000110_11111100_0;
      patterns[62985] = 25'b11110110_00000111_11111101_0;
      patterns[62986] = 25'b11110110_00001000_11111110_0;
      patterns[62987] = 25'b11110110_00001001_11111111_0;
      patterns[62988] = 25'b11110110_00001010_00000000_1;
      patterns[62989] = 25'b11110110_00001011_00000001_1;
      patterns[62990] = 25'b11110110_00001100_00000010_1;
      patterns[62991] = 25'b11110110_00001101_00000011_1;
      patterns[62992] = 25'b11110110_00001110_00000100_1;
      patterns[62993] = 25'b11110110_00001111_00000101_1;
      patterns[62994] = 25'b11110110_00010000_00000110_1;
      patterns[62995] = 25'b11110110_00010001_00000111_1;
      patterns[62996] = 25'b11110110_00010010_00001000_1;
      patterns[62997] = 25'b11110110_00010011_00001001_1;
      patterns[62998] = 25'b11110110_00010100_00001010_1;
      patterns[62999] = 25'b11110110_00010101_00001011_1;
      patterns[63000] = 25'b11110110_00010110_00001100_1;
      patterns[63001] = 25'b11110110_00010111_00001101_1;
      patterns[63002] = 25'b11110110_00011000_00001110_1;
      patterns[63003] = 25'b11110110_00011001_00001111_1;
      patterns[63004] = 25'b11110110_00011010_00010000_1;
      patterns[63005] = 25'b11110110_00011011_00010001_1;
      patterns[63006] = 25'b11110110_00011100_00010010_1;
      patterns[63007] = 25'b11110110_00011101_00010011_1;
      patterns[63008] = 25'b11110110_00011110_00010100_1;
      patterns[63009] = 25'b11110110_00011111_00010101_1;
      patterns[63010] = 25'b11110110_00100000_00010110_1;
      patterns[63011] = 25'b11110110_00100001_00010111_1;
      patterns[63012] = 25'b11110110_00100010_00011000_1;
      patterns[63013] = 25'b11110110_00100011_00011001_1;
      patterns[63014] = 25'b11110110_00100100_00011010_1;
      patterns[63015] = 25'b11110110_00100101_00011011_1;
      patterns[63016] = 25'b11110110_00100110_00011100_1;
      patterns[63017] = 25'b11110110_00100111_00011101_1;
      patterns[63018] = 25'b11110110_00101000_00011110_1;
      patterns[63019] = 25'b11110110_00101001_00011111_1;
      patterns[63020] = 25'b11110110_00101010_00100000_1;
      patterns[63021] = 25'b11110110_00101011_00100001_1;
      patterns[63022] = 25'b11110110_00101100_00100010_1;
      patterns[63023] = 25'b11110110_00101101_00100011_1;
      patterns[63024] = 25'b11110110_00101110_00100100_1;
      patterns[63025] = 25'b11110110_00101111_00100101_1;
      patterns[63026] = 25'b11110110_00110000_00100110_1;
      patterns[63027] = 25'b11110110_00110001_00100111_1;
      patterns[63028] = 25'b11110110_00110010_00101000_1;
      patterns[63029] = 25'b11110110_00110011_00101001_1;
      patterns[63030] = 25'b11110110_00110100_00101010_1;
      patterns[63031] = 25'b11110110_00110101_00101011_1;
      patterns[63032] = 25'b11110110_00110110_00101100_1;
      patterns[63033] = 25'b11110110_00110111_00101101_1;
      patterns[63034] = 25'b11110110_00111000_00101110_1;
      patterns[63035] = 25'b11110110_00111001_00101111_1;
      patterns[63036] = 25'b11110110_00111010_00110000_1;
      patterns[63037] = 25'b11110110_00111011_00110001_1;
      patterns[63038] = 25'b11110110_00111100_00110010_1;
      patterns[63039] = 25'b11110110_00111101_00110011_1;
      patterns[63040] = 25'b11110110_00111110_00110100_1;
      patterns[63041] = 25'b11110110_00111111_00110101_1;
      patterns[63042] = 25'b11110110_01000000_00110110_1;
      patterns[63043] = 25'b11110110_01000001_00110111_1;
      patterns[63044] = 25'b11110110_01000010_00111000_1;
      patterns[63045] = 25'b11110110_01000011_00111001_1;
      patterns[63046] = 25'b11110110_01000100_00111010_1;
      patterns[63047] = 25'b11110110_01000101_00111011_1;
      patterns[63048] = 25'b11110110_01000110_00111100_1;
      patterns[63049] = 25'b11110110_01000111_00111101_1;
      patterns[63050] = 25'b11110110_01001000_00111110_1;
      patterns[63051] = 25'b11110110_01001001_00111111_1;
      patterns[63052] = 25'b11110110_01001010_01000000_1;
      patterns[63053] = 25'b11110110_01001011_01000001_1;
      patterns[63054] = 25'b11110110_01001100_01000010_1;
      patterns[63055] = 25'b11110110_01001101_01000011_1;
      patterns[63056] = 25'b11110110_01001110_01000100_1;
      patterns[63057] = 25'b11110110_01001111_01000101_1;
      patterns[63058] = 25'b11110110_01010000_01000110_1;
      patterns[63059] = 25'b11110110_01010001_01000111_1;
      patterns[63060] = 25'b11110110_01010010_01001000_1;
      patterns[63061] = 25'b11110110_01010011_01001001_1;
      patterns[63062] = 25'b11110110_01010100_01001010_1;
      patterns[63063] = 25'b11110110_01010101_01001011_1;
      patterns[63064] = 25'b11110110_01010110_01001100_1;
      patterns[63065] = 25'b11110110_01010111_01001101_1;
      patterns[63066] = 25'b11110110_01011000_01001110_1;
      patterns[63067] = 25'b11110110_01011001_01001111_1;
      patterns[63068] = 25'b11110110_01011010_01010000_1;
      patterns[63069] = 25'b11110110_01011011_01010001_1;
      patterns[63070] = 25'b11110110_01011100_01010010_1;
      patterns[63071] = 25'b11110110_01011101_01010011_1;
      patterns[63072] = 25'b11110110_01011110_01010100_1;
      patterns[63073] = 25'b11110110_01011111_01010101_1;
      patterns[63074] = 25'b11110110_01100000_01010110_1;
      patterns[63075] = 25'b11110110_01100001_01010111_1;
      patterns[63076] = 25'b11110110_01100010_01011000_1;
      patterns[63077] = 25'b11110110_01100011_01011001_1;
      patterns[63078] = 25'b11110110_01100100_01011010_1;
      patterns[63079] = 25'b11110110_01100101_01011011_1;
      patterns[63080] = 25'b11110110_01100110_01011100_1;
      patterns[63081] = 25'b11110110_01100111_01011101_1;
      patterns[63082] = 25'b11110110_01101000_01011110_1;
      patterns[63083] = 25'b11110110_01101001_01011111_1;
      patterns[63084] = 25'b11110110_01101010_01100000_1;
      patterns[63085] = 25'b11110110_01101011_01100001_1;
      patterns[63086] = 25'b11110110_01101100_01100010_1;
      patterns[63087] = 25'b11110110_01101101_01100011_1;
      patterns[63088] = 25'b11110110_01101110_01100100_1;
      patterns[63089] = 25'b11110110_01101111_01100101_1;
      patterns[63090] = 25'b11110110_01110000_01100110_1;
      patterns[63091] = 25'b11110110_01110001_01100111_1;
      patterns[63092] = 25'b11110110_01110010_01101000_1;
      patterns[63093] = 25'b11110110_01110011_01101001_1;
      patterns[63094] = 25'b11110110_01110100_01101010_1;
      patterns[63095] = 25'b11110110_01110101_01101011_1;
      patterns[63096] = 25'b11110110_01110110_01101100_1;
      patterns[63097] = 25'b11110110_01110111_01101101_1;
      patterns[63098] = 25'b11110110_01111000_01101110_1;
      patterns[63099] = 25'b11110110_01111001_01101111_1;
      patterns[63100] = 25'b11110110_01111010_01110000_1;
      patterns[63101] = 25'b11110110_01111011_01110001_1;
      patterns[63102] = 25'b11110110_01111100_01110010_1;
      patterns[63103] = 25'b11110110_01111101_01110011_1;
      patterns[63104] = 25'b11110110_01111110_01110100_1;
      patterns[63105] = 25'b11110110_01111111_01110101_1;
      patterns[63106] = 25'b11110110_10000000_01110110_1;
      patterns[63107] = 25'b11110110_10000001_01110111_1;
      patterns[63108] = 25'b11110110_10000010_01111000_1;
      patterns[63109] = 25'b11110110_10000011_01111001_1;
      patterns[63110] = 25'b11110110_10000100_01111010_1;
      patterns[63111] = 25'b11110110_10000101_01111011_1;
      patterns[63112] = 25'b11110110_10000110_01111100_1;
      patterns[63113] = 25'b11110110_10000111_01111101_1;
      patterns[63114] = 25'b11110110_10001000_01111110_1;
      patterns[63115] = 25'b11110110_10001001_01111111_1;
      patterns[63116] = 25'b11110110_10001010_10000000_1;
      patterns[63117] = 25'b11110110_10001011_10000001_1;
      patterns[63118] = 25'b11110110_10001100_10000010_1;
      patterns[63119] = 25'b11110110_10001101_10000011_1;
      patterns[63120] = 25'b11110110_10001110_10000100_1;
      patterns[63121] = 25'b11110110_10001111_10000101_1;
      patterns[63122] = 25'b11110110_10010000_10000110_1;
      patterns[63123] = 25'b11110110_10010001_10000111_1;
      patterns[63124] = 25'b11110110_10010010_10001000_1;
      patterns[63125] = 25'b11110110_10010011_10001001_1;
      patterns[63126] = 25'b11110110_10010100_10001010_1;
      patterns[63127] = 25'b11110110_10010101_10001011_1;
      patterns[63128] = 25'b11110110_10010110_10001100_1;
      patterns[63129] = 25'b11110110_10010111_10001101_1;
      patterns[63130] = 25'b11110110_10011000_10001110_1;
      patterns[63131] = 25'b11110110_10011001_10001111_1;
      patterns[63132] = 25'b11110110_10011010_10010000_1;
      patterns[63133] = 25'b11110110_10011011_10010001_1;
      patterns[63134] = 25'b11110110_10011100_10010010_1;
      patterns[63135] = 25'b11110110_10011101_10010011_1;
      patterns[63136] = 25'b11110110_10011110_10010100_1;
      patterns[63137] = 25'b11110110_10011111_10010101_1;
      patterns[63138] = 25'b11110110_10100000_10010110_1;
      patterns[63139] = 25'b11110110_10100001_10010111_1;
      patterns[63140] = 25'b11110110_10100010_10011000_1;
      patterns[63141] = 25'b11110110_10100011_10011001_1;
      patterns[63142] = 25'b11110110_10100100_10011010_1;
      patterns[63143] = 25'b11110110_10100101_10011011_1;
      patterns[63144] = 25'b11110110_10100110_10011100_1;
      patterns[63145] = 25'b11110110_10100111_10011101_1;
      patterns[63146] = 25'b11110110_10101000_10011110_1;
      patterns[63147] = 25'b11110110_10101001_10011111_1;
      patterns[63148] = 25'b11110110_10101010_10100000_1;
      patterns[63149] = 25'b11110110_10101011_10100001_1;
      patterns[63150] = 25'b11110110_10101100_10100010_1;
      patterns[63151] = 25'b11110110_10101101_10100011_1;
      patterns[63152] = 25'b11110110_10101110_10100100_1;
      patterns[63153] = 25'b11110110_10101111_10100101_1;
      patterns[63154] = 25'b11110110_10110000_10100110_1;
      patterns[63155] = 25'b11110110_10110001_10100111_1;
      patterns[63156] = 25'b11110110_10110010_10101000_1;
      patterns[63157] = 25'b11110110_10110011_10101001_1;
      patterns[63158] = 25'b11110110_10110100_10101010_1;
      patterns[63159] = 25'b11110110_10110101_10101011_1;
      patterns[63160] = 25'b11110110_10110110_10101100_1;
      patterns[63161] = 25'b11110110_10110111_10101101_1;
      patterns[63162] = 25'b11110110_10111000_10101110_1;
      patterns[63163] = 25'b11110110_10111001_10101111_1;
      patterns[63164] = 25'b11110110_10111010_10110000_1;
      patterns[63165] = 25'b11110110_10111011_10110001_1;
      patterns[63166] = 25'b11110110_10111100_10110010_1;
      patterns[63167] = 25'b11110110_10111101_10110011_1;
      patterns[63168] = 25'b11110110_10111110_10110100_1;
      patterns[63169] = 25'b11110110_10111111_10110101_1;
      patterns[63170] = 25'b11110110_11000000_10110110_1;
      patterns[63171] = 25'b11110110_11000001_10110111_1;
      patterns[63172] = 25'b11110110_11000010_10111000_1;
      patterns[63173] = 25'b11110110_11000011_10111001_1;
      patterns[63174] = 25'b11110110_11000100_10111010_1;
      patterns[63175] = 25'b11110110_11000101_10111011_1;
      patterns[63176] = 25'b11110110_11000110_10111100_1;
      patterns[63177] = 25'b11110110_11000111_10111101_1;
      patterns[63178] = 25'b11110110_11001000_10111110_1;
      patterns[63179] = 25'b11110110_11001001_10111111_1;
      patterns[63180] = 25'b11110110_11001010_11000000_1;
      patterns[63181] = 25'b11110110_11001011_11000001_1;
      patterns[63182] = 25'b11110110_11001100_11000010_1;
      patterns[63183] = 25'b11110110_11001101_11000011_1;
      patterns[63184] = 25'b11110110_11001110_11000100_1;
      patterns[63185] = 25'b11110110_11001111_11000101_1;
      patterns[63186] = 25'b11110110_11010000_11000110_1;
      patterns[63187] = 25'b11110110_11010001_11000111_1;
      patterns[63188] = 25'b11110110_11010010_11001000_1;
      patterns[63189] = 25'b11110110_11010011_11001001_1;
      patterns[63190] = 25'b11110110_11010100_11001010_1;
      patterns[63191] = 25'b11110110_11010101_11001011_1;
      patterns[63192] = 25'b11110110_11010110_11001100_1;
      patterns[63193] = 25'b11110110_11010111_11001101_1;
      patterns[63194] = 25'b11110110_11011000_11001110_1;
      patterns[63195] = 25'b11110110_11011001_11001111_1;
      patterns[63196] = 25'b11110110_11011010_11010000_1;
      patterns[63197] = 25'b11110110_11011011_11010001_1;
      patterns[63198] = 25'b11110110_11011100_11010010_1;
      patterns[63199] = 25'b11110110_11011101_11010011_1;
      patterns[63200] = 25'b11110110_11011110_11010100_1;
      patterns[63201] = 25'b11110110_11011111_11010101_1;
      patterns[63202] = 25'b11110110_11100000_11010110_1;
      patterns[63203] = 25'b11110110_11100001_11010111_1;
      patterns[63204] = 25'b11110110_11100010_11011000_1;
      patterns[63205] = 25'b11110110_11100011_11011001_1;
      patterns[63206] = 25'b11110110_11100100_11011010_1;
      patterns[63207] = 25'b11110110_11100101_11011011_1;
      patterns[63208] = 25'b11110110_11100110_11011100_1;
      patterns[63209] = 25'b11110110_11100111_11011101_1;
      patterns[63210] = 25'b11110110_11101000_11011110_1;
      patterns[63211] = 25'b11110110_11101001_11011111_1;
      patterns[63212] = 25'b11110110_11101010_11100000_1;
      patterns[63213] = 25'b11110110_11101011_11100001_1;
      patterns[63214] = 25'b11110110_11101100_11100010_1;
      patterns[63215] = 25'b11110110_11101101_11100011_1;
      patterns[63216] = 25'b11110110_11101110_11100100_1;
      patterns[63217] = 25'b11110110_11101111_11100101_1;
      patterns[63218] = 25'b11110110_11110000_11100110_1;
      patterns[63219] = 25'b11110110_11110001_11100111_1;
      patterns[63220] = 25'b11110110_11110010_11101000_1;
      patterns[63221] = 25'b11110110_11110011_11101001_1;
      patterns[63222] = 25'b11110110_11110100_11101010_1;
      patterns[63223] = 25'b11110110_11110101_11101011_1;
      patterns[63224] = 25'b11110110_11110110_11101100_1;
      patterns[63225] = 25'b11110110_11110111_11101101_1;
      patterns[63226] = 25'b11110110_11111000_11101110_1;
      patterns[63227] = 25'b11110110_11111001_11101111_1;
      patterns[63228] = 25'b11110110_11111010_11110000_1;
      patterns[63229] = 25'b11110110_11111011_11110001_1;
      patterns[63230] = 25'b11110110_11111100_11110010_1;
      patterns[63231] = 25'b11110110_11111101_11110011_1;
      patterns[63232] = 25'b11110110_11111110_11110100_1;
      patterns[63233] = 25'b11110110_11111111_11110101_1;
      patterns[63234] = 25'b11110111_00000000_11110111_0;
      patterns[63235] = 25'b11110111_00000001_11111000_0;
      patterns[63236] = 25'b11110111_00000010_11111001_0;
      patterns[63237] = 25'b11110111_00000011_11111010_0;
      patterns[63238] = 25'b11110111_00000100_11111011_0;
      patterns[63239] = 25'b11110111_00000101_11111100_0;
      patterns[63240] = 25'b11110111_00000110_11111101_0;
      patterns[63241] = 25'b11110111_00000111_11111110_0;
      patterns[63242] = 25'b11110111_00001000_11111111_0;
      patterns[63243] = 25'b11110111_00001001_00000000_1;
      patterns[63244] = 25'b11110111_00001010_00000001_1;
      patterns[63245] = 25'b11110111_00001011_00000010_1;
      patterns[63246] = 25'b11110111_00001100_00000011_1;
      patterns[63247] = 25'b11110111_00001101_00000100_1;
      patterns[63248] = 25'b11110111_00001110_00000101_1;
      patterns[63249] = 25'b11110111_00001111_00000110_1;
      patterns[63250] = 25'b11110111_00010000_00000111_1;
      patterns[63251] = 25'b11110111_00010001_00001000_1;
      patterns[63252] = 25'b11110111_00010010_00001001_1;
      patterns[63253] = 25'b11110111_00010011_00001010_1;
      patterns[63254] = 25'b11110111_00010100_00001011_1;
      patterns[63255] = 25'b11110111_00010101_00001100_1;
      patterns[63256] = 25'b11110111_00010110_00001101_1;
      patterns[63257] = 25'b11110111_00010111_00001110_1;
      patterns[63258] = 25'b11110111_00011000_00001111_1;
      patterns[63259] = 25'b11110111_00011001_00010000_1;
      patterns[63260] = 25'b11110111_00011010_00010001_1;
      patterns[63261] = 25'b11110111_00011011_00010010_1;
      patterns[63262] = 25'b11110111_00011100_00010011_1;
      patterns[63263] = 25'b11110111_00011101_00010100_1;
      patterns[63264] = 25'b11110111_00011110_00010101_1;
      patterns[63265] = 25'b11110111_00011111_00010110_1;
      patterns[63266] = 25'b11110111_00100000_00010111_1;
      patterns[63267] = 25'b11110111_00100001_00011000_1;
      patterns[63268] = 25'b11110111_00100010_00011001_1;
      patterns[63269] = 25'b11110111_00100011_00011010_1;
      patterns[63270] = 25'b11110111_00100100_00011011_1;
      patterns[63271] = 25'b11110111_00100101_00011100_1;
      patterns[63272] = 25'b11110111_00100110_00011101_1;
      patterns[63273] = 25'b11110111_00100111_00011110_1;
      patterns[63274] = 25'b11110111_00101000_00011111_1;
      patterns[63275] = 25'b11110111_00101001_00100000_1;
      patterns[63276] = 25'b11110111_00101010_00100001_1;
      patterns[63277] = 25'b11110111_00101011_00100010_1;
      patterns[63278] = 25'b11110111_00101100_00100011_1;
      patterns[63279] = 25'b11110111_00101101_00100100_1;
      patterns[63280] = 25'b11110111_00101110_00100101_1;
      patterns[63281] = 25'b11110111_00101111_00100110_1;
      patterns[63282] = 25'b11110111_00110000_00100111_1;
      patterns[63283] = 25'b11110111_00110001_00101000_1;
      patterns[63284] = 25'b11110111_00110010_00101001_1;
      patterns[63285] = 25'b11110111_00110011_00101010_1;
      patterns[63286] = 25'b11110111_00110100_00101011_1;
      patterns[63287] = 25'b11110111_00110101_00101100_1;
      patterns[63288] = 25'b11110111_00110110_00101101_1;
      patterns[63289] = 25'b11110111_00110111_00101110_1;
      patterns[63290] = 25'b11110111_00111000_00101111_1;
      patterns[63291] = 25'b11110111_00111001_00110000_1;
      patterns[63292] = 25'b11110111_00111010_00110001_1;
      patterns[63293] = 25'b11110111_00111011_00110010_1;
      patterns[63294] = 25'b11110111_00111100_00110011_1;
      patterns[63295] = 25'b11110111_00111101_00110100_1;
      patterns[63296] = 25'b11110111_00111110_00110101_1;
      patterns[63297] = 25'b11110111_00111111_00110110_1;
      patterns[63298] = 25'b11110111_01000000_00110111_1;
      patterns[63299] = 25'b11110111_01000001_00111000_1;
      patterns[63300] = 25'b11110111_01000010_00111001_1;
      patterns[63301] = 25'b11110111_01000011_00111010_1;
      patterns[63302] = 25'b11110111_01000100_00111011_1;
      patterns[63303] = 25'b11110111_01000101_00111100_1;
      patterns[63304] = 25'b11110111_01000110_00111101_1;
      patterns[63305] = 25'b11110111_01000111_00111110_1;
      patterns[63306] = 25'b11110111_01001000_00111111_1;
      patterns[63307] = 25'b11110111_01001001_01000000_1;
      patterns[63308] = 25'b11110111_01001010_01000001_1;
      patterns[63309] = 25'b11110111_01001011_01000010_1;
      patterns[63310] = 25'b11110111_01001100_01000011_1;
      patterns[63311] = 25'b11110111_01001101_01000100_1;
      patterns[63312] = 25'b11110111_01001110_01000101_1;
      patterns[63313] = 25'b11110111_01001111_01000110_1;
      patterns[63314] = 25'b11110111_01010000_01000111_1;
      patterns[63315] = 25'b11110111_01010001_01001000_1;
      patterns[63316] = 25'b11110111_01010010_01001001_1;
      patterns[63317] = 25'b11110111_01010011_01001010_1;
      patterns[63318] = 25'b11110111_01010100_01001011_1;
      patterns[63319] = 25'b11110111_01010101_01001100_1;
      patterns[63320] = 25'b11110111_01010110_01001101_1;
      patterns[63321] = 25'b11110111_01010111_01001110_1;
      patterns[63322] = 25'b11110111_01011000_01001111_1;
      patterns[63323] = 25'b11110111_01011001_01010000_1;
      patterns[63324] = 25'b11110111_01011010_01010001_1;
      patterns[63325] = 25'b11110111_01011011_01010010_1;
      patterns[63326] = 25'b11110111_01011100_01010011_1;
      patterns[63327] = 25'b11110111_01011101_01010100_1;
      patterns[63328] = 25'b11110111_01011110_01010101_1;
      patterns[63329] = 25'b11110111_01011111_01010110_1;
      patterns[63330] = 25'b11110111_01100000_01010111_1;
      patterns[63331] = 25'b11110111_01100001_01011000_1;
      patterns[63332] = 25'b11110111_01100010_01011001_1;
      patterns[63333] = 25'b11110111_01100011_01011010_1;
      patterns[63334] = 25'b11110111_01100100_01011011_1;
      patterns[63335] = 25'b11110111_01100101_01011100_1;
      patterns[63336] = 25'b11110111_01100110_01011101_1;
      patterns[63337] = 25'b11110111_01100111_01011110_1;
      patterns[63338] = 25'b11110111_01101000_01011111_1;
      patterns[63339] = 25'b11110111_01101001_01100000_1;
      patterns[63340] = 25'b11110111_01101010_01100001_1;
      patterns[63341] = 25'b11110111_01101011_01100010_1;
      patterns[63342] = 25'b11110111_01101100_01100011_1;
      patterns[63343] = 25'b11110111_01101101_01100100_1;
      patterns[63344] = 25'b11110111_01101110_01100101_1;
      patterns[63345] = 25'b11110111_01101111_01100110_1;
      patterns[63346] = 25'b11110111_01110000_01100111_1;
      patterns[63347] = 25'b11110111_01110001_01101000_1;
      patterns[63348] = 25'b11110111_01110010_01101001_1;
      patterns[63349] = 25'b11110111_01110011_01101010_1;
      patterns[63350] = 25'b11110111_01110100_01101011_1;
      patterns[63351] = 25'b11110111_01110101_01101100_1;
      patterns[63352] = 25'b11110111_01110110_01101101_1;
      patterns[63353] = 25'b11110111_01110111_01101110_1;
      patterns[63354] = 25'b11110111_01111000_01101111_1;
      patterns[63355] = 25'b11110111_01111001_01110000_1;
      patterns[63356] = 25'b11110111_01111010_01110001_1;
      patterns[63357] = 25'b11110111_01111011_01110010_1;
      patterns[63358] = 25'b11110111_01111100_01110011_1;
      patterns[63359] = 25'b11110111_01111101_01110100_1;
      patterns[63360] = 25'b11110111_01111110_01110101_1;
      patterns[63361] = 25'b11110111_01111111_01110110_1;
      patterns[63362] = 25'b11110111_10000000_01110111_1;
      patterns[63363] = 25'b11110111_10000001_01111000_1;
      patterns[63364] = 25'b11110111_10000010_01111001_1;
      patterns[63365] = 25'b11110111_10000011_01111010_1;
      patterns[63366] = 25'b11110111_10000100_01111011_1;
      patterns[63367] = 25'b11110111_10000101_01111100_1;
      patterns[63368] = 25'b11110111_10000110_01111101_1;
      patterns[63369] = 25'b11110111_10000111_01111110_1;
      patterns[63370] = 25'b11110111_10001000_01111111_1;
      patterns[63371] = 25'b11110111_10001001_10000000_1;
      patterns[63372] = 25'b11110111_10001010_10000001_1;
      patterns[63373] = 25'b11110111_10001011_10000010_1;
      patterns[63374] = 25'b11110111_10001100_10000011_1;
      patterns[63375] = 25'b11110111_10001101_10000100_1;
      patterns[63376] = 25'b11110111_10001110_10000101_1;
      patterns[63377] = 25'b11110111_10001111_10000110_1;
      patterns[63378] = 25'b11110111_10010000_10000111_1;
      patterns[63379] = 25'b11110111_10010001_10001000_1;
      patterns[63380] = 25'b11110111_10010010_10001001_1;
      patterns[63381] = 25'b11110111_10010011_10001010_1;
      patterns[63382] = 25'b11110111_10010100_10001011_1;
      patterns[63383] = 25'b11110111_10010101_10001100_1;
      patterns[63384] = 25'b11110111_10010110_10001101_1;
      patterns[63385] = 25'b11110111_10010111_10001110_1;
      patterns[63386] = 25'b11110111_10011000_10001111_1;
      patterns[63387] = 25'b11110111_10011001_10010000_1;
      patterns[63388] = 25'b11110111_10011010_10010001_1;
      patterns[63389] = 25'b11110111_10011011_10010010_1;
      patterns[63390] = 25'b11110111_10011100_10010011_1;
      patterns[63391] = 25'b11110111_10011101_10010100_1;
      patterns[63392] = 25'b11110111_10011110_10010101_1;
      patterns[63393] = 25'b11110111_10011111_10010110_1;
      patterns[63394] = 25'b11110111_10100000_10010111_1;
      patterns[63395] = 25'b11110111_10100001_10011000_1;
      patterns[63396] = 25'b11110111_10100010_10011001_1;
      patterns[63397] = 25'b11110111_10100011_10011010_1;
      patterns[63398] = 25'b11110111_10100100_10011011_1;
      patterns[63399] = 25'b11110111_10100101_10011100_1;
      patterns[63400] = 25'b11110111_10100110_10011101_1;
      patterns[63401] = 25'b11110111_10100111_10011110_1;
      patterns[63402] = 25'b11110111_10101000_10011111_1;
      patterns[63403] = 25'b11110111_10101001_10100000_1;
      patterns[63404] = 25'b11110111_10101010_10100001_1;
      patterns[63405] = 25'b11110111_10101011_10100010_1;
      patterns[63406] = 25'b11110111_10101100_10100011_1;
      patterns[63407] = 25'b11110111_10101101_10100100_1;
      patterns[63408] = 25'b11110111_10101110_10100101_1;
      patterns[63409] = 25'b11110111_10101111_10100110_1;
      patterns[63410] = 25'b11110111_10110000_10100111_1;
      patterns[63411] = 25'b11110111_10110001_10101000_1;
      patterns[63412] = 25'b11110111_10110010_10101001_1;
      patterns[63413] = 25'b11110111_10110011_10101010_1;
      patterns[63414] = 25'b11110111_10110100_10101011_1;
      patterns[63415] = 25'b11110111_10110101_10101100_1;
      patterns[63416] = 25'b11110111_10110110_10101101_1;
      patterns[63417] = 25'b11110111_10110111_10101110_1;
      patterns[63418] = 25'b11110111_10111000_10101111_1;
      patterns[63419] = 25'b11110111_10111001_10110000_1;
      patterns[63420] = 25'b11110111_10111010_10110001_1;
      patterns[63421] = 25'b11110111_10111011_10110010_1;
      patterns[63422] = 25'b11110111_10111100_10110011_1;
      patterns[63423] = 25'b11110111_10111101_10110100_1;
      patterns[63424] = 25'b11110111_10111110_10110101_1;
      patterns[63425] = 25'b11110111_10111111_10110110_1;
      patterns[63426] = 25'b11110111_11000000_10110111_1;
      patterns[63427] = 25'b11110111_11000001_10111000_1;
      patterns[63428] = 25'b11110111_11000010_10111001_1;
      patterns[63429] = 25'b11110111_11000011_10111010_1;
      patterns[63430] = 25'b11110111_11000100_10111011_1;
      patterns[63431] = 25'b11110111_11000101_10111100_1;
      patterns[63432] = 25'b11110111_11000110_10111101_1;
      patterns[63433] = 25'b11110111_11000111_10111110_1;
      patterns[63434] = 25'b11110111_11001000_10111111_1;
      patterns[63435] = 25'b11110111_11001001_11000000_1;
      patterns[63436] = 25'b11110111_11001010_11000001_1;
      patterns[63437] = 25'b11110111_11001011_11000010_1;
      patterns[63438] = 25'b11110111_11001100_11000011_1;
      patterns[63439] = 25'b11110111_11001101_11000100_1;
      patterns[63440] = 25'b11110111_11001110_11000101_1;
      patterns[63441] = 25'b11110111_11001111_11000110_1;
      patterns[63442] = 25'b11110111_11010000_11000111_1;
      patterns[63443] = 25'b11110111_11010001_11001000_1;
      patterns[63444] = 25'b11110111_11010010_11001001_1;
      patterns[63445] = 25'b11110111_11010011_11001010_1;
      patterns[63446] = 25'b11110111_11010100_11001011_1;
      patterns[63447] = 25'b11110111_11010101_11001100_1;
      patterns[63448] = 25'b11110111_11010110_11001101_1;
      patterns[63449] = 25'b11110111_11010111_11001110_1;
      patterns[63450] = 25'b11110111_11011000_11001111_1;
      patterns[63451] = 25'b11110111_11011001_11010000_1;
      patterns[63452] = 25'b11110111_11011010_11010001_1;
      patterns[63453] = 25'b11110111_11011011_11010010_1;
      patterns[63454] = 25'b11110111_11011100_11010011_1;
      patterns[63455] = 25'b11110111_11011101_11010100_1;
      patterns[63456] = 25'b11110111_11011110_11010101_1;
      patterns[63457] = 25'b11110111_11011111_11010110_1;
      patterns[63458] = 25'b11110111_11100000_11010111_1;
      patterns[63459] = 25'b11110111_11100001_11011000_1;
      patterns[63460] = 25'b11110111_11100010_11011001_1;
      patterns[63461] = 25'b11110111_11100011_11011010_1;
      patterns[63462] = 25'b11110111_11100100_11011011_1;
      patterns[63463] = 25'b11110111_11100101_11011100_1;
      patterns[63464] = 25'b11110111_11100110_11011101_1;
      patterns[63465] = 25'b11110111_11100111_11011110_1;
      patterns[63466] = 25'b11110111_11101000_11011111_1;
      patterns[63467] = 25'b11110111_11101001_11100000_1;
      patterns[63468] = 25'b11110111_11101010_11100001_1;
      patterns[63469] = 25'b11110111_11101011_11100010_1;
      patterns[63470] = 25'b11110111_11101100_11100011_1;
      patterns[63471] = 25'b11110111_11101101_11100100_1;
      patterns[63472] = 25'b11110111_11101110_11100101_1;
      patterns[63473] = 25'b11110111_11101111_11100110_1;
      patterns[63474] = 25'b11110111_11110000_11100111_1;
      patterns[63475] = 25'b11110111_11110001_11101000_1;
      patterns[63476] = 25'b11110111_11110010_11101001_1;
      patterns[63477] = 25'b11110111_11110011_11101010_1;
      patterns[63478] = 25'b11110111_11110100_11101011_1;
      patterns[63479] = 25'b11110111_11110101_11101100_1;
      patterns[63480] = 25'b11110111_11110110_11101101_1;
      patterns[63481] = 25'b11110111_11110111_11101110_1;
      patterns[63482] = 25'b11110111_11111000_11101111_1;
      patterns[63483] = 25'b11110111_11111001_11110000_1;
      patterns[63484] = 25'b11110111_11111010_11110001_1;
      patterns[63485] = 25'b11110111_11111011_11110010_1;
      patterns[63486] = 25'b11110111_11111100_11110011_1;
      patterns[63487] = 25'b11110111_11111101_11110100_1;
      patterns[63488] = 25'b11110111_11111110_11110101_1;
      patterns[63489] = 25'b11110111_11111111_11110110_1;
      patterns[63490] = 25'b11111000_00000000_11111000_0;
      patterns[63491] = 25'b11111000_00000001_11111001_0;
      patterns[63492] = 25'b11111000_00000010_11111010_0;
      patterns[63493] = 25'b11111000_00000011_11111011_0;
      patterns[63494] = 25'b11111000_00000100_11111100_0;
      patterns[63495] = 25'b11111000_00000101_11111101_0;
      patterns[63496] = 25'b11111000_00000110_11111110_0;
      patterns[63497] = 25'b11111000_00000111_11111111_0;
      patterns[63498] = 25'b11111000_00001000_00000000_1;
      patterns[63499] = 25'b11111000_00001001_00000001_1;
      patterns[63500] = 25'b11111000_00001010_00000010_1;
      patterns[63501] = 25'b11111000_00001011_00000011_1;
      patterns[63502] = 25'b11111000_00001100_00000100_1;
      patterns[63503] = 25'b11111000_00001101_00000101_1;
      patterns[63504] = 25'b11111000_00001110_00000110_1;
      patterns[63505] = 25'b11111000_00001111_00000111_1;
      patterns[63506] = 25'b11111000_00010000_00001000_1;
      patterns[63507] = 25'b11111000_00010001_00001001_1;
      patterns[63508] = 25'b11111000_00010010_00001010_1;
      patterns[63509] = 25'b11111000_00010011_00001011_1;
      patterns[63510] = 25'b11111000_00010100_00001100_1;
      patterns[63511] = 25'b11111000_00010101_00001101_1;
      patterns[63512] = 25'b11111000_00010110_00001110_1;
      patterns[63513] = 25'b11111000_00010111_00001111_1;
      patterns[63514] = 25'b11111000_00011000_00010000_1;
      patterns[63515] = 25'b11111000_00011001_00010001_1;
      patterns[63516] = 25'b11111000_00011010_00010010_1;
      patterns[63517] = 25'b11111000_00011011_00010011_1;
      patterns[63518] = 25'b11111000_00011100_00010100_1;
      patterns[63519] = 25'b11111000_00011101_00010101_1;
      patterns[63520] = 25'b11111000_00011110_00010110_1;
      patterns[63521] = 25'b11111000_00011111_00010111_1;
      patterns[63522] = 25'b11111000_00100000_00011000_1;
      patterns[63523] = 25'b11111000_00100001_00011001_1;
      patterns[63524] = 25'b11111000_00100010_00011010_1;
      patterns[63525] = 25'b11111000_00100011_00011011_1;
      patterns[63526] = 25'b11111000_00100100_00011100_1;
      patterns[63527] = 25'b11111000_00100101_00011101_1;
      patterns[63528] = 25'b11111000_00100110_00011110_1;
      patterns[63529] = 25'b11111000_00100111_00011111_1;
      patterns[63530] = 25'b11111000_00101000_00100000_1;
      patterns[63531] = 25'b11111000_00101001_00100001_1;
      patterns[63532] = 25'b11111000_00101010_00100010_1;
      patterns[63533] = 25'b11111000_00101011_00100011_1;
      patterns[63534] = 25'b11111000_00101100_00100100_1;
      patterns[63535] = 25'b11111000_00101101_00100101_1;
      patterns[63536] = 25'b11111000_00101110_00100110_1;
      patterns[63537] = 25'b11111000_00101111_00100111_1;
      patterns[63538] = 25'b11111000_00110000_00101000_1;
      patterns[63539] = 25'b11111000_00110001_00101001_1;
      patterns[63540] = 25'b11111000_00110010_00101010_1;
      patterns[63541] = 25'b11111000_00110011_00101011_1;
      patterns[63542] = 25'b11111000_00110100_00101100_1;
      patterns[63543] = 25'b11111000_00110101_00101101_1;
      patterns[63544] = 25'b11111000_00110110_00101110_1;
      patterns[63545] = 25'b11111000_00110111_00101111_1;
      patterns[63546] = 25'b11111000_00111000_00110000_1;
      patterns[63547] = 25'b11111000_00111001_00110001_1;
      patterns[63548] = 25'b11111000_00111010_00110010_1;
      patterns[63549] = 25'b11111000_00111011_00110011_1;
      patterns[63550] = 25'b11111000_00111100_00110100_1;
      patterns[63551] = 25'b11111000_00111101_00110101_1;
      patterns[63552] = 25'b11111000_00111110_00110110_1;
      patterns[63553] = 25'b11111000_00111111_00110111_1;
      patterns[63554] = 25'b11111000_01000000_00111000_1;
      patterns[63555] = 25'b11111000_01000001_00111001_1;
      patterns[63556] = 25'b11111000_01000010_00111010_1;
      patterns[63557] = 25'b11111000_01000011_00111011_1;
      patterns[63558] = 25'b11111000_01000100_00111100_1;
      patterns[63559] = 25'b11111000_01000101_00111101_1;
      patterns[63560] = 25'b11111000_01000110_00111110_1;
      patterns[63561] = 25'b11111000_01000111_00111111_1;
      patterns[63562] = 25'b11111000_01001000_01000000_1;
      patterns[63563] = 25'b11111000_01001001_01000001_1;
      patterns[63564] = 25'b11111000_01001010_01000010_1;
      patterns[63565] = 25'b11111000_01001011_01000011_1;
      patterns[63566] = 25'b11111000_01001100_01000100_1;
      patterns[63567] = 25'b11111000_01001101_01000101_1;
      patterns[63568] = 25'b11111000_01001110_01000110_1;
      patterns[63569] = 25'b11111000_01001111_01000111_1;
      patterns[63570] = 25'b11111000_01010000_01001000_1;
      patterns[63571] = 25'b11111000_01010001_01001001_1;
      patterns[63572] = 25'b11111000_01010010_01001010_1;
      patterns[63573] = 25'b11111000_01010011_01001011_1;
      patterns[63574] = 25'b11111000_01010100_01001100_1;
      patterns[63575] = 25'b11111000_01010101_01001101_1;
      patterns[63576] = 25'b11111000_01010110_01001110_1;
      patterns[63577] = 25'b11111000_01010111_01001111_1;
      patterns[63578] = 25'b11111000_01011000_01010000_1;
      patterns[63579] = 25'b11111000_01011001_01010001_1;
      patterns[63580] = 25'b11111000_01011010_01010010_1;
      patterns[63581] = 25'b11111000_01011011_01010011_1;
      patterns[63582] = 25'b11111000_01011100_01010100_1;
      patterns[63583] = 25'b11111000_01011101_01010101_1;
      patterns[63584] = 25'b11111000_01011110_01010110_1;
      patterns[63585] = 25'b11111000_01011111_01010111_1;
      patterns[63586] = 25'b11111000_01100000_01011000_1;
      patterns[63587] = 25'b11111000_01100001_01011001_1;
      patterns[63588] = 25'b11111000_01100010_01011010_1;
      patterns[63589] = 25'b11111000_01100011_01011011_1;
      patterns[63590] = 25'b11111000_01100100_01011100_1;
      patterns[63591] = 25'b11111000_01100101_01011101_1;
      patterns[63592] = 25'b11111000_01100110_01011110_1;
      patterns[63593] = 25'b11111000_01100111_01011111_1;
      patterns[63594] = 25'b11111000_01101000_01100000_1;
      patterns[63595] = 25'b11111000_01101001_01100001_1;
      patterns[63596] = 25'b11111000_01101010_01100010_1;
      patterns[63597] = 25'b11111000_01101011_01100011_1;
      patterns[63598] = 25'b11111000_01101100_01100100_1;
      patterns[63599] = 25'b11111000_01101101_01100101_1;
      patterns[63600] = 25'b11111000_01101110_01100110_1;
      patterns[63601] = 25'b11111000_01101111_01100111_1;
      patterns[63602] = 25'b11111000_01110000_01101000_1;
      patterns[63603] = 25'b11111000_01110001_01101001_1;
      patterns[63604] = 25'b11111000_01110010_01101010_1;
      patterns[63605] = 25'b11111000_01110011_01101011_1;
      patterns[63606] = 25'b11111000_01110100_01101100_1;
      patterns[63607] = 25'b11111000_01110101_01101101_1;
      patterns[63608] = 25'b11111000_01110110_01101110_1;
      patterns[63609] = 25'b11111000_01110111_01101111_1;
      patterns[63610] = 25'b11111000_01111000_01110000_1;
      patterns[63611] = 25'b11111000_01111001_01110001_1;
      patterns[63612] = 25'b11111000_01111010_01110010_1;
      patterns[63613] = 25'b11111000_01111011_01110011_1;
      patterns[63614] = 25'b11111000_01111100_01110100_1;
      patterns[63615] = 25'b11111000_01111101_01110101_1;
      patterns[63616] = 25'b11111000_01111110_01110110_1;
      patterns[63617] = 25'b11111000_01111111_01110111_1;
      patterns[63618] = 25'b11111000_10000000_01111000_1;
      patterns[63619] = 25'b11111000_10000001_01111001_1;
      patterns[63620] = 25'b11111000_10000010_01111010_1;
      patterns[63621] = 25'b11111000_10000011_01111011_1;
      patterns[63622] = 25'b11111000_10000100_01111100_1;
      patterns[63623] = 25'b11111000_10000101_01111101_1;
      patterns[63624] = 25'b11111000_10000110_01111110_1;
      patterns[63625] = 25'b11111000_10000111_01111111_1;
      patterns[63626] = 25'b11111000_10001000_10000000_1;
      patterns[63627] = 25'b11111000_10001001_10000001_1;
      patterns[63628] = 25'b11111000_10001010_10000010_1;
      patterns[63629] = 25'b11111000_10001011_10000011_1;
      patterns[63630] = 25'b11111000_10001100_10000100_1;
      patterns[63631] = 25'b11111000_10001101_10000101_1;
      patterns[63632] = 25'b11111000_10001110_10000110_1;
      patterns[63633] = 25'b11111000_10001111_10000111_1;
      patterns[63634] = 25'b11111000_10010000_10001000_1;
      patterns[63635] = 25'b11111000_10010001_10001001_1;
      patterns[63636] = 25'b11111000_10010010_10001010_1;
      patterns[63637] = 25'b11111000_10010011_10001011_1;
      patterns[63638] = 25'b11111000_10010100_10001100_1;
      patterns[63639] = 25'b11111000_10010101_10001101_1;
      patterns[63640] = 25'b11111000_10010110_10001110_1;
      patterns[63641] = 25'b11111000_10010111_10001111_1;
      patterns[63642] = 25'b11111000_10011000_10010000_1;
      patterns[63643] = 25'b11111000_10011001_10010001_1;
      patterns[63644] = 25'b11111000_10011010_10010010_1;
      patterns[63645] = 25'b11111000_10011011_10010011_1;
      patterns[63646] = 25'b11111000_10011100_10010100_1;
      patterns[63647] = 25'b11111000_10011101_10010101_1;
      patterns[63648] = 25'b11111000_10011110_10010110_1;
      patterns[63649] = 25'b11111000_10011111_10010111_1;
      patterns[63650] = 25'b11111000_10100000_10011000_1;
      patterns[63651] = 25'b11111000_10100001_10011001_1;
      patterns[63652] = 25'b11111000_10100010_10011010_1;
      patterns[63653] = 25'b11111000_10100011_10011011_1;
      patterns[63654] = 25'b11111000_10100100_10011100_1;
      patterns[63655] = 25'b11111000_10100101_10011101_1;
      patterns[63656] = 25'b11111000_10100110_10011110_1;
      patterns[63657] = 25'b11111000_10100111_10011111_1;
      patterns[63658] = 25'b11111000_10101000_10100000_1;
      patterns[63659] = 25'b11111000_10101001_10100001_1;
      patterns[63660] = 25'b11111000_10101010_10100010_1;
      patterns[63661] = 25'b11111000_10101011_10100011_1;
      patterns[63662] = 25'b11111000_10101100_10100100_1;
      patterns[63663] = 25'b11111000_10101101_10100101_1;
      patterns[63664] = 25'b11111000_10101110_10100110_1;
      patterns[63665] = 25'b11111000_10101111_10100111_1;
      patterns[63666] = 25'b11111000_10110000_10101000_1;
      patterns[63667] = 25'b11111000_10110001_10101001_1;
      patterns[63668] = 25'b11111000_10110010_10101010_1;
      patterns[63669] = 25'b11111000_10110011_10101011_1;
      patterns[63670] = 25'b11111000_10110100_10101100_1;
      patterns[63671] = 25'b11111000_10110101_10101101_1;
      patterns[63672] = 25'b11111000_10110110_10101110_1;
      patterns[63673] = 25'b11111000_10110111_10101111_1;
      patterns[63674] = 25'b11111000_10111000_10110000_1;
      patterns[63675] = 25'b11111000_10111001_10110001_1;
      patterns[63676] = 25'b11111000_10111010_10110010_1;
      patterns[63677] = 25'b11111000_10111011_10110011_1;
      patterns[63678] = 25'b11111000_10111100_10110100_1;
      patterns[63679] = 25'b11111000_10111101_10110101_1;
      patterns[63680] = 25'b11111000_10111110_10110110_1;
      patterns[63681] = 25'b11111000_10111111_10110111_1;
      patterns[63682] = 25'b11111000_11000000_10111000_1;
      patterns[63683] = 25'b11111000_11000001_10111001_1;
      patterns[63684] = 25'b11111000_11000010_10111010_1;
      patterns[63685] = 25'b11111000_11000011_10111011_1;
      patterns[63686] = 25'b11111000_11000100_10111100_1;
      patterns[63687] = 25'b11111000_11000101_10111101_1;
      patterns[63688] = 25'b11111000_11000110_10111110_1;
      patterns[63689] = 25'b11111000_11000111_10111111_1;
      patterns[63690] = 25'b11111000_11001000_11000000_1;
      patterns[63691] = 25'b11111000_11001001_11000001_1;
      patterns[63692] = 25'b11111000_11001010_11000010_1;
      patterns[63693] = 25'b11111000_11001011_11000011_1;
      patterns[63694] = 25'b11111000_11001100_11000100_1;
      patterns[63695] = 25'b11111000_11001101_11000101_1;
      patterns[63696] = 25'b11111000_11001110_11000110_1;
      patterns[63697] = 25'b11111000_11001111_11000111_1;
      patterns[63698] = 25'b11111000_11010000_11001000_1;
      patterns[63699] = 25'b11111000_11010001_11001001_1;
      patterns[63700] = 25'b11111000_11010010_11001010_1;
      patterns[63701] = 25'b11111000_11010011_11001011_1;
      patterns[63702] = 25'b11111000_11010100_11001100_1;
      patterns[63703] = 25'b11111000_11010101_11001101_1;
      patterns[63704] = 25'b11111000_11010110_11001110_1;
      patterns[63705] = 25'b11111000_11010111_11001111_1;
      patterns[63706] = 25'b11111000_11011000_11010000_1;
      patterns[63707] = 25'b11111000_11011001_11010001_1;
      patterns[63708] = 25'b11111000_11011010_11010010_1;
      patterns[63709] = 25'b11111000_11011011_11010011_1;
      patterns[63710] = 25'b11111000_11011100_11010100_1;
      patterns[63711] = 25'b11111000_11011101_11010101_1;
      patterns[63712] = 25'b11111000_11011110_11010110_1;
      patterns[63713] = 25'b11111000_11011111_11010111_1;
      patterns[63714] = 25'b11111000_11100000_11011000_1;
      patterns[63715] = 25'b11111000_11100001_11011001_1;
      patterns[63716] = 25'b11111000_11100010_11011010_1;
      patterns[63717] = 25'b11111000_11100011_11011011_1;
      patterns[63718] = 25'b11111000_11100100_11011100_1;
      patterns[63719] = 25'b11111000_11100101_11011101_1;
      patterns[63720] = 25'b11111000_11100110_11011110_1;
      patterns[63721] = 25'b11111000_11100111_11011111_1;
      patterns[63722] = 25'b11111000_11101000_11100000_1;
      patterns[63723] = 25'b11111000_11101001_11100001_1;
      patterns[63724] = 25'b11111000_11101010_11100010_1;
      patterns[63725] = 25'b11111000_11101011_11100011_1;
      patterns[63726] = 25'b11111000_11101100_11100100_1;
      patterns[63727] = 25'b11111000_11101101_11100101_1;
      patterns[63728] = 25'b11111000_11101110_11100110_1;
      patterns[63729] = 25'b11111000_11101111_11100111_1;
      patterns[63730] = 25'b11111000_11110000_11101000_1;
      patterns[63731] = 25'b11111000_11110001_11101001_1;
      patterns[63732] = 25'b11111000_11110010_11101010_1;
      patterns[63733] = 25'b11111000_11110011_11101011_1;
      patterns[63734] = 25'b11111000_11110100_11101100_1;
      patterns[63735] = 25'b11111000_11110101_11101101_1;
      patterns[63736] = 25'b11111000_11110110_11101110_1;
      patterns[63737] = 25'b11111000_11110111_11101111_1;
      patterns[63738] = 25'b11111000_11111000_11110000_1;
      patterns[63739] = 25'b11111000_11111001_11110001_1;
      patterns[63740] = 25'b11111000_11111010_11110010_1;
      patterns[63741] = 25'b11111000_11111011_11110011_1;
      patterns[63742] = 25'b11111000_11111100_11110100_1;
      patterns[63743] = 25'b11111000_11111101_11110101_1;
      patterns[63744] = 25'b11111000_11111110_11110110_1;
      patterns[63745] = 25'b11111000_11111111_11110111_1;
      patterns[63746] = 25'b11111001_00000000_11111001_0;
      patterns[63747] = 25'b11111001_00000001_11111010_0;
      patterns[63748] = 25'b11111001_00000010_11111011_0;
      patterns[63749] = 25'b11111001_00000011_11111100_0;
      patterns[63750] = 25'b11111001_00000100_11111101_0;
      patterns[63751] = 25'b11111001_00000101_11111110_0;
      patterns[63752] = 25'b11111001_00000110_11111111_0;
      patterns[63753] = 25'b11111001_00000111_00000000_1;
      patterns[63754] = 25'b11111001_00001000_00000001_1;
      patterns[63755] = 25'b11111001_00001001_00000010_1;
      patterns[63756] = 25'b11111001_00001010_00000011_1;
      patterns[63757] = 25'b11111001_00001011_00000100_1;
      patterns[63758] = 25'b11111001_00001100_00000101_1;
      patterns[63759] = 25'b11111001_00001101_00000110_1;
      patterns[63760] = 25'b11111001_00001110_00000111_1;
      patterns[63761] = 25'b11111001_00001111_00001000_1;
      patterns[63762] = 25'b11111001_00010000_00001001_1;
      patterns[63763] = 25'b11111001_00010001_00001010_1;
      patterns[63764] = 25'b11111001_00010010_00001011_1;
      patterns[63765] = 25'b11111001_00010011_00001100_1;
      patterns[63766] = 25'b11111001_00010100_00001101_1;
      patterns[63767] = 25'b11111001_00010101_00001110_1;
      patterns[63768] = 25'b11111001_00010110_00001111_1;
      patterns[63769] = 25'b11111001_00010111_00010000_1;
      patterns[63770] = 25'b11111001_00011000_00010001_1;
      patterns[63771] = 25'b11111001_00011001_00010010_1;
      patterns[63772] = 25'b11111001_00011010_00010011_1;
      patterns[63773] = 25'b11111001_00011011_00010100_1;
      patterns[63774] = 25'b11111001_00011100_00010101_1;
      patterns[63775] = 25'b11111001_00011101_00010110_1;
      patterns[63776] = 25'b11111001_00011110_00010111_1;
      patterns[63777] = 25'b11111001_00011111_00011000_1;
      patterns[63778] = 25'b11111001_00100000_00011001_1;
      patterns[63779] = 25'b11111001_00100001_00011010_1;
      patterns[63780] = 25'b11111001_00100010_00011011_1;
      patterns[63781] = 25'b11111001_00100011_00011100_1;
      patterns[63782] = 25'b11111001_00100100_00011101_1;
      patterns[63783] = 25'b11111001_00100101_00011110_1;
      patterns[63784] = 25'b11111001_00100110_00011111_1;
      patterns[63785] = 25'b11111001_00100111_00100000_1;
      patterns[63786] = 25'b11111001_00101000_00100001_1;
      patterns[63787] = 25'b11111001_00101001_00100010_1;
      patterns[63788] = 25'b11111001_00101010_00100011_1;
      patterns[63789] = 25'b11111001_00101011_00100100_1;
      patterns[63790] = 25'b11111001_00101100_00100101_1;
      patterns[63791] = 25'b11111001_00101101_00100110_1;
      patterns[63792] = 25'b11111001_00101110_00100111_1;
      patterns[63793] = 25'b11111001_00101111_00101000_1;
      patterns[63794] = 25'b11111001_00110000_00101001_1;
      patterns[63795] = 25'b11111001_00110001_00101010_1;
      patterns[63796] = 25'b11111001_00110010_00101011_1;
      patterns[63797] = 25'b11111001_00110011_00101100_1;
      patterns[63798] = 25'b11111001_00110100_00101101_1;
      patterns[63799] = 25'b11111001_00110101_00101110_1;
      patterns[63800] = 25'b11111001_00110110_00101111_1;
      patterns[63801] = 25'b11111001_00110111_00110000_1;
      patterns[63802] = 25'b11111001_00111000_00110001_1;
      patterns[63803] = 25'b11111001_00111001_00110010_1;
      patterns[63804] = 25'b11111001_00111010_00110011_1;
      patterns[63805] = 25'b11111001_00111011_00110100_1;
      patterns[63806] = 25'b11111001_00111100_00110101_1;
      patterns[63807] = 25'b11111001_00111101_00110110_1;
      patterns[63808] = 25'b11111001_00111110_00110111_1;
      patterns[63809] = 25'b11111001_00111111_00111000_1;
      patterns[63810] = 25'b11111001_01000000_00111001_1;
      patterns[63811] = 25'b11111001_01000001_00111010_1;
      patterns[63812] = 25'b11111001_01000010_00111011_1;
      patterns[63813] = 25'b11111001_01000011_00111100_1;
      patterns[63814] = 25'b11111001_01000100_00111101_1;
      patterns[63815] = 25'b11111001_01000101_00111110_1;
      patterns[63816] = 25'b11111001_01000110_00111111_1;
      patterns[63817] = 25'b11111001_01000111_01000000_1;
      patterns[63818] = 25'b11111001_01001000_01000001_1;
      patterns[63819] = 25'b11111001_01001001_01000010_1;
      patterns[63820] = 25'b11111001_01001010_01000011_1;
      patterns[63821] = 25'b11111001_01001011_01000100_1;
      patterns[63822] = 25'b11111001_01001100_01000101_1;
      patterns[63823] = 25'b11111001_01001101_01000110_1;
      patterns[63824] = 25'b11111001_01001110_01000111_1;
      patterns[63825] = 25'b11111001_01001111_01001000_1;
      patterns[63826] = 25'b11111001_01010000_01001001_1;
      patterns[63827] = 25'b11111001_01010001_01001010_1;
      patterns[63828] = 25'b11111001_01010010_01001011_1;
      patterns[63829] = 25'b11111001_01010011_01001100_1;
      patterns[63830] = 25'b11111001_01010100_01001101_1;
      patterns[63831] = 25'b11111001_01010101_01001110_1;
      patterns[63832] = 25'b11111001_01010110_01001111_1;
      patterns[63833] = 25'b11111001_01010111_01010000_1;
      patterns[63834] = 25'b11111001_01011000_01010001_1;
      patterns[63835] = 25'b11111001_01011001_01010010_1;
      patterns[63836] = 25'b11111001_01011010_01010011_1;
      patterns[63837] = 25'b11111001_01011011_01010100_1;
      patterns[63838] = 25'b11111001_01011100_01010101_1;
      patterns[63839] = 25'b11111001_01011101_01010110_1;
      patterns[63840] = 25'b11111001_01011110_01010111_1;
      patterns[63841] = 25'b11111001_01011111_01011000_1;
      patterns[63842] = 25'b11111001_01100000_01011001_1;
      patterns[63843] = 25'b11111001_01100001_01011010_1;
      patterns[63844] = 25'b11111001_01100010_01011011_1;
      patterns[63845] = 25'b11111001_01100011_01011100_1;
      patterns[63846] = 25'b11111001_01100100_01011101_1;
      patterns[63847] = 25'b11111001_01100101_01011110_1;
      patterns[63848] = 25'b11111001_01100110_01011111_1;
      patterns[63849] = 25'b11111001_01100111_01100000_1;
      patterns[63850] = 25'b11111001_01101000_01100001_1;
      patterns[63851] = 25'b11111001_01101001_01100010_1;
      patterns[63852] = 25'b11111001_01101010_01100011_1;
      patterns[63853] = 25'b11111001_01101011_01100100_1;
      patterns[63854] = 25'b11111001_01101100_01100101_1;
      patterns[63855] = 25'b11111001_01101101_01100110_1;
      patterns[63856] = 25'b11111001_01101110_01100111_1;
      patterns[63857] = 25'b11111001_01101111_01101000_1;
      patterns[63858] = 25'b11111001_01110000_01101001_1;
      patterns[63859] = 25'b11111001_01110001_01101010_1;
      patterns[63860] = 25'b11111001_01110010_01101011_1;
      patterns[63861] = 25'b11111001_01110011_01101100_1;
      patterns[63862] = 25'b11111001_01110100_01101101_1;
      patterns[63863] = 25'b11111001_01110101_01101110_1;
      patterns[63864] = 25'b11111001_01110110_01101111_1;
      patterns[63865] = 25'b11111001_01110111_01110000_1;
      patterns[63866] = 25'b11111001_01111000_01110001_1;
      patterns[63867] = 25'b11111001_01111001_01110010_1;
      patterns[63868] = 25'b11111001_01111010_01110011_1;
      patterns[63869] = 25'b11111001_01111011_01110100_1;
      patterns[63870] = 25'b11111001_01111100_01110101_1;
      patterns[63871] = 25'b11111001_01111101_01110110_1;
      patterns[63872] = 25'b11111001_01111110_01110111_1;
      patterns[63873] = 25'b11111001_01111111_01111000_1;
      patterns[63874] = 25'b11111001_10000000_01111001_1;
      patterns[63875] = 25'b11111001_10000001_01111010_1;
      patterns[63876] = 25'b11111001_10000010_01111011_1;
      patterns[63877] = 25'b11111001_10000011_01111100_1;
      patterns[63878] = 25'b11111001_10000100_01111101_1;
      patterns[63879] = 25'b11111001_10000101_01111110_1;
      patterns[63880] = 25'b11111001_10000110_01111111_1;
      patterns[63881] = 25'b11111001_10000111_10000000_1;
      patterns[63882] = 25'b11111001_10001000_10000001_1;
      patterns[63883] = 25'b11111001_10001001_10000010_1;
      patterns[63884] = 25'b11111001_10001010_10000011_1;
      patterns[63885] = 25'b11111001_10001011_10000100_1;
      patterns[63886] = 25'b11111001_10001100_10000101_1;
      patterns[63887] = 25'b11111001_10001101_10000110_1;
      patterns[63888] = 25'b11111001_10001110_10000111_1;
      patterns[63889] = 25'b11111001_10001111_10001000_1;
      patterns[63890] = 25'b11111001_10010000_10001001_1;
      patterns[63891] = 25'b11111001_10010001_10001010_1;
      patterns[63892] = 25'b11111001_10010010_10001011_1;
      patterns[63893] = 25'b11111001_10010011_10001100_1;
      patterns[63894] = 25'b11111001_10010100_10001101_1;
      patterns[63895] = 25'b11111001_10010101_10001110_1;
      patterns[63896] = 25'b11111001_10010110_10001111_1;
      patterns[63897] = 25'b11111001_10010111_10010000_1;
      patterns[63898] = 25'b11111001_10011000_10010001_1;
      patterns[63899] = 25'b11111001_10011001_10010010_1;
      patterns[63900] = 25'b11111001_10011010_10010011_1;
      patterns[63901] = 25'b11111001_10011011_10010100_1;
      patterns[63902] = 25'b11111001_10011100_10010101_1;
      patterns[63903] = 25'b11111001_10011101_10010110_1;
      patterns[63904] = 25'b11111001_10011110_10010111_1;
      patterns[63905] = 25'b11111001_10011111_10011000_1;
      patterns[63906] = 25'b11111001_10100000_10011001_1;
      patterns[63907] = 25'b11111001_10100001_10011010_1;
      patterns[63908] = 25'b11111001_10100010_10011011_1;
      patterns[63909] = 25'b11111001_10100011_10011100_1;
      patterns[63910] = 25'b11111001_10100100_10011101_1;
      patterns[63911] = 25'b11111001_10100101_10011110_1;
      patterns[63912] = 25'b11111001_10100110_10011111_1;
      patterns[63913] = 25'b11111001_10100111_10100000_1;
      patterns[63914] = 25'b11111001_10101000_10100001_1;
      patterns[63915] = 25'b11111001_10101001_10100010_1;
      patterns[63916] = 25'b11111001_10101010_10100011_1;
      patterns[63917] = 25'b11111001_10101011_10100100_1;
      patterns[63918] = 25'b11111001_10101100_10100101_1;
      patterns[63919] = 25'b11111001_10101101_10100110_1;
      patterns[63920] = 25'b11111001_10101110_10100111_1;
      patterns[63921] = 25'b11111001_10101111_10101000_1;
      patterns[63922] = 25'b11111001_10110000_10101001_1;
      patterns[63923] = 25'b11111001_10110001_10101010_1;
      patterns[63924] = 25'b11111001_10110010_10101011_1;
      patterns[63925] = 25'b11111001_10110011_10101100_1;
      patterns[63926] = 25'b11111001_10110100_10101101_1;
      patterns[63927] = 25'b11111001_10110101_10101110_1;
      patterns[63928] = 25'b11111001_10110110_10101111_1;
      patterns[63929] = 25'b11111001_10110111_10110000_1;
      patterns[63930] = 25'b11111001_10111000_10110001_1;
      patterns[63931] = 25'b11111001_10111001_10110010_1;
      patterns[63932] = 25'b11111001_10111010_10110011_1;
      patterns[63933] = 25'b11111001_10111011_10110100_1;
      patterns[63934] = 25'b11111001_10111100_10110101_1;
      patterns[63935] = 25'b11111001_10111101_10110110_1;
      patterns[63936] = 25'b11111001_10111110_10110111_1;
      patterns[63937] = 25'b11111001_10111111_10111000_1;
      patterns[63938] = 25'b11111001_11000000_10111001_1;
      patterns[63939] = 25'b11111001_11000001_10111010_1;
      patterns[63940] = 25'b11111001_11000010_10111011_1;
      patterns[63941] = 25'b11111001_11000011_10111100_1;
      patterns[63942] = 25'b11111001_11000100_10111101_1;
      patterns[63943] = 25'b11111001_11000101_10111110_1;
      patterns[63944] = 25'b11111001_11000110_10111111_1;
      patterns[63945] = 25'b11111001_11000111_11000000_1;
      patterns[63946] = 25'b11111001_11001000_11000001_1;
      patterns[63947] = 25'b11111001_11001001_11000010_1;
      patterns[63948] = 25'b11111001_11001010_11000011_1;
      patterns[63949] = 25'b11111001_11001011_11000100_1;
      patterns[63950] = 25'b11111001_11001100_11000101_1;
      patterns[63951] = 25'b11111001_11001101_11000110_1;
      patterns[63952] = 25'b11111001_11001110_11000111_1;
      patterns[63953] = 25'b11111001_11001111_11001000_1;
      patterns[63954] = 25'b11111001_11010000_11001001_1;
      patterns[63955] = 25'b11111001_11010001_11001010_1;
      patterns[63956] = 25'b11111001_11010010_11001011_1;
      patterns[63957] = 25'b11111001_11010011_11001100_1;
      patterns[63958] = 25'b11111001_11010100_11001101_1;
      patterns[63959] = 25'b11111001_11010101_11001110_1;
      patterns[63960] = 25'b11111001_11010110_11001111_1;
      patterns[63961] = 25'b11111001_11010111_11010000_1;
      patterns[63962] = 25'b11111001_11011000_11010001_1;
      patterns[63963] = 25'b11111001_11011001_11010010_1;
      patterns[63964] = 25'b11111001_11011010_11010011_1;
      patterns[63965] = 25'b11111001_11011011_11010100_1;
      patterns[63966] = 25'b11111001_11011100_11010101_1;
      patterns[63967] = 25'b11111001_11011101_11010110_1;
      patterns[63968] = 25'b11111001_11011110_11010111_1;
      patterns[63969] = 25'b11111001_11011111_11011000_1;
      patterns[63970] = 25'b11111001_11100000_11011001_1;
      patterns[63971] = 25'b11111001_11100001_11011010_1;
      patterns[63972] = 25'b11111001_11100010_11011011_1;
      patterns[63973] = 25'b11111001_11100011_11011100_1;
      patterns[63974] = 25'b11111001_11100100_11011101_1;
      patterns[63975] = 25'b11111001_11100101_11011110_1;
      patterns[63976] = 25'b11111001_11100110_11011111_1;
      patterns[63977] = 25'b11111001_11100111_11100000_1;
      patterns[63978] = 25'b11111001_11101000_11100001_1;
      patterns[63979] = 25'b11111001_11101001_11100010_1;
      patterns[63980] = 25'b11111001_11101010_11100011_1;
      patterns[63981] = 25'b11111001_11101011_11100100_1;
      patterns[63982] = 25'b11111001_11101100_11100101_1;
      patterns[63983] = 25'b11111001_11101101_11100110_1;
      patterns[63984] = 25'b11111001_11101110_11100111_1;
      patterns[63985] = 25'b11111001_11101111_11101000_1;
      patterns[63986] = 25'b11111001_11110000_11101001_1;
      patterns[63987] = 25'b11111001_11110001_11101010_1;
      patterns[63988] = 25'b11111001_11110010_11101011_1;
      patterns[63989] = 25'b11111001_11110011_11101100_1;
      patterns[63990] = 25'b11111001_11110100_11101101_1;
      patterns[63991] = 25'b11111001_11110101_11101110_1;
      patterns[63992] = 25'b11111001_11110110_11101111_1;
      patterns[63993] = 25'b11111001_11110111_11110000_1;
      patterns[63994] = 25'b11111001_11111000_11110001_1;
      patterns[63995] = 25'b11111001_11111001_11110010_1;
      patterns[63996] = 25'b11111001_11111010_11110011_1;
      patterns[63997] = 25'b11111001_11111011_11110100_1;
      patterns[63998] = 25'b11111001_11111100_11110101_1;
      patterns[63999] = 25'b11111001_11111101_11110110_1;
      patterns[64000] = 25'b11111001_11111110_11110111_1;
      patterns[64001] = 25'b11111001_11111111_11111000_1;
      patterns[64002] = 25'b11111010_00000000_11111010_0;
      patterns[64003] = 25'b11111010_00000001_11111011_0;
      patterns[64004] = 25'b11111010_00000010_11111100_0;
      patterns[64005] = 25'b11111010_00000011_11111101_0;
      patterns[64006] = 25'b11111010_00000100_11111110_0;
      patterns[64007] = 25'b11111010_00000101_11111111_0;
      patterns[64008] = 25'b11111010_00000110_00000000_1;
      patterns[64009] = 25'b11111010_00000111_00000001_1;
      patterns[64010] = 25'b11111010_00001000_00000010_1;
      patterns[64011] = 25'b11111010_00001001_00000011_1;
      patterns[64012] = 25'b11111010_00001010_00000100_1;
      patterns[64013] = 25'b11111010_00001011_00000101_1;
      patterns[64014] = 25'b11111010_00001100_00000110_1;
      patterns[64015] = 25'b11111010_00001101_00000111_1;
      patterns[64016] = 25'b11111010_00001110_00001000_1;
      patterns[64017] = 25'b11111010_00001111_00001001_1;
      patterns[64018] = 25'b11111010_00010000_00001010_1;
      patterns[64019] = 25'b11111010_00010001_00001011_1;
      patterns[64020] = 25'b11111010_00010010_00001100_1;
      patterns[64021] = 25'b11111010_00010011_00001101_1;
      patterns[64022] = 25'b11111010_00010100_00001110_1;
      patterns[64023] = 25'b11111010_00010101_00001111_1;
      patterns[64024] = 25'b11111010_00010110_00010000_1;
      patterns[64025] = 25'b11111010_00010111_00010001_1;
      patterns[64026] = 25'b11111010_00011000_00010010_1;
      patterns[64027] = 25'b11111010_00011001_00010011_1;
      patterns[64028] = 25'b11111010_00011010_00010100_1;
      patterns[64029] = 25'b11111010_00011011_00010101_1;
      patterns[64030] = 25'b11111010_00011100_00010110_1;
      patterns[64031] = 25'b11111010_00011101_00010111_1;
      patterns[64032] = 25'b11111010_00011110_00011000_1;
      patterns[64033] = 25'b11111010_00011111_00011001_1;
      patterns[64034] = 25'b11111010_00100000_00011010_1;
      patterns[64035] = 25'b11111010_00100001_00011011_1;
      patterns[64036] = 25'b11111010_00100010_00011100_1;
      patterns[64037] = 25'b11111010_00100011_00011101_1;
      patterns[64038] = 25'b11111010_00100100_00011110_1;
      patterns[64039] = 25'b11111010_00100101_00011111_1;
      patterns[64040] = 25'b11111010_00100110_00100000_1;
      patterns[64041] = 25'b11111010_00100111_00100001_1;
      patterns[64042] = 25'b11111010_00101000_00100010_1;
      patterns[64043] = 25'b11111010_00101001_00100011_1;
      patterns[64044] = 25'b11111010_00101010_00100100_1;
      patterns[64045] = 25'b11111010_00101011_00100101_1;
      patterns[64046] = 25'b11111010_00101100_00100110_1;
      patterns[64047] = 25'b11111010_00101101_00100111_1;
      patterns[64048] = 25'b11111010_00101110_00101000_1;
      patterns[64049] = 25'b11111010_00101111_00101001_1;
      patterns[64050] = 25'b11111010_00110000_00101010_1;
      patterns[64051] = 25'b11111010_00110001_00101011_1;
      patterns[64052] = 25'b11111010_00110010_00101100_1;
      patterns[64053] = 25'b11111010_00110011_00101101_1;
      patterns[64054] = 25'b11111010_00110100_00101110_1;
      patterns[64055] = 25'b11111010_00110101_00101111_1;
      patterns[64056] = 25'b11111010_00110110_00110000_1;
      patterns[64057] = 25'b11111010_00110111_00110001_1;
      patterns[64058] = 25'b11111010_00111000_00110010_1;
      patterns[64059] = 25'b11111010_00111001_00110011_1;
      patterns[64060] = 25'b11111010_00111010_00110100_1;
      patterns[64061] = 25'b11111010_00111011_00110101_1;
      patterns[64062] = 25'b11111010_00111100_00110110_1;
      patterns[64063] = 25'b11111010_00111101_00110111_1;
      patterns[64064] = 25'b11111010_00111110_00111000_1;
      patterns[64065] = 25'b11111010_00111111_00111001_1;
      patterns[64066] = 25'b11111010_01000000_00111010_1;
      patterns[64067] = 25'b11111010_01000001_00111011_1;
      patterns[64068] = 25'b11111010_01000010_00111100_1;
      patterns[64069] = 25'b11111010_01000011_00111101_1;
      patterns[64070] = 25'b11111010_01000100_00111110_1;
      patterns[64071] = 25'b11111010_01000101_00111111_1;
      patterns[64072] = 25'b11111010_01000110_01000000_1;
      patterns[64073] = 25'b11111010_01000111_01000001_1;
      patterns[64074] = 25'b11111010_01001000_01000010_1;
      patterns[64075] = 25'b11111010_01001001_01000011_1;
      patterns[64076] = 25'b11111010_01001010_01000100_1;
      patterns[64077] = 25'b11111010_01001011_01000101_1;
      patterns[64078] = 25'b11111010_01001100_01000110_1;
      patterns[64079] = 25'b11111010_01001101_01000111_1;
      patterns[64080] = 25'b11111010_01001110_01001000_1;
      patterns[64081] = 25'b11111010_01001111_01001001_1;
      patterns[64082] = 25'b11111010_01010000_01001010_1;
      patterns[64083] = 25'b11111010_01010001_01001011_1;
      patterns[64084] = 25'b11111010_01010010_01001100_1;
      patterns[64085] = 25'b11111010_01010011_01001101_1;
      patterns[64086] = 25'b11111010_01010100_01001110_1;
      patterns[64087] = 25'b11111010_01010101_01001111_1;
      patterns[64088] = 25'b11111010_01010110_01010000_1;
      patterns[64089] = 25'b11111010_01010111_01010001_1;
      patterns[64090] = 25'b11111010_01011000_01010010_1;
      patterns[64091] = 25'b11111010_01011001_01010011_1;
      patterns[64092] = 25'b11111010_01011010_01010100_1;
      patterns[64093] = 25'b11111010_01011011_01010101_1;
      patterns[64094] = 25'b11111010_01011100_01010110_1;
      patterns[64095] = 25'b11111010_01011101_01010111_1;
      patterns[64096] = 25'b11111010_01011110_01011000_1;
      patterns[64097] = 25'b11111010_01011111_01011001_1;
      patterns[64098] = 25'b11111010_01100000_01011010_1;
      patterns[64099] = 25'b11111010_01100001_01011011_1;
      patterns[64100] = 25'b11111010_01100010_01011100_1;
      patterns[64101] = 25'b11111010_01100011_01011101_1;
      patterns[64102] = 25'b11111010_01100100_01011110_1;
      patterns[64103] = 25'b11111010_01100101_01011111_1;
      patterns[64104] = 25'b11111010_01100110_01100000_1;
      patterns[64105] = 25'b11111010_01100111_01100001_1;
      patterns[64106] = 25'b11111010_01101000_01100010_1;
      patterns[64107] = 25'b11111010_01101001_01100011_1;
      patterns[64108] = 25'b11111010_01101010_01100100_1;
      patterns[64109] = 25'b11111010_01101011_01100101_1;
      patterns[64110] = 25'b11111010_01101100_01100110_1;
      patterns[64111] = 25'b11111010_01101101_01100111_1;
      patterns[64112] = 25'b11111010_01101110_01101000_1;
      patterns[64113] = 25'b11111010_01101111_01101001_1;
      patterns[64114] = 25'b11111010_01110000_01101010_1;
      patterns[64115] = 25'b11111010_01110001_01101011_1;
      patterns[64116] = 25'b11111010_01110010_01101100_1;
      patterns[64117] = 25'b11111010_01110011_01101101_1;
      patterns[64118] = 25'b11111010_01110100_01101110_1;
      patterns[64119] = 25'b11111010_01110101_01101111_1;
      patterns[64120] = 25'b11111010_01110110_01110000_1;
      patterns[64121] = 25'b11111010_01110111_01110001_1;
      patterns[64122] = 25'b11111010_01111000_01110010_1;
      patterns[64123] = 25'b11111010_01111001_01110011_1;
      patterns[64124] = 25'b11111010_01111010_01110100_1;
      patterns[64125] = 25'b11111010_01111011_01110101_1;
      patterns[64126] = 25'b11111010_01111100_01110110_1;
      patterns[64127] = 25'b11111010_01111101_01110111_1;
      patterns[64128] = 25'b11111010_01111110_01111000_1;
      patterns[64129] = 25'b11111010_01111111_01111001_1;
      patterns[64130] = 25'b11111010_10000000_01111010_1;
      patterns[64131] = 25'b11111010_10000001_01111011_1;
      patterns[64132] = 25'b11111010_10000010_01111100_1;
      patterns[64133] = 25'b11111010_10000011_01111101_1;
      patterns[64134] = 25'b11111010_10000100_01111110_1;
      patterns[64135] = 25'b11111010_10000101_01111111_1;
      patterns[64136] = 25'b11111010_10000110_10000000_1;
      patterns[64137] = 25'b11111010_10000111_10000001_1;
      patterns[64138] = 25'b11111010_10001000_10000010_1;
      patterns[64139] = 25'b11111010_10001001_10000011_1;
      patterns[64140] = 25'b11111010_10001010_10000100_1;
      patterns[64141] = 25'b11111010_10001011_10000101_1;
      patterns[64142] = 25'b11111010_10001100_10000110_1;
      patterns[64143] = 25'b11111010_10001101_10000111_1;
      patterns[64144] = 25'b11111010_10001110_10001000_1;
      patterns[64145] = 25'b11111010_10001111_10001001_1;
      patterns[64146] = 25'b11111010_10010000_10001010_1;
      patterns[64147] = 25'b11111010_10010001_10001011_1;
      patterns[64148] = 25'b11111010_10010010_10001100_1;
      patterns[64149] = 25'b11111010_10010011_10001101_1;
      patterns[64150] = 25'b11111010_10010100_10001110_1;
      patterns[64151] = 25'b11111010_10010101_10001111_1;
      patterns[64152] = 25'b11111010_10010110_10010000_1;
      patterns[64153] = 25'b11111010_10010111_10010001_1;
      patterns[64154] = 25'b11111010_10011000_10010010_1;
      patterns[64155] = 25'b11111010_10011001_10010011_1;
      patterns[64156] = 25'b11111010_10011010_10010100_1;
      patterns[64157] = 25'b11111010_10011011_10010101_1;
      patterns[64158] = 25'b11111010_10011100_10010110_1;
      patterns[64159] = 25'b11111010_10011101_10010111_1;
      patterns[64160] = 25'b11111010_10011110_10011000_1;
      patterns[64161] = 25'b11111010_10011111_10011001_1;
      patterns[64162] = 25'b11111010_10100000_10011010_1;
      patterns[64163] = 25'b11111010_10100001_10011011_1;
      patterns[64164] = 25'b11111010_10100010_10011100_1;
      patterns[64165] = 25'b11111010_10100011_10011101_1;
      patterns[64166] = 25'b11111010_10100100_10011110_1;
      patterns[64167] = 25'b11111010_10100101_10011111_1;
      patterns[64168] = 25'b11111010_10100110_10100000_1;
      patterns[64169] = 25'b11111010_10100111_10100001_1;
      patterns[64170] = 25'b11111010_10101000_10100010_1;
      patterns[64171] = 25'b11111010_10101001_10100011_1;
      patterns[64172] = 25'b11111010_10101010_10100100_1;
      patterns[64173] = 25'b11111010_10101011_10100101_1;
      patterns[64174] = 25'b11111010_10101100_10100110_1;
      patterns[64175] = 25'b11111010_10101101_10100111_1;
      patterns[64176] = 25'b11111010_10101110_10101000_1;
      patterns[64177] = 25'b11111010_10101111_10101001_1;
      patterns[64178] = 25'b11111010_10110000_10101010_1;
      patterns[64179] = 25'b11111010_10110001_10101011_1;
      patterns[64180] = 25'b11111010_10110010_10101100_1;
      patterns[64181] = 25'b11111010_10110011_10101101_1;
      patterns[64182] = 25'b11111010_10110100_10101110_1;
      patterns[64183] = 25'b11111010_10110101_10101111_1;
      patterns[64184] = 25'b11111010_10110110_10110000_1;
      patterns[64185] = 25'b11111010_10110111_10110001_1;
      patterns[64186] = 25'b11111010_10111000_10110010_1;
      patterns[64187] = 25'b11111010_10111001_10110011_1;
      patterns[64188] = 25'b11111010_10111010_10110100_1;
      patterns[64189] = 25'b11111010_10111011_10110101_1;
      patterns[64190] = 25'b11111010_10111100_10110110_1;
      patterns[64191] = 25'b11111010_10111101_10110111_1;
      patterns[64192] = 25'b11111010_10111110_10111000_1;
      patterns[64193] = 25'b11111010_10111111_10111001_1;
      patterns[64194] = 25'b11111010_11000000_10111010_1;
      patterns[64195] = 25'b11111010_11000001_10111011_1;
      patterns[64196] = 25'b11111010_11000010_10111100_1;
      patterns[64197] = 25'b11111010_11000011_10111101_1;
      patterns[64198] = 25'b11111010_11000100_10111110_1;
      patterns[64199] = 25'b11111010_11000101_10111111_1;
      patterns[64200] = 25'b11111010_11000110_11000000_1;
      patterns[64201] = 25'b11111010_11000111_11000001_1;
      patterns[64202] = 25'b11111010_11001000_11000010_1;
      patterns[64203] = 25'b11111010_11001001_11000011_1;
      patterns[64204] = 25'b11111010_11001010_11000100_1;
      patterns[64205] = 25'b11111010_11001011_11000101_1;
      patterns[64206] = 25'b11111010_11001100_11000110_1;
      patterns[64207] = 25'b11111010_11001101_11000111_1;
      patterns[64208] = 25'b11111010_11001110_11001000_1;
      patterns[64209] = 25'b11111010_11001111_11001001_1;
      patterns[64210] = 25'b11111010_11010000_11001010_1;
      patterns[64211] = 25'b11111010_11010001_11001011_1;
      patterns[64212] = 25'b11111010_11010010_11001100_1;
      patterns[64213] = 25'b11111010_11010011_11001101_1;
      patterns[64214] = 25'b11111010_11010100_11001110_1;
      patterns[64215] = 25'b11111010_11010101_11001111_1;
      patterns[64216] = 25'b11111010_11010110_11010000_1;
      patterns[64217] = 25'b11111010_11010111_11010001_1;
      patterns[64218] = 25'b11111010_11011000_11010010_1;
      patterns[64219] = 25'b11111010_11011001_11010011_1;
      patterns[64220] = 25'b11111010_11011010_11010100_1;
      patterns[64221] = 25'b11111010_11011011_11010101_1;
      patterns[64222] = 25'b11111010_11011100_11010110_1;
      patterns[64223] = 25'b11111010_11011101_11010111_1;
      patterns[64224] = 25'b11111010_11011110_11011000_1;
      patterns[64225] = 25'b11111010_11011111_11011001_1;
      patterns[64226] = 25'b11111010_11100000_11011010_1;
      patterns[64227] = 25'b11111010_11100001_11011011_1;
      patterns[64228] = 25'b11111010_11100010_11011100_1;
      patterns[64229] = 25'b11111010_11100011_11011101_1;
      patterns[64230] = 25'b11111010_11100100_11011110_1;
      patterns[64231] = 25'b11111010_11100101_11011111_1;
      patterns[64232] = 25'b11111010_11100110_11100000_1;
      patterns[64233] = 25'b11111010_11100111_11100001_1;
      patterns[64234] = 25'b11111010_11101000_11100010_1;
      patterns[64235] = 25'b11111010_11101001_11100011_1;
      patterns[64236] = 25'b11111010_11101010_11100100_1;
      patterns[64237] = 25'b11111010_11101011_11100101_1;
      patterns[64238] = 25'b11111010_11101100_11100110_1;
      patterns[64239] = 25'b11111010_11101101_11100111_1;
      patterns[64240] = 25'b11111010_11101110_11101000_1;
      patterns[64241] = 25'b11111010_11101111_11101001_1;
      patterns[64242] = 25'b11111010_11110000_11101010_1;
      patterns[64243] = 25'b11111010_11110001_11101011_1;
      patterns[64244] = 25'b11111010_11110010_11101100_1;
      patterns[64245] = 25'b11111010_11110011_11101101_1;
      patterns[64246] = 25'b11111010_11110100_11101110_1;
      patterns[64247] = 25'b11111010_11110101_11101111_1;
      patterns[64248] = 25'b11111010_11110110_11110000_1;
      patterns[64249] = 25'b11111010_11110111_11110001_1;
      patterns[64250] = 25'b11111010_11111000_11110010_1;
      patterns[64251] = 25'b11111010_11111001_11110011_1;
      patterns[64252] = 25'b11111010_11111010_11110100_1;
      patterns[64253] = 25'b11111010_11111011_11110101_1;
      patterns[64254] = 25'b11111010_11111100_11110110_1;
      patterns[64255] = 25'b11111010_11111101_11110111_1;
      patterns[64256] = 25'b11111010_11111110_11111000_1;
      patterns[64257] = 25'b11111010_11111111_11111001_1;
      patterns[64258] = 25'b11111011_00000000_11111011_0;
      patterns[64259] = 25'b11111011_00000001_11111100_0;
      patterns[64260] = 25'b11111011_00000010_11111101_0;
      patterns[64261] = 25'b11111011_00000011_11111110_0;
      patterns[64262] = 25'b11111011_00000100_11111111_0;
      patterns[64263] = 25'b11111011_00000101_00000000_1;
      patterns[64264] = 25'b11111011_00000110_00000001_1;
      patterns[64265] = 25'b11111011_00000111_00000010_1;
      patterns[64266] = 25'b11111011_00001000_00000011_1;
      patterns[64267] = 25'b11111011_00001001_00000100_1;
      patterns[64268] = 25'b11111011_00001010_00000101_1;
      patterns[64269] = 25'b11111011_00001011_00000110_1;
      patterns[64270] = 25'b11111011_00001100_00000111_1;
      patterns[64271] = 25'b11111011_00001101_00001000_1;
      patterns[64272] = 25'b11111011_00001110_00001001_1;
      patterns[64273] = 25'b11111011_00001111_00001010_1;
      patterns[64274] = 25'b11111011_00010000_00001011_1;
      patterns[64275] = 25'b11111011_00010001_00001100_1;
      patterns[64276] = 25'b11111011_00010010_00001101_1;
      patterns[64277] = 25'b11111011_00010011_00001110_1;
      patterns[64278] = 25'b11111011_00010100_00001111_1;
      patterns[64279] = 25'b11111011_00010101_00010000_1;
      patterns[64280] = 25'b11111011_00010110_00010001_1;
      patterns[64281] = 25'b11111011_00010111_00010010_1;
      patterns[64282] = 25'b11111011_00011000_00010011_1;
      patterns[64283] = 25'b11111011_00011001_00010100_1;
      patterns[64284] = 25'b11111011_00011010_00010101_1;
      patterns[64285] = 25'b11111011_00011011_00010110_1;
      patterns[64286] = 25'b11111011_00011100_00010111_1;
      patterns[64287] = 25'b11111011_00011101_00011000_1;
      patterns[64288] = 25'b11111011_00011110_00011001_1;
      patterns[64289] = 25'b11111011_00011111_00011010_1;
      patterns[64290] = 25'b11111011_00100000_00011011_1;
      patterns[64291] = 25'b11111011_00100001_00011100_1;
      patterns[64292] = 25'b11111011_00100010_00011101_1;
      patterns[64293] = 25'b11111011_00100011_00011110_1;
      patterns[64294] = 25'b11111011_00100100_00011111_1;
      patterns[64295] = 25'b11111011_00100101_00100000_1;
      patterns[64296] = 25'b11111011_00100110_00100001_1;
      patterns[64297] = 25'b11111011_00100111_00100010_1;
      patterns[64298] = 25'b11111011_00101000_00100011_1;
      patterns[64299] = 25'b11111011_00101001_00100100_1;
      patterns[64300] = 25'b11111011_00101010_00100101_1;
      patterns[64301] = 25'b11111011_00101011_00100110_1;
      patterns[64302] = 25'b11111011_00101100_00100111_1;
      patterns[64303] = 25'b11111011_00101101_00101000_1;
      patterns[64304] = 25'b11111011_00101110_00101001_1;
      patterns[64305] = 25'b11111011_00101111_00101010_1;
      patterns[64306] = 25'b11111011_00110000_00101011_1;
      patterns[64307] = 25'b11111011_00110001_00101100_1;
      patterns[64308] = 25'b11111011_00110010_00101101_1;
      patterns[64309] = 25'b11111011_00110011_00101110_1;
      patterns[64310] = 25'b11111011_00110100_00101111_1;
      patterns[64311] = 25'b11111011_00110101_00110000_1;
      patterns[64312] = 25'b11111011_00110110_00110001_1;
      patterns[64313] = 25'b11111011_00110111_00110010_1;
      patterns[64314] = 25'b11111011_00111000_00110011_1;
      patterns[64315] = 25'b11111011_00111001_00110100_1;
      patterns[64316] = 25'b11111011_00111010_00110101_1;
      patterns[64317] = 25'b11111011_00111011_00110110_1;
      patterns[64318] = 25'b11111011_00111100_00110111_1;
      patterns[64319] = 25'b11111011_00111101_00111000_1;
      patterns[64320] = 25'b11111011_00111110_00111001_1;
      patterns[64321] = 25'b11111011_00111111_00111010_1;
      patterns[64322] = 25'b11111011_01000000_00111011_1;
      patterns[64323] = 25'b11111011_01000001_00111100_1;
      patterns[64324] = 25'b11111011_01000010_00111101_1;
      patterns[64325] = 25'b11111011_01000011_00111110_1;
      patterns[64326] = 25'b11111011_01000100_00111111_1;
      patterns[64327] = 25'b11111011_01000101_01000000_1;
      patterns[64328] = 25'b11111011_01000110_01000001_1;
      patterns[64329] = 25'b11111011_01000111_01000010_1;
      patterns[64330] = 25'b11111011_01001000_01000011_1;
      patterns[64331] = 25'b11111011_01001001_01000100_1;
      patterns[64332] = 25'b11111011_01001010_01000101_1;
      patterns[64333] = 25'b11111011_01001011_01000110_1;
      patterns[64334] = 25'b11111011_01001100_01000111_1;
      patterns[64335] = 25'b11111011_01001101_01001000_1;
      patterns[64336] = 25'b11111011_01001110_01001001_1;
      patterns[64337] = 25'b11111011_01001111_01001010_1;
      patterns[64338] = 25'b11111011_01010000_01001011_1;
      patterns[64339] = 25'b11111011_01010001_01001100_1;
      patterns[64340] = 25'b11111011_01010010_01001101_1;
      patterns[64341] = 25'b11111011_01010011_01001110_1;
      patterns[64342] = 25'b11111011_01010100_01001111_1;
      patterns[64343] = 25'b11111011_01010101_01010000_1;
      patterns[64344] = 25'b11111011_01010110_01010001_1;
      patterns[64345] = 25'b11111011_01010111_01010010_1;
      patterns[64346] = 25'b11111011_01011000_01010011_1;
      patterns[64347] = 25'b11111011_01011001_01010100_1;
      patterns[64348] = 25'b11111011_01011010_01010101_1;
      patterns[64349] = 25'b11111011_01011011_01010110_1;
      patterns[64350] = 25'b11111011_01011100_01010111_1;
      patterns[64351] = 25'b11111011_01011101_01011000_1;
      patterns[64352] = 25'b11111011_01011110_01011001_1;
      patterns[64353] = 25'b11111011_01011111_01011010_1;
      patterns[64354] = 25'b11111011_01100000_01011011_1;
      patterns[64355] = 25'b11111011_01100001_01011100_1;
      patterns[64356] = 25'b11111011_01100010_01011101_1;
      patterns[64357] = 25'b11111011_01100011_01011110_1;
      patterns[64358] = 25'b11111011_01100100_01011111_1;
      patterns[64359] = 25'b11111011_01100101_01100000_1;
      patterns[64360] = 25'b11111011_01100110_01100001_1;
      patterns[64361] = 25'b11111011_01100111_01100010_1;
      patterns[64362] = 25'b11111011_01101000_01100011_1;
      patterns[64363] = 25'b11111011_01101001_01100100_1;
      patterns[64364] = 25'b11111011_01101010_01100101_1;
      patterns[64365] = 25'b11111011_01101011_01100110_1;
      patterns[64366] = 25'b11111011_01101100_01100111_1;
      patterns[64367] = 25'b11111011_01101101_01101000_1;
      patterns[64368] = 25'b11111011_01101110_01101001_1;
      patterns[64369] = 25'b11111011_01101111_01101010_1;
      patterns[64370] = 25'b11111011_01110000_01101011_1;
      patterns[64371] = 25'b11111011_01110001_01101100_1;
      patterns[64372] = 25'b11111011_01110010_01101101_1;
      patterns[64373] = 25'b11111011_01110011_01101110_1;
      patterns[64374] = 25'b11111011_01110100_01101111_1;
      patterns[64375] = 25'b11111011_01110101_01110000_1;
      patterns[64376] = 25'b11111011_01110110_01110001_1;
      patterns[64377] = 25'b11111011_01110111_01110010_1;
      patterns[64378] = 25'b11111011_01111000_01110011_1;
      patterns[64379] = 25'b11111011_01111001_01110100_1;
      patterns[64380] = 25'b11111011_01111010_01110101_1;
      patterns[64381] = 25'b11111011_01111011_01110110_1;
      patterns[64382] = 25'b11111011_01111100_01110111_1;
      patterns[64383] = 25'b11111011_01111101_01111000_1;
      patterns[64384] = 25'b11111011_01111110_01111001_1;
      patterns[64385] = 25'b11111011_01111111_01111010_1;
      patterns[64386] = 25'b11111011_10000000_01111011_1;
      patterns[64387] = 25'b11111011_10000001_01111100_1;
      patterns[64388] = 25'b11111011_10000010_01111101_1;
      patterns[64389] = 25'b11111011_10000011_01111110_1;
      patterns[64390] = 25'b11111011_10000100_01111111_1;
      patterns[64391] = 25'b11111011_10000101_10000000_1;
      patterns[64392] = 25'b11111011_10000110_10000001_1;
      patterns[64393] = 25'b11111011_10000111_10000010_1;
      patterns[64394] = 25'b11111011_10001000_10000011_1;
      patterns[64395] = 25'b11111011_10001001_10000100_1;
      patterns[64396] = 25'b11111011_10001010_10000101_1;
      patterns[64397] = 25'b11111011_10001011_10000110_1;
      patterns[64398] = 25'b11111011_10001100_10000111_1;
      patterns[64399] = 25'b11111011_10001101_10001000_1;
      patterns[64400] = 25'b11111011_10001110_10001001_1;
      patterns[64401] = 25'b11111011_10001111_10001010_1;
      patterns[64402] = 25'b11111011_10010000_10001011_1;
      patterns[64403] = 25'b11111011_10010001_10001100_1;
      patterns[64404] = 25'b11111011_10010010_10001101_1;
      patterns[64405] = 25'b11111011_10010011_10001110_1;
      patterns[64406] = 25'b11111011_10010100_10001111_1;
      patterns[64407] = 25'b11111011_10010101_10010000_1;
      patterns[64408] = 25'b11111011_10010110_10010001_1;
      patterns[64409] = 25'b11111011_10010111_10010010_1;
      patterns[64410] = 25'b11111011_10011000_10010011_1;
      patterns[64411] = 25'b11111011_10011001_10010100_1;
      patterns[64412] = 25'b11111011_10011010_10010101_1;
      patterns[64413] = 25'b11111011_10011011_10010110_1;
      patterns[64414] = 25'b11111011_10011100_10010111_1;
      patterns[64415] = 25'b11111011_10011101_10011000_1;
      patterns[64416] = 25'b11111011_10011110_10011001_1;
      patterns[64417] = 25'b11111011_10011111_10011010_1;
      patterns[64418] = 25'b11111011_10100000_10011011_1;
      patterns[64419] = 25'b11111011_10100001_10011100_1;
      patterns[64420] = 25'b11111011_10100010_10011101_1;
      patterns[64421] = 25'b11111011_10100011_10011110_1;
      patterns[64422] = 25'b11111011_10100100_10011111_1;
      patterns[64423] = 25'b11111011_10100101_10100000_1;
      patterns[64424] = 25'b11111011_10100110_10100001_1;
      patterns[64425] = 25'b11111011_10100111_10100010_1;
      patterns[64426] = 25'b11111011_10101000_10100011_1;
      patterns[64427] = 25'b11111011_10101001_10100100_1;
      patterns[64428] = 25'b11111011_10101010_10100101_1;
      patterns[64429] = 25'b11111011_10101011_10100110_1;
      patterns[64430] = 25'b11111011_10101100_10100111_1;
      patterns[64431] = 25'b11111011_10101101_10101000_1;
      patterns[64432] = 25'b11111011_10101110_10101001_1;
      patterns[64433] = 25'b11111011_10101111_10101010_1;
      patterns[64434] = 25'b11111011_10110000_10101011_1;
      patterns[64435] = 25'b11111011_10110001_10101100_1;
      patterns[64436] = 25'b11111011_10110010_10101101_1;
      patterns[64437] = 25'b11111011_10110011_10101110_1;
      patterns[64438] = 25'b11111011_10110100_10101111_1;
      patterns[64439] = 25'b11111011_10110101_10110000_1;
      patterns[64440] = 25'b11111011_10110110_10110001_1;
      patterns[64441] = 25'b11111011_10110111_10110010_1;
      patterns[64442] = 25'b11111011_10111000_10110011_1;
      patterns[64443] = 25'b11111011_10111001_10110100_1;
      patterns[64444] = 25'b11111011_10111010_10110101_1;
      patterns[64445] = 25'b11111011_10111011_10110110_1;
      patterns[64446] = 25'b11111011_10111100_10110111_1;
      patterns[64447] = 25'b11111011_10111101_10111000_1;
      patterns[64448] = 25'b11111011_10111110_10111001_1;
      patterns[64449] = 25'b11111011_10111111_10111010_1;
      patterns[64450] = 25'b11111011_11000000_10111011_1;
      patterns[64451] = 25'b11111011_11000001_10111100_1;
      patterns[64452] = 25'b11111011_11000010_10111101_1;
      patterns[64453] = 25'b11111011_11000011_10111110_1;
      patterns[64454] = 25'b11111011_11000100_10111111_1;
      patterns[64455] = 25'b11111011_11000101_11000000_1;
      patterns[64456] = 25'b11111011_11000110_11000001_1;
      patterns[64457] = 25'b11111011_11000111_11000010_1;
      patterns[64458] = 25'b11111011_11001000_11000011_1;
      patterns[64459] = 25'b11111011_11001001_11000100_1;
      patterns[64460] = 25'b11111011_11001010_11000101_1;
      patterns[64461] = 25'b11111011_11001011_11000110_1;
      patterns[64462] = 25'b11111011_11001100_11000111_1;
      patterns[64463] = 25'b11111011_11001101_11001000_1;
      patterns[64464] = 25'b11111011_11001110_11001001_1;
      patterns[64465] = 25'b11111011_11001111_11001010_1;
      patterns[64466] = 25'b11111011_11010000_11001011_1;
      patterns[64467] = 25'b11111011_11010001_11001100_1;
      patterns[64468] = 25'b11111011_11010010_11001101_1;
      patterns[64469] = 25'b11111011_11010011_11001110_1;
      patterns[64470] = 25'b11111011_11010100_11001111_1;
      patterns[64471] = 25'b11111011_11010101_11010000_1;
      patterns[64472] = 25'b11111011_11010110_11010001_1;
      patterns[64473] = 25'b11111011_11010111_11010010_1;
      patterns[64474] = 25'b11111011_11011000_11010011_1;
      patterns[64475] = 25'b11111011_11011001_11010100_1;
      patterns[64476] = 25'b11111011_11011010_11010101_1;
      patterns[64477] = 25'b11111011_11011011_11010110_1;
      patterns[64478] = 25'b11111011_11011100_11010111_1;
      patterns[64479] = 25'b11111011_11011101_11011000_1;
      patterns[64480] = 25'b11111011_11011110_11011001_1;
      patterns[64481] = 25'b11111011_11011111_11011010_1;
      patterns[64482] = 25'b11111011_11100000_11011011_1;
      patterns[64483] = 25'b11111011_11100001_11011100_1;
      patterns[64484] = 25'b11111011_11100010_11011101_1;
      patterns[64485] = 25'b11111011_11100011_11011110_1;
      patterns[64486] = 25'b11111011_11100100_11011111_1;
      patterns[64487] = 25'b11111011_11100101_11100000_1;
      patterns[64488] = 25'b11111011_11100110_11100001_1;
      patterns[64489] = 25'b11111011_11100111_11100010_1;
      patterns[64490] = 25'b11111011_11101000_11100011_1;
      patterns[64491] = 25'b11111011_11101001_11100100_1;
      patterns[64492] = 25'b11111011_11101010_11100101_1;
      patterns[64493] = 25'b11111011_11101011_11100110_1;
      patterns[64494] = 25'b11111011_11101100_11100111_1;
      patterns[64495] = 25'b11111011_11101101_11101000_1;
      patterns[64496] = 25'b11111011_11101110_11101001_1;
      patterns[64497] = 25'b11111011_11101111_11101010_1;
      patterns[64498] = 25'b11111011_11110000_11101011_1;
      patterns[64499] = 25'b11111011_11110001_11101100_1;
      patterns[64500] = 25'b11111011_11110010_11101101_1;
      patterns[64501] = 25'b11111011_11110011_11101110_1;
      patterns[64502] = 25'b11111011_11110100_11101111_1;
      patterns[64503] = 25'b11111011_11110101_11110000_1;
      patterns[64504] = 25'b11111011_11110110_11110001_1;
      patterns[64505] = 25'b11111011_11110111_11110010_1;
      patterns[64506] = 25'b11111011_11111000_11110011_1;
      patterns[64507] = 25'b11111011_11111001_11110100_1;
      patterns[64508] = 25'b11111011_11111010_11110101_1;
      patterns[64509] = 25'b11111011_11111011_11110110_1;
      patterns[64510] = 25'b11111011_11111100_11110111_1;
      patterns[64511] = 25'b11111011_11111101_11111000_1;
      patterns[64512] = 25'b11111011_11111110_11111001_1;
      patterns[64513] = 25'b11111011_11111111_11111010_1;
      patterns[64514] = 25'b11111100_00000000_11111100_0;
      patterns[64515] = 25'b11111100_00000001_11111101_0;
      patterns[64516] = 25'b11111100_00000010_11111110_0;
      patterns[64517] = 25'b11111100_00000011_11111111_0;
      patterns[64518] = 25'b11111100_00000100_00000000_1;
      patterns[64519] = 25'b11111100_00000101_00000001_1;
      patterns[64520] = 25'b11111100_00000110_00000010_1;
      patterns[64521] = 25'b11111100_00000111_00000011_1;
      patterns[64522] = 25'b11111100_00001000_00000100_1;
      patterns[64523] = 25'b11111100_00001001_00000101_1;
      patterns[64524] = 25'b11111100_00001010_00000110_1;
      patterns[64525] = 25'b11111100_00001011_00000111_1;
      patterns[64526] = 25'b11111100_00001100_00001000_1;
      patterns[64527] = 25'b11111100_00001101_00001001_1;
      patterns[64528] = 25'b11111100_00001110_00001010_1;
      patterns[64529] = 25'b11111100_00001111_00001011_1;
      patterns[64530] = 25'b11111100_00010000_00001100_1;
      patterns[64531] = 25'b11111100_00010001_00001101_1;
      patterns[64532] = 25'b11111100_00010010_00001110_1;
      patterns[64533] = 25'b11111100_00010011_00001111_1;
      patterns[64534] = 25'b11111100_00010100_00010000_1;
      patterns[64535] = 25'b11111100_00010101_00010001_1;
      patterns[64536] = 25'b11111100_00010110_00010010_1;
      patterns[64537] = 25'b11111100_00010111_00010011_1;
      patterns[64538] = 25'b11111100_00011000_00010100_1;
      patterns[64539] = 25'b11111100_00011001_00010101_1;
      patterns[64540] = 25'b11111100_00011010_00010110_1;
      patterns[64541] = 25'b11111100_00011011_00010111_1;
      patterns[64542] = 25'b11111100_00011100_00011000_1;
      patterns[64543] = 25'b11111100_00011101_00011001_1;
      patterns[64544] = 25'b11111100_00011110_00011010_1;
      patterns[64545] = 25'b11111100_00011111_00011011_1;
      patterns[64546] = 25'b11111100_00100000_00011100_1;
      patterns[64547] = 25'b11111100_00100001_00011101_1;
      patterns[64548] = 25'b11111100_00100010_00011110_1;
      patterns[64549] = 25'b11111100_00100011_00011111_1;
      patterns[64550] = 25'b11111100_00100100_00100000_1;
      patterns[64551] = 25'b11111100_00100101_00100001_1;
      patterns[64552] = 25'b11111100_00100110_00100010_1;
      patterns[64553] = 25'b11111100_00100111_00100011_1;
      patterns[64554] = 25'b11111100_00101000_00100100_1;
      patterns[64555] = 25'b11111100_00101001_00100101_1;
      patterns[64556] = 25'b11111100_00101010_00100110_1;
      patterns[64557] = 25'b11111100_00101011_00100111_1;
      patterns[64558] = 25'b11111100_00101100_00101000_1;
      patterns[64559] = 25'b11111100_00101101_00101001_1;
      patterns[64560] = 25'b11111100_00101110_00101010_1;
      patterns[64561] = 25'b11111100_00101111_00101011_1;
      patterns[64562] = 25'b11111100_00110000_00101100_1;
      patterns[64563] = 25'b11111100_00110001_00101101_1;
      patterns[64564] = 25'b11111100_00110010_00101110_1;
      patterns[64565] = 25'b11111100_00110011_00101111_1;
      patterns[64566] = 25'b11111100_00110100_00110000_1;
      patterns[64567] = 25'b11111100_00110101_00110001_1;
      patterns[64568] = 25'b11111100_00110110_00110010_1;
      patterns[64569] = 25'b11111100_00110111_00110011_1;
      patterns[64570] = 25'b11111100_00111000_00110100_1;
      patterns[64571] = 25'b11111100_00111001_00110101_1;
      patterns[64572] = 25'b11111100_00111010_00110110_1;
      patterns[64573] = 25'b11111100_00111011_00110111_1;
      patterns[64574] = 25'b11111100_00111100_00111000_1;
      patterns[64575] = 25'b11111100_00111101_00111001_1;
      patterns[64576] = 25'b11111100_00111110_00111010_1;
      patterns[64577] = 25'b11111100_00111111_00111011_1;
      patterns[64578] = 25'b11111100_01000000_00111100_1;
      patterns[64579] = 25'b11111100_01000001_00111101_1;
      patterns[64580] = 25'b11111100_01000010_00111110_1;
      patterns[64581] = 25'b11111100_01000011_00111111_1;
      patterns[64582] = 25'b11111100_01000100_01000000_1;
      patterns[64583] = 25'b11111100_01000101_01000001_1;
      patterns[64584] = 25'b11111100_01000110_01000010_1;
      patterns[64585] = 25'b11111100_01000111_01000011_1;
      patterns[64586] = 25'b11111100_01001000_01000100_1;
      patterns[64587] = 25'b11111100_01001001_01000101_1;
      patterns[64588] = 25'b11111100_01001010_01000110_1;
      patterns[64589] = 25'b11111100_01001011_01000111_1;
      patterns[64590] = 25'b11111100_01001100_01001000_1;
      patterns[64591] = 25'b11111100_01001101_01001001_1;
      patterns[64592] = 25'b11111100_01001110_01001010_1;
      patterns[64593] = 25'b11111100_01001111_01001011_1;
      patterns[64594] = 25'b11111100_01010000_01001100_1;
      patterns[64595] = 25'b11111100_01010001_01001101_1;
      patterns[64596] = 25'b11111100_01010010_01001110_1;
      patterns[64597] = 25'b11111100_01010011_01001111_1;
      patterns[64598] = 25'b11111100_01010100_01010000_1;
      patterns[64599] = 25'b11111100_01010101_01010001_1;
      patterns[64600] = 25'b11111100_01010110_01010010_1;
      patterns[64601] = 25'b11111100_01010111_01010011_1;
      patterns[64602] = 25'b11111100_01011000_01010100_1;
      patterns[64603] = 25'b11111100_01011001_01010101_1;
      patterns[64604] = 25'b11111100_01011010_01010110_1;
      patterns[64605] = 25'b11111100_01011011_01010111_1;
      patterns[64606] = 25'b11111100_01011100_01011000_1;
      patterns[64607] = 25'b11111100_01011101_01011001_1;
      patterns[64608] = 25'b11111100_01011110_01011010_1;
      patterns[64609] = 25'b11111100_01011111_01011011_1;
      patterns[64610] = 25'b11111100_01100000_01011100_1;
      patterns[64611] = 25'b11111100_01100001_01011101_1;
      patterns[64612] = 25'b11111100_01100010_01011110_1;
      patterns[64613] = 25'b11111100_01100011_01011111_1;
      patterns[64614] = 25'b11111100_01100100_01100000_1;
      patterns[64615] = 25'b11111100_01100101_01100001_1;
      patterns[64616] = 25'b11111100_01100110_01100010_1;
      patterns[64617] = 25'b11111100_01100111_01100011_1;
      patterns[64618] = 25'b11111100_01101000_01100100_1;
      patterns[64619] = 25'b11111100_01101001_01100101_1;
      patterns[64620] = 25'b11111100_01101010_01100110_1;
      patterns[64621] = 25'b11111100_01101011_01100111_1;
      patterns[64622] = 25'b11111100_01101100_01101000_1;
      patterns[64623] = 25'b11111100_01101101_01101001_1;
      patterns[64624] = 25'b11111100_01101110_01101010_1;
      patterns[64625] = 25'b11111100_01101111_01101011_1;
      patterns[64626] = 25'b11111100_01110000_01101100_1;
      patterns[64627] = 25'b11111100_01110001_01101101_1;
      patterns[64628] = 25'b11111100_01110010_01101110_1;
      patterns[64629] = 25'b11111100_01110011_01101111_1;
      patterns[64630] = 25'b11111100_01110100_01110000_1;
      patterns[64631] = 25'b11111100_01110101_01110001_1;
      patterns[64632] = 25'b11111100_01110110_01110010_1;
      patterns[64633] = 25'b11111100_01110111_01110011_1;
      patterns[64634] = 25'b11111100_01111000_01110100_1;
      patterns[64635] = 25'b11111100_01111001_01110101_1;
      patterns[64636] = 25'b11111100_01111010_01110110_1;
      patterns[64637] = 25'b11111100_01111011_01110111_1;
      patterns[64638] = 25'b11111100_01111100_01111000_1;
      patterns[64639] = 25'b11111100_01111101_01111001_1;
      patterns[64640] = 25'b11111100_01111110_01111010_1;
      patterns[64641] = 25'b11111100_01111111_01111011_1;
      patterns[64642] = 25'b11111100_10000000_01111100_1;
      patterns[64643] = 25'b11111100_10000001_01111101_1;
      patterns[64644] = 25'b11111100_10000010_01111110_1;
      patterns[64645] = 25'b11111100_10000011_01111111_1;
      patterns[64646] = 25'b11111100_10000100_10000000_1;
      patterns[64647] = 25'b11111100_10000101_10000001_1;
      patterns[64648] = 25'b11111100_10000110_10000010_1;
      patterns[64649] = 25'b11111100_10000111_10000011_1;
      patterns[64650] = 25'b11111100_10001000_10000100_1;
      patterns[64651] = 25'b11111100_10001001_10000101_1;
      patterns[64652] = 25'b11111100_10001010_10000110_1;
      patterns[64653] = 25'b11111100_10001011_10000111_1;
      patterns[64654] = 25'b11111100_10001100_10001000_1;
      patterns[64655] = 25'b11111100_10001101_10001001_1;
      patterns[64656] = 25'b11111100_10001110_10001010_1;
      patterns[64657] = 25'b11111100_10001111_10001011_1;
      patterns[64658] = 25'b11111100_10010000_10001100_1;
      patterns[64659] = 25'b11111100_10010001_10001101_1;
      patterns[64660] = 25'b11111100_10010010_10001110_1;
      patterns[64661] = 25'b11111100_10010011_10001111_1;
      patterns[64662] = 25'b11111100_10010100_10010000_1;
      patterns[64663] = 25'b11111100_10010101_10010001_1;
      patterns[64664] = 25'b11111100_10010110_10010010_1;
      patterns[64665] = 25'b11111100_10010111_10010011_1;
      patterns[64666] = 25'b11111100_10011000_10010100_1;
      patterns[64667] = 25'b11111100_10011001_10010101_1;
      patterns[64668] = 25'b11111100_10011010_10010110_1;
      patterns[64669] = 25'b11111100_10011011_10010111_1;
      patterns[64670] = 25'b11111100_10011100_10011000_1;
      patterns[64671] = 25'b11111100_10011101_10011001_1;
      patterns[64672] = 25'b11111100_10011110_10011010_1;
      patterns[64673] = 25'b11111100_10011111_10011011_1;
      patterns[64674] = 25'b11111100_10100000_10011100_1;
      patterns[64675] = 25'b11111100_10100001_10011101_1;
      patterns[64676] = 25'b11111100_10100010_10011110_1;
      patterns[64677] = 25'b11111100_10100011_10011111_1;
      patterns[64678] = 25'b11111100_10100100_10100000_1;
      patterns[64679] = 25'b11111100_10100101_10100001_1;
      patterns[64680] = 25'b11111100_10100110_10100010_1;
      patterns[64681] = 25'b11111100_10100111_10100011_1;
      patterns[64682] = 25'b11111100_10101000_10100100_1;
      patterns[64683] = 25'b11111100_10101001_10100101_1;
      patterns[64684] = 25'b11111100_10101010_10100110_1;
      patterns[64685] = 25'b11111100_10101011_10100111_1;
      patterns[64686] = 25'b11111100_10101100_10101000_1;
      patterns[64687] = 25'b11111100_10101101_10101001_1;
      patterns[64688] = 25'b11111100_10101110_10101010_1;
      patterns[64689] = 25'b11111100_10101111_10101011_1;
      patterns[64690] = 25'b11111100_10110000_10101100_1;
      patterns[64691] = 25'b11111100_10110001_10101101_1;
      patterns[64692] = 25'b11111100_10110010_10101110_1;
      patterns[64693] = 25'b11111100_10110011_10101111_1;
      patterns[64694] = 25'b11111100_10110100_10110000_1;
      patterns[64695] = 25'b11111100_10110101_10110001_1;
      patterns[64696] = 25'b11111100_10110110_10110010_1;
      patterns[64697] = 25'b11111100_10110111_10110011_1;
      patterns[64698] = 25'b11111100_10111000_10110100_1;
      patterns[64699] = 25'b11111100_10111001_10110101_1;
      patterns[64700] = 25'b11111100_10111010_10110110_1;
      patterns[64701] = 25'b11111100_10111011_10110111_1;
      patterns[64702] = 25'b11111100_10111100_10111000_1;
      patterns[64703] = 25'b11111100_10111101_10111001_1;
      patterns[64704] = 25'b11111100_10111110_10111010_1;
      patterns[64705] = 25'b11111100_10111111_10111011_1;
      patterns[64706] = 25'b11111100_11000000_10111100_1;
      patterns[64707] = 25'b11111100_11000001_10111101_1;
      patterns[64708] = 25'b11111100_11000010_10111110_1;
      patterns[64709] = 25'b11111100_11000011_10111111_1;
      patterns[64710] = 25'b11111100_11000100_11000000_1;
      patterns[64711] = 25'b11111100_11000101_11000001_1;
      patterns[64712] = 25'b11111100_11000110_11000010_1;
      patterns[64713] = 25'b11111100_11000111_11000011_1;
      patterns[64714] = 25'b11111100_11001000_11000100_1;
      patterns[64715] = 25'b11111100_11001001_11000101_1;
      patterns[64716] = 25'b11111100_11001010_11000110_1;
      patterns[64717] = 25'b11111100_11001011_11000111_1;
      patterns[64718] = 25'b11111100_11001100_11001000_1;
      patterns[64719] = 25'b11111100_11001101_11001001_1;
      patterns[64720] = 25'b11111100_11001110_11001010_1;
      patterns[64721] = 25'b11111100_11001111_11001011_1;
      patterns[64722] = 25'b11111100_11010000_11001100_1;
      patterns[64723] = 25'b11111100_11010001_11001101_1;
      patterns[64724] = 25'b11111100_11010010_11001110_1;
      patterns[64725] = 25'b11111100_11010011_11001111_1;
      patterns[64726] = 25'b11111100_11010100_11010000_1;
      patterns[64727] = 25'b11111100_11010101_11010001_1;
      patterns[64728] = 25'b11111100_11010110_11010010_1;
      patterns[64729] = 25'b11111100_11010111_11010011_1;
      patterns[64730] = 25'b11111100_11011000_11010100_1;
      patterns[64731] = 25'b11111100_11011001_11010101_1;
      patterns[64732] = 25'b11111100_11011010_11010110_1;
      patterns[64733] = 25'b11111100_11011011_11010111_1;
      patterns[64734] = 25'b11111100_11011100_11011000_1;
      patterns[64735] = 25'b11111100_11011101_11011001_1;
      patterns[64736] = 25'b11111100_11011110_11011010_1;
      patterns[64737] = 25'b11111100_11011111_11011011_1;
      patterns[64738] = 25'b11111100_11100000_11011100_1;
      patterns[64739] = 25'b11111100_11100001_11011101_1;
      patterns[64740] = 25'b11111100_11100010_11011110_1;
      patterns[64741] = 25'b11111100_11100011_11011111_1;
      patterns[64742] = 25'b11111100_11100100_11100000_1;
      patterns[64743] = 25'b11111100_11100101_11100001_1;
      patterns[64744] = 25'b11111100_11100110_11100010_1;
      patterns[64745] = 25'b11111100_11100111_11100011_1;
      patterns[64746] = 25'b11111100_11101000_11100100_1;
      patterns[64747] = 25'b11111100_11101001_11100101_1;
      patterns[64748] = 25'b11111100_11101010_11100110_1;
      patterns[64749] = 25'b11111100_11101011_11100111_1;
      patterns[64750] = 25'b11111100_11101100_11101000_1;
      patterns[64751] = 25'b11111100_11101101_11101001_1;
      patterns[64752] = 25'b11111100_11101110_11101010_1;
      patterns[64753] = 25'b11111100_11101111_11101011_1;
      patterns[64754] = 25'b11111100_11110000_11101100_1;
      patterns[64755] = 25'b11111100_11110001_11101101_1;
      patterns[64756] = 25'b11111100_11110010_11101110_1;
      patterns[64757] = 25'b11111100_11110011_11101111_1;
      patterns[64758] = 25'b11111100_11110100_11110000_1;
      patterns[64759] = 25'b11111100_11110101_11110001_1;
      patterns[64760] = 25'b11111100_11110110_11110010_1;
      patterns[64761] = 25'b11111100_11110111_11110011_1;
      patterns[64762] = 25'b11111100_11111000_11110100_1;
      patterns[64763] = 25'b11111100_11111001_11110101_1;
      patterns[64764] = 25'b11111100_11111010_11110110_1;
      patterns[64765] = 25'b11111100_11111011_11110111_1;
      patterns[64766] = 25'b11111100_11111100_11111000_1;
      patterns[64767] = 25'b11111100_11111101_11111001_1;
      patterns[64768] = 25'b11111100_11111110_11111010_1;
      patterns[64769] = 25'b11111100_11111111_11111011_1;
      patterns[64770] = 25'b11111101_00000000_11111101_0;
      patterns[64771] = 25'b11111101_00000001_11111110_0;
      patterns[64772] = 25'b11111101_00000010_11111111_0;
      patterns[64773] = 25'b11111101_00000011_00000000_1;
      patterns[64774] = 25'b11111101_00000100_00000001_1;
      patterns[64775] = 25'b11111101_00000101_00000010_1;
      patterns[64776] = 25'b11111101_00000110_00000011_1;
      patterns[64777] = 25'b11111101_00000111_00000100_1;
      patterns[64778] = 25'b11111101_00001000_00000101_1;
      patterns[64779] = 25'b11111101_00001001_00000110_1;
      patterns[64780] = 25'b11111101_00001010_00000111_1;
      patterns[64781] = 25'b11111101_00001011_00001000_1;
      patterns[64782] = 25'b11111101_00001100_00001001_1;
      patterns[64783] = 25'b11111101_00001101_00001010_1;
      patterns[64784] = 25'b11111101_00001110_00001011_1;
      patterns[64785] = 25'b11111101_00001111_00001100_1;
      patterns[64786] = 25'b11111101_00010000_00001101_1;
      patterns[64787] = 25'b11111101_00010001_00001110_1;
      patterns[64788] = 25'b11111101_00010010_00001111_1;
      patterns[64789] = 25'b11111101_00010011_00010000_1;
      patterns[64790] = 25'b11111101_00010100_00010001_1;
      patterns[64791] = 25'b11111101_00010101_00010010_1;
      patterns[64792] = 25'b11111101_00010110_00010011_1;
      patterns[64793] = 25'b11111101_00010111_00010100_1;
      patterns[64794] = 25'b11111101_00011000_00010101_1;
      patterns[64795] = 25'b11111101_00011001_00010110_1;
      patterns[64796] = 25'b11111101_00011010_00010111_1;
      patterns[64797] = 25'b11111101_00011011_00011000_1;
      patterns[64798] = 25'b11111101_00011100_00011001_1;
      patterns[64799] = 25'b11111101_00011101_00011010_1;
      patterns[64800] = 25'b11111101_00011110_00011011_1;
      patterns[64801] = 25'b11111101_00011111_00011100_1;
      patterns[64802] = 25'b11111101_00100000_00011101_1;
      patterns[64803] = 25'b11111101_00100001_00011110_1;
      patterns[64804] = 25'b11111101_00100010_00011111_1;
      patterns[64805] = 25'b11111101_00100011_00100000_1;
      patterns[64806] = 25'b11111101_00100100_00100001_1;
      patterns[64807] = 25'b11111101_00100101_00100010_1;
      patterns[64808] = 25'b11111101_00100110_00100011_1;
      patterns[64809] = 25'b11111101_00100111_00100100_1;
      patterns[64810] = 25'b11111101_00101000_00100101_1;
      patterns[64811] = 25'b11111101_00101001_00100110_1;
      patterns[64812] = 25'b11111101_00101010_00100111_1;
      patterns[64813] = 25'b11111101_00101011_00101000_1;
      patterns[64814] = 25'b11111101_00101100_00101001_1;
      patterns[64815] = 25'b11111101_00101101_00101010_1;
      patterns[64816] = 25'b11111101_00101110_00101011_1;
      patterns[64817] = 25'b11111101_00101111_00101100_1;
      patterns[64818] = 25'b11111101_00110000_00101101_1;
      patterns[64819] = 25'b11111101_00110001_00101110_1;
      patterns[64820] = 25'b11111101_00110010_00101111_1;
      patterns[64821] = 25'b11111101_00110011_00110000_1;
      patterns[64822] = 25'b11111101_00110100_00110001_1;
      patterns[64823] = 25'b11111101_00110101_00110010_1;
      patterns[64824] = 25'b11111101_00110110_00110011_1;
      patterns[64825] = 25'b11111101_00110111_00110100_1;
      patterns[64826] = 25'b11111101_00111000_00110101_1;
      patterns[64827] = 25'b11111101_00111001_00110110_1;
      patterns[64828] = 25'b11111101_00111010_00110111_1;
      patterns[64829] = 25'b11111101_00111011_00111000_1;
      patterns[64830] = 25'b11111101_00111100_00111001_1;
      patterns[64831] = 25'b11111101_00111101_00111010_1;
      patterns[64832] = 25'b11111101_00111110_00111011_1;
      patterns[64833] = 25'b11111101_00111111_00111100_1;
      patterns[64834] = 25'b11111101_01000000_00111101_1;
      patterns[64835] = 25'b11111101_01000001_00111110_1;
      patterns[64836] = 25'b11111101_01000010_00111111_1;
      patterns[64837] = 25'b11111101_01000011_01000000_1;
      patterns[64838] = 25'b11111101_01000100_01000001_1;
      patterns[64839] = 25'b11111101_01000101_01000010_1;
      patterns[64840] = 25'b11111101_01000110_01000011_1;
      patterns[64841] = 25'b11111101_01000111_01000100_1;
      patterns[64842] = 25'b11111101_01001000_01000101_1;
      patterns[64843] = 25'b11111101_01001001_01000110_1;
      patterns[64844] = 25'b11111101_01001010_01000111_1;
      patterns[64845] = 25'b11111101_01001011_01001000_1;
      patterns[64846] = 25'b11111101_01001100_01001001_1;
      patterns[64847] = 25'b11111101_01001101_01001010_1;
      patterns[64848] = 25'b11111101_01001110_01001011_1;
      patterns[64849] = 25'b11111101_01001111_01001100_1;
      patterns[64850] = 25'b11111101_01010000_01001101_1;
      patterns[64851] = 25'b11111101_01010001_01001110_1;
      patterns[64852] = 25'b11111101_01010010_01001111_1;
      patterns[64853] = 25'b11111101_01010011_01010000_1;
      patterns[64854] = 25'b11111101_01010100_01010001_1;
      patterns[64855] = 25'b11111101_01010101_01010010_1;
      patterns[64856] = 25'b11111101_01010110_01010011_1;
      patterns[64857] = 25'b11111101_01010111_01010100_1;
      patterns[64858] = 25'b11111101_01011000_01010101_1;
      patterns[64859] = 25'b11111101_01011001_01010110_1;
      patterns[64860] = 25'b11111101_01011010_01010111_1;
      patterns[64861] = 25'b11111101_01011011_01011000_1;
      patterns[64862] = 25'b11111101_01011100_01011001_1;
      patterns[64863] = 25'b11111101_01011101_01011010_1;
      patterns[64864] = 25'b11111101_01011110_01011011_1;
      patterns[64865] = 25'b11111101_01011111_01011100_1;
      patterns[64866] = 25'b11111101_01100000_01011101_1;
      patterns[64867] = 25'b11111101_01100001_01011110_1;
      patterns[64868] = 25'b11111101_01100010_01011111_1;
      patterns[64869] = 25'b11111101_01100011_01100000_1;
      patterns[64870] = 25'b11111101_01100100_01100001_1;
      patterns[64871] = 25'b11111101_01100101_01100010_1;
      patterns[64872] = 25'b11111101_01100110_01100011_1;
      patterns[64873] = 25'b11111101_01100111_01100100_1;
      patterns[64874] = 25'b11111101_01101000_01100101_1;
      patterns[64875] = 25'b11111101_01101001_01100110_1;
      patterns[64876] = 25'b11111101_01101010_01100111_1;
      patterns[64877] = 25'b11111101_01101011_01101000_1;
      patterns[64878] = 25'b11111101_01101100_01101001_1;
      patterns[64879] = 25'b11111101_01101101_01101010_1;
      patterns[64880] = 25'b11111101_01101110_01101011_1;
      patterns[64881] = 25'b11111101_01101111_01101100_1;
      patterns[64882] = 25'b11111101_01110000_01101101_1;
      patterns[64883] = 25'b11111101_01110001_01101110_1;
      patterns[64884] = 25'b11111101_01110010_01101111_1;
      patterns[64885] = 25'b11111101_01110011_01110000_1;
      patterns[64886] = 25'b11111101_01110100_01110001_1;
      patterns[64887] = 25'b11111101_01110101_01110010_1;
      patterns[64888] = 25'b11111101_01110110_01110011_1;
      patterns[64889] = 25'b11111101_01110111_01110100_1;
      patterns[64890] = 25'b11111101_01111000_01110101_1;
      patterns[64891] = 25'b11111101_01111001_01110110_1;
      patterns[64892] = 25'b11111101_01111010_01110111_1;
      patterns[64893] = 25'b11111101_01111011_01111000_1;
      patterns[64894] = 25'b11111101_01111100_01111001_1;
      patterns[64895] = 25'b11111101_01111101_01111010_1;
      patterns[64896] = 25'b11111101_01111110_01111011_1;
      patterns[64897] = 25'b11111101_01111111_01111100_1;
      patterns[64898] = 25'b11111101_10000000_01111101_1;
      patterns[64899] = 25'b11111101_10000001_01111110_1;
      patterns[64900] = 25'b11111101_10000010_01111111_1;
      patterns[64901] = 25'b11111101_10000011_10000000_1;
      patterns[64902] = 25'b11111101_10000100_10000001_1;
      patterns[64903] = 25'b11111101_10000101_10000010_1;
      patterns[64904] = 25'b11111101_10000110_10000011_1;
      patterns[64905] = 25'b11111101_10000111_10000100_1;
      patterns[64906] = 25'b11111101_10001000_10000101_1;
      patterns[64907] = 25'b11111101_10001001_10000110_1;
      patterns[64908] = 25'b11111101_10001010_10000111_1;
      patterns[64909] = 25'b11111101_10001011_10001000_1;
      patterns[64910] = 25'b11111101_10001100_10001001_1;
      patterns[64911] = 25'b11111101_10001101_10001010_1;
      patterns[64912] = 25'b11111101_10001110_10001011_1;
      patterns[64913] = 25'b11111101_10001111_10001100_1;
      patterns[64914] = 25'b11111101_10010000_10001101_1;
      patterns[64915] = 25'b11111101_10010001_10001110_1;
      patterns[64916] = 25'b11111101_10010010_10001111_1;
      patterns[64917] = 25'b11111101_10010011_10010000_1;
      patterns[64918] = 25'b11111101_10010100_10010001_1;
      patterns[64919] = 25'b11111101_10010101_10010010_1;
      patterns[64920] = 25'b11111101_10010110_10010011_1;
      patterns[64921] = 25'b11111101_10010111_10010100_1;
      patterns[64922] = 25'b11111101_10011000_10010101_1;
      patterns[64923] = 25'b11111101_10011001_10010110_1;
      patterns[64924] = 25'b11111101_10011010_10010111_1;
      patterns[64925] = 25'b11111101_10011011_10011000_1;
      patterns[64926] = 25'b11111101_10011100_10011001_1;
      patterns[64927] = 25'b11111101_10011101_10011010_1;
      patterns[64928] = 25'b11111101_10011110_10011011_1;
      patterns[64929] = 25'b11111101_10011111_10011100_1;
      patterns[64930] = 25'b11111101_10100000_10011101_1;
      patterns[64931] = 25'b11111101_10100001_10011110_1;
      patterns[64932] = 25'b11111101_10100010_10011111_1;
      patterns[64933] = 25'b11111101_10100011_10100000_1;
      patterns[64934] = 25'b11111101_10100100_10100001_1;
      patterns[64935] = 25'b11111101_10100101_10100010_1;
      patterns[64936] = 25'b11111101_10100110_10100011_1;
      patterns[64937] = 25'b11111101_10100111_10100100_1;
      patterns[64938] = 25'b11111101_10101000_10100101_1;
      patterns[64939] = 25'b11111101_10101001_10100110_1;
      patterns[64940] = 25'b11111101_10101010_10100111_1;
      patterns[64941] = 25'b11111101_10101011_10101000_1;
      patterns[64942] = 25'b11111101_10101100_10101001_1;
      patterns[64943] = 25'b11111101_10101101_10101010_1;
      patterns[64944] = 25'b11111101_10101110_10101011_1;
      patterns[64945] = 25'b11111101_10101111_10101100_1;
      patterns[64946] = 25'b11111101_10110000_10101101_1;
      patterns[64947] = 25'b11111101_10110001_10101110_1;
      patterns[64948] = 25'b11111101_10110010_10101111_1;
      patterns[64949] = 25'b11111101_10110011_10110000_1;
      patterns[64950] = 25'b11111101_10110100_10110001_1;
      patterns[64951] = 25'b11111101_10110101_10110010_1;
      patterns[64952] = 25'b11111101_10110110_10110011_1;
      patterns[64953] = 25'b11111101_10110111_10110100_1;
      patterns[64954] = 25'b11111101_10111000_10110101_1;
      patterns[64955] = 25'b11111101_10111001_10110110_1;
      patterns[64956] = 25'b11111101_10111010_10110111_1;
      patterns[64957] = 25'b11111101_10111011_10111000_1;
      patterns[64958] = 25'b11111101_10111100_10111001_1;
      patterns[64959] = 25'b11111101_10111101_10111010_1;
      patterns[64960] = 25'b11111101_10111110_10111011_1;
      patterns[64961] = 25'b11111101_10111111_10111100_1;
      patterns[64962] = 25'b11111101_11000000_10111101_1;
      patterns[64963] = 25'b11111101_11000001_10111110_1;
      patterns[64964] = 25'b11111101_11000010_10111111_1;
      patterns[64965] = 25'b11111101_11000011_11000000_1;
      patterns[64966] = 25'b11111101_11000100_11000001_1;
      patterns[64967] = 25'b11111101_11000101_11000010_1;
      patterns[64968] = 25'b11111101_11000110_11000011_1;
      patterns[64969] = 25'b11111101_11000111_11000100_1;
      patterns[64970] = 25'b11111101_11001000_11000101_1;
      patterns[64971] = 25'b11111101_11001001_11000110_1;
      patterns[64972] = 25'b11111101_11001010_11000111_1;
      patterns[64973] = 25'b11111101_11001011_11001000_1;
      patterns[64974] = 25'b11111101_11001100_11001001_1;
      patterns[64975] = 25'b11111101_11001101_11001010_1;
      patterns[64976] = 25'b11111101_11001110_11001011_1;
      patterns[64977] = 25'b11111101_11001111_11001100_1;
      patterns[64978] = 25'b11111101_11010000_11001101_1;
      patterns[64979] = 25'b11111101_11010001_11001110_1;
      patterns[64980] = 25'b11111101_11010010_11001111_1;
      patterns[64981] = 25'b11111101_11010011_11010000_1;
      patterns[64982] = 25'b11111101_11010100_11010001_1;
      patterns[64983] = 25'b11111101_11010101_11010010_1;
      patterns[64984] = 25'b11111101_11010110_11010011_1;
      patterns[64985] = 25'b11111101_11010111_11010100_1;
      patterns[64986] = 25'b11111101_11011000_11010101_1;
      patterns[64987] = 25'b11111101_11011001_11010110_1;
      patterns[64988] = 25'b11111101_11011010_11010111_1;
      patterns[64989] = 25'b11111101_11011011_11011000_1;
      patterns[64990] = 25'b11111101_11011100_11011001_1;
      patterns[64991] = 25'b11111101_11011101_11011010_1;
      patterns[64992] = 25'b11111101_11011110_11011011_1;
      patterns[64993] = 25'b11111101_11011111_11011100_1;
      patterns[64994] = 25'b11111101_11100000_11011101_1;
      patterns[64995] = 25'b11111101_11100001_11011110_1;
      patterns[64996] = 25'b11111101_11100010_11011111_1;
      patterns[64997] = 25'b11111101_11100011_11100000_1;
      patterns[64998] = 25'b11111101_11100100_11100001_1;
      patterns[64999] = 25'b11111101_11100101_11100010_1;
      patterns[65000] = 25'b11111101_11100110_11100011_1;
      patterns[65001] = 25'b11111101_11100111_11100100_1;
      patterns[65002] = 25'b11111101_11101000_11100101_1;
      patterns[65003] = 25'b11111101_11101001_11100110_1;
      patterns[65004] = 25'b11111101_11101010_11100111_1;
      patterns[65005] = 25'b11111101_11101011_11101000_1;
      patterns[65006] = 25'b11111101_11101100_11101001_1;
      patterns[65007] = 25'b11111101_11101101_11101010_1;
      patterns[65008] = 25'b11111101_11101110_11101011_1;
      patterns[65009] = 25'b11111101_11101111_11101100_1;
      patterns[65010] = 25'b11111101_11110000_11101101_1;
      patterns[65011] = 25'b11111101_11110001_11101110_1;
      patterns[65012] = 25'b11111101_11110010_11101111_1;
      patterns[65013] = 25'b11111101_11110011_11110000_1;
      patterns[65014] = 25'b11111101_11110100_11110001_1;
      patterns[65015] = 25'b11111101_11110101_11110010_1;
      patterns[65016] = 25'b11111101_11110110_11110011_1;
      patterns[65017] = 25'b11111101_11110111_11110100_1;
      patterns[65018] = 25'b11111101_11111000_11110101_1;
      patterns[65019] = 25'b11111101_11111001_11110110_1;
      patterns[65020] = 25'b11111101_11111010_11110111_1;
      patterns[65021] = 25'b11111101_11111011_11111000_1;
      patterns[65022] = 25'b11111101_11111100_11111001_1;
      patterns[65023] = 25'b11111101_11111101_11111010_1;
      patterns[65024] = 25'b11111101_11111110_11111011_1;
      patterns[65025] = 25'b11111101_11111111_11111100_1;
      patterns[65026] = 25'b11111110_00000000_11111110_0;
      patterns[65027] = 25'b11111110_00000001_11111111_0;
      patterns[65028] = 25'b11111110_00000010_00000000_1;
      patterns[65029] = 25'b11111110_00000011_00000001_1;
      patterns[65030] = 25'b11111110_00000100_00000010_1;
      patterns[65031] = 25'b11111110_00000101_00000011_1;
      patterns[65032] = 25'b11111110_00000110_00000100_1;
      patterns[65033] = 25'b11111110_00000111_00000101_1;
      patterns[65034] = 25'b11111110_00001000_00000110_1;
      patterns[65035] = 25'b11111110_00001001_00000111_1;
      patterns[65036] = 25'b11111110_00001010_00001000_1;
      patterns[65037] = 25'b11111110_00001011_00001001_1;
      patterns[65038] = 25'b11111110_00001100_00001010_1;
      patterns[65039] = 25'b11111110_00001101_00001011_1;
      patterns[65040] = 25'b11111110_00001110_00001100_1;
      patterns[65041] = 25'b11111110_00001111_00001101_1;
      patterns[65042] = 25'b11111110_00010000_00001110_1;
      patterns[65043] = 25'b11111110_00010001_00001111_1;
      patterns[65044] = 25'b11111110_00010010_00010000_1;
      patterns[65045] = 25'b11111110_00010011_00010001_1;
      patterns[65046] = 25'b11111110_00010100_00010010_1;
      patterns[65047] = 25'b11111110_00010101_00010011_1;
      patterns[65048] = 25'b11111110_00010110_00010100_1;
      patterns[65049] = 25'b11111110_00010111_00010101_1;
      patterns[65050] = 25'b11111110_00011000_00010110_1;
      patterns[65051] = 25'b11111110_00011001_00010111_1;
      patterns[65052] = 25'b11111110_00011010_00011000_1;
      patterns[65053] = 25'b11111110_00011011_00011001_1;
      patterns[65054] = 25'b11111110_00011100_00011010_1;
      patterns[65055] = 25'b11111110_00011101_00011011_1;
      patterns[65056] = 25'b11111110_00011110_00011100_1;
      patterns[65057] = 25'b11111110_00011111_00011101_1;
      patterns[65058] = 25'b11111110_00100000_00011110_1;
      patterns[65059] = 25'b11111110_00100001_00011111_1;
      patterns[65060] = 25'b11111110_00100010_00100000_1;
      patterns[65061] = 25'b11111110_00100011_00100001_1;
      patterns[65062] = 25'b11111110_00100100_00100010_1;
      patterns[65063] = 25'b11111110_00100101_00100011_1;
      patterns[65064] = 25'b11111110_00100110_00100100_1;
      patterns[65065] = 25'b11111110_00100111_00100101_1;
      patterns[65066] = 25'b11111110_00101000_00100110_1;
      patterns[65067] = 25'b11111110_00101001_00100111_1;
      patterns[65068] = 25'b11111110_00101010_00101000_1;
      patterns[65069] = 25'b11111110_00101011_00101001_1;
      patterns[65070] = 25'b11111110_00101100_00101010_1;
      patterns[65071] = 25'b11111110_00101101_00101011_1;
      patterns[65072] = 25'b11111110_00101110_00101100_1;
      patterns[65073] = 25'b11111110_00101111_00101101_1;
      patterns[65074] = 25'b11111110_00110000_00101110_1;
      patterns[65075] = 25'b11111110_00110001_00101111_1;
      patterns[65076] = 25'b11111110_00110010_00110000_1;
      patterns[65077] = 25'b11111110_00110011_00110001_1;
      patterns[65078] = 25'b11111110_00110100_00110010_1;
      patterns[65079] = 25'b11111110_00110101_00110011_1;
      patterns[65080] = 25'b11111110_00110110_00110100_1;
      patterns[65081] = 25'b11111110_00110111_00110101_1;
      patterns[65082] = 25'b11111110_00111000_00110110_1;
      patterns[65083] = 25'b11111110_00111001_00110111_1;
      patterns[65084] = 25'b11111110_00111010_00111000_1;
      patterns[65085] = 25'b11111110_00111011_00111001_1;
      patterns[65086] = 25'b11111110_00111100_00111010_1;
      patterns[65087] = 25'b11111110_00111101_00111011_1;
      patterns[65088] = 25'b11111110_00111110_00111100_1;
      patterns[65089] = 25'b11111110_00111111_00111101_1;
      patterns[65090] = 25'b11111110_01000000_00111110_1;
      patterns[65091] = 25'b11111110_01000001_00111111_1;
      patterns[65092] = 25'b11111110_01000010_01000000_1;
      patterns[65093] = 25'b11111110_01000011_01000001_1;
      patterns[65094] = 25'b11111110_01000100_01000010_1;
      patterns[65095] = 25'b11111110_01000101_01000011_1;
      patterns[65096] = 25'b11111110_01000110_01000100_1;
      patterns[65097] = 25'b11111110_01000111_01000101_1;
      patterns[65098] = 25'b11111110_01001000_01000110_1;
      patterns[65099] = 25'b11111110_01001001_01000111_1;
      patterns[65100] = 25'b11111110_01001010_01001000_1;
      patterns[65101] = 25'b11111110_01001011_01001001_1;
      patterns[65102] = 25'b11111110_01001100_01001010_1;
      patterns[65103] = 25'b11111110_01001101_01001011_1;
      patterns[65104] = 25'b11111110_01001110_01001100_1;
      patterns[65105] = 25'b11111110_01001111_01001101_1;
      patterns[65106] = 25'b11111110_01010000_01001110_1;
      patterns[65107] = 25'b11111110_01010001_01001111_1;
      patterns[65108] = 25'b11111110_01010010_01010000_1;
      patterns[65109] = 25'b11111110_01010011_01010001_1;
      patterns[65110] = 25'b11111110_01010100_01010010_1;
      patterns[65111] = 25'b11111110_01010101_01010011_1;
      patterns[65112] = 25'b11111110_01010110_01010100_1;
      patterns[65113] = 25'b11111110_01010111_01010101_1;
      patterns[65114] = 25'b11111110_01011000_01010110_1;
      patterns[65115] = 25'b11111110_01011001_01010111_1;
      patterns[65116] = 25'b11111110_01011010_01011000_1;
      patterns[65117] = 25'b11111110_01011011_01011001_1;
      patterns[65118] = 25'b11111110_01011100_01011010_1;
      patterns[65119] = 25'b11111110_01011101_01011011_1;
      patterns[65120] = 25'b11111110_01011110_01011100_1;
      patterns[65121] = 25'b11111110_01011111_01011101_1;
      patterns[65122] = 25'b11111110_01100000_01011110_1;
      patterns[65123] = 25'b11111110_01100001_01011111_1;
      patterns[65124] = 25'b11111110_01100010_01100000_1;
      patterns[65125] = 25'b11111110_01100011_01100001_1;
      patterns[65126] = 25'b11111110_01100100_01100010_1;
      patterns[65127] = 25'b11111110_01100101_01100011_1;
      patterns[65128] = 25'b11111110_01100110_01100100_1;
      patterns[65129] = 25'b11111110_01100111_01100101_1;
      patterns[65130] = 25'b11111110_01101000_01100110_1;
      patterns[65131] = 25'b11111110_01101001_01100111_1;
      patterns[65132] = 25'b11111110_01101010_01101000_1;
      patterns[65133] = 25'b11111110_01101011_01101001_1;
      patterns[65134] = 25'b11111110_01101100_01101010_1;
      patterns[65135] = 25'b11111110_01101101_01101011_1;
      patterns[65136] = 25'b11111110_01101110_01101100_1;
      patterns[65137] = 25'b11111110_01101111_01101101_1;
      patterns[65138] = 25'b11111110_01110000_01101110_1;
      patterns[65139] = 25'b11111110_01110001_01101111_1;
      patterns[65140] = 25'b11111110_01110010_01110000_1;
      patterns[65141] = 25'b11111110_01110011_01110001_1;
      patterns[65142] = 25'b11111110_01110100_01110010_1;
      patterns[65143] = 25'b11111110_01110101_01110011_1;
      patterns[65144] = 25'b11111110_01110110_01110100_1;
      patterns[65145] = 25'b11111110_01110111_01110101_1;
      patterns[65146] = 25'b11111110_01111000_01110110_1;
      patterns[65147] = 25'b11111110_01111001_01110111_1;
      patterns[65148] = 25'b11111110_01111010_01111000_1;
      patterns[65149] = 25'b11111110_01111011_01111001_1;
      patterns[65150] = 25'b11111110_01111100_01111010_1;
      patterns[65151] = 25'b11111110_01111101_01111011_1;
      patterns[65152] = 25'b11111110_01111110_01111100_1;
      patterns[65153] = 25'b11111110_01111111_01111101_1;
      patterns[65154] = 25'b11111110_10000000_01111110_1;
      patterns[65155] = 25'b11111110_10000001_01111111_1;
      patterns[65156] = 25'b11111110_10000010_10000000_1;
      patterns[65157] = 25'b11111110_10000011_10000001_1;
      patterns[65158] = 25'b11111110_10000100_10000010_1;
      patterns[65159] = 25'b11111110_10000101_10000011_1;
      patterns[65160] = 25'b11111110_10000110_10000100_1;
      patterns[65161] = 25'b11111110_10000111_10000101_1;
      patterns[65162] = 25'b11111110_10001000_10000110_1;
      patterns[65163] = 25'b11111110_10001001_10000111_1;
      patterns[65164] = 25'b11111110_10001010_10001000_1;
      patterns[65165] = 25'b11111110_10001011_10001001_1;
      patterns[65166] = 25'b11111110_10001100_10001010_1;
      patterns[65167] = 25'b11111110_10001101_10001011_1;
      patterns[65168] = 25'b11111110_10001110_10001100_1;
      patterns[65169] = 25'b11111110_10001111_10001101_1;
      patterns[65170] = 25'b11111110_10010000_10001110_1;
      patterns[65171] = 25'b11111110_10010001_10001111_1;
      patterns[65172] = 25'b11111110_10010010_10010000_1;
      patterns[65173] = 25'b11111110_10010011_10010001_1;
      patterns[65174] = 25'b11111110_10010100_10010010_1;
      patterns[65175] = 25'b11111110_10010101_10010011_1;
      patterns[65176] = 25'b11111110_10010110_10010100_1;
      patterns[65177] = 25'b11111110_10010111_10010101_1;
      patterns[65178] = 25'b11111110_10011000_10010110_1;
      patterns[65179] = 25'b11111110_10011001_10010111_1;
      patterns[65180] = 25'b11111110_10011010_10011000_1;
      patterns[65181] = 25'b11111110_10011011_10011001_1;
      patterns[65182] = 25'b11111110_10011100_10011010_1;
      patterns[65183] = 25'b11111110_10011101_10011011_1;
      patterns[65184] = 25'b11111110_10011110_10011100_1;
      patterns[65185] = 25'b11111110_10011111_10011101_1;
      patterns[65186] = 25'b11111110_10100000_10011110_1;
      patterns[65187] = 25'b11111110_10100001_10011111_1;
      patterns[65188] = 25'b11111110_10100010_10100000_1;
      patterns[65189] = 25'b11111110_10100011_10100001_1;
      patterns[65190] = 25'b11111110_10100100_10100010_1;
      patterns[65191] = 25'b11111110_10100101_10100011_1;
      patterns[65192] = 25'b11111110_10100110_10100100_1;
      patterns[65193] = 25'b11111110_10100111_10100101_1;
      patterns[65194] = 25'b11111110_10101000_10100110_1;
      patterns[65195] = 25'b11111110_10101001_10100111_1;
      patterns[65196] = 25'b11111110_10101010_10101000_1;
      patterns[65197] = 25'b11111110_10101011_10101001_1;
      patterns[65198] = 25'b11111110_10101100_10101010_1;
      patterns[65199] = 25'b11111110_10101101_10101011_1;
      patterns[65200] = 25'b11111110_10101110_10101100_1;
      patterns[65201] = 25'b11111110_10101111_10101101_1;
      patterns[65202] = 25'b11111110_10110000_10101110_1;
      patterns[65203] = 25'b11111110_10110001_10101111_1;
      patterns[65204] = 25'b11111110_10110010_10110000_1;
      patterns[65205] = 25'b11111110_10110011_10110001_1;
      patterns[65206] = 25'b11111110_10110100_10110010_1;
      patterns[65207] = 25'b11111110_10110101_10110011_1;
      patterns[65208] = 25'b11111110_10110110_10110100_1;
      patterns[65209] = 25'b11111110_10110111_10110101_1;
      patterns[65210] = 25'b11111110_10111000_10110110_1;
      patterns[65211] = 25'b11111110_10111001_10110111_1;
      patterns[65212] = 25'b11111110_10111010_10111000_1;
      patterns[65213] = 25'b11111110_10111011_10111001_1;
      patterns[65214] = 25'b11111110_10111100_10111010_1;
      patterns[65215] = 25'b11111110_10111101_10111011_1;
      patterns[65216] = 25'b11111110_10111110_10111100_1;
      patterns[65217] = 25'b11111110_10111111_10111101_1;
      patterns[65218] = 25'b11111110_11000000_10111110_1;
      patterns[65219] = 25'b11111110_11000001_10111111_1;
      patterns[65220] = 25'b11111110_11000010_11000000_1;
      patterns[65221] = 25'b11111110_11000011_11000001_1;
      patterns[65222] = 25'b11111110_11000100_11000010_1;
      patterns[65223] = 25'b11111110_11000101_11000011_1;
      patterns[65224] = 25'b11111110_11000110_11000100_1;
      patterns[65225] = 25'b11111110_11000111_11000101_1;
      patterns[65226] = 25'b11111110_11001000_11000110_1;
      patterns[65227] = 25'b11111110_11001001_11000111_1;
      patterns[65228] = 25'b11111110_11001010_11001000_1;
      patterns[65229] = 25'b11111110_11001011_11001001_1;
      patterns[65230] = 25'b11111110_11001100_11001010_1;
      patterns[65231] = 25'b11111110_11001101_11001011_1;
      patterns[65232] = 25'b11111110_11001110_11001100_1;
      patterns[65233] = 25'b11111110_11001111_11001101_1;
      patterns[65234] = 25'b11111110_11010000_11001110_1;
      patterns[65235] = 25'b11111110_11010001_11001111_1;
      patterns[65236] = 25'b11111110_11010010_11010000_1;
      patterns[65237] = 25'b11111110_11010011_11010001_1;
      patterns[65238] = 25'b11111110_11010100_11010010_1;
      patterns[65239] = 25'b11111110_11010101_11010011_1;
      patterns[65240] = 25'b11111110_11010110_11010100_1;
      patterns[65241] = 25'b11111110_11010111_11010101_1;
      patterns[65242] = 25'b11111110_11011000_11010110_1;
      patterns[65243] = 25'b11111110_11011001_11010111_1;
      patterns[65244] = 25'b11111110_11011010_11011000_1;
      patterns[65245] = 25'b11111110_11011011_11011001_1;
      patterns[65246] = 25'b11111110_11011100_11011010_1;
      patterns[65247] = 25'b11111110_11011101_11011011_1;
      patterns[65248] = 25'b11111110_11011110_11011100_1;
      patterns[65249] = 25'b11111110_11011111_11011101_1;
      patterns[65250] = 25'b11111110_11100000_11011110_1;
      patterns[65251] = 25'b11111110_11100001_11011111_1;
      patterns[65252] = 25'b11111110_11100010_11100000_1;
      patterns[65253] = 25'b11111110_11100011_11100001_1;
      patterns[65254] = 25'b11111110_11100100_11100010_1;
      patterns[65255] = 25'b11111110_11100101_11100011_1;
      patterns[65256] = 25'b11111110_11100110_11100100_1;
      patterns[65257] = 25'b11111110_11100111_11100101_1;
      patterns[65258] = 25'b11111110_11101000_11100110_1;
      patterns[65259] = 25'b11111110_11101001_11100111_1;
      patterns[65260] = 25'b11111110_11101010_11101000_1;
      patterns[65261] = 25'b11111110_11101011_11101001_1;
      patterns[65262] = 25'b11111110_11101100_11101010_1;
      patterns[65263] = 25'b11111110_11101101_11101011_1;
      patterns[65264] = 25'b11111110_11101110_11101100_1;
      patterns[65265] = 25'b11111110_11101111_11101101_1;
      patterns[65266] = 25'b11111110_11110000_11101110_1;
      patterns[65267] = 25'b11111110_11110001_11101111_1;
      patterns[65268] = 25'b11111110_11110010_11110000_1;
      patterns[65269] = 25'b11111110_11110011_11110001_1;
      patterns[65270] = 25'b11111110_11110100_11110010_1;
      patterns[65271] = 25'b11111110_11110101_11110011_1;
      patterns[65272] = 25'b11111110_11110110_11110100_1;
      patterns[65273] = 25'b11111110_11110111_11110101_1;
      patterns[65274] = 25'b11111110_11111000_11110110_1;
      patterns[65275] = 25'b11111110_11111001_11110111_1;
      patterns[65276] = 25'b11111110_11111010_11111000_1;
      patterns[65277] = 25'b11111110_11111011_11111001_1;
      patterns[65278] = 25'b11111110_11111100_11111010_1;
      patterns[65279] = 25'b11111110_11111101_11111011_1;
      patterns[65280] = 25'b11111110_11111110_11111100_1;
      patterns[65281] = 25'b11111110_11111111_11111101_1;
      patterns[65282] = 25'b11111111_00000000_11111111_0;
      patterns[65283] = 25'b11111111_00000001_00000000_1;
      patterns[65284] = 25'b11111111_00000010_00000001_1;
      patterns[65285] = 25'b11111111_00000011_00000010_1;
      patterns[65286] = 25'b11111111_00000100_00000011_1;
      patterns[65287] = 25'b11111111_00000101_00000100_1;
      patterns[65288] = 25'b11111111_00000110_00000101_1;
      patterns[65289] = 25'b11111111_00000111_00000110_1;
      patterns[65290] = 25'b11111111_00001000_00000111_1;
      patterns[65291] = 25'b11111111_00001001_00001000_1;
      patterns[65292] = 25'b11111111_00001010_00001001_1;
      patterns[65293] = 25'b11111111_00001011_00001010_1;
      patterns[65294] = 25'b11111111_00001100_00001011_1;
      patterns[65295] = 25'b11111111_00001101_00001100_1;
      patterns[65296] = 25'b11111111_00001110_00001101_1;
      patterns[65297] = 25'b11111111_00001111_00001110_1;
      patterns[65298] = 25'b11111111_00010000_00001111_1;
      patterns[65299] = 25'b11111111_00010001_00010000_1;
      patterns[65300] = 25'b11111111_00010010_00010001_1;
      patterns[65301] = 25'b11111111_00010011_00010010_1;
      patterns[65302] = 25'b11111111_00010100_00010011_1;
      patterns[65303] = 25'b11111111_00010101_00010100_1;
      patterns[65304] = 25'b11111111_00010110_00010101_1;
      patterns[65305] = 25'b11111111_00010111_00010110_1;
      patterns[65306] = 25'b11111111_00011000_00010111_1;
      patterns[65307] = 25'b11111111_00011001_00011000_1;
      patterns[65308] = 25'b11111111_00011010_00011001_1;
      patterns[65309] = 25'b11111111_00011011_00011010_1;
      patterns[65310] = 25'b11111111_00011100_00011011_1;
      patterns[65311] = 25'b11111111_00011101_00011100_1;
      patterns[65312] = 25'b11111111_00011110_00011101_1;
      patterns[65313] = 25'b11111111_00011111_00011110_1;
      patterns[65314] = 25'b11111111_00100000_00011111_1;
      patterns[65315] = 25'b11111111_00100001_00100000_1;
      patterns[65316] = 25'b11111111_00100010_00100001_1;
      patterns[65317] = 25'b11111111_00100011_00100010_1;
      patterns[65318] = 25'b11111111_00100100_00100011_1;
      patterns[65319] = 25'b11111111_00100101_00100100_1;
      patterns[65320] = 25'b11111111_00100110_00100101_1;
      patterns[65321] = 25'b11111111_00100111_00100110_1;
      patterns[65322] = 25'b11111111_00101000_00100111_1;
      patterns[65323] = 25'b11111111_00101001_00101000_1;
      patterns[65324] = 25'b11111111_00101010_00101001_1;
      patterns[65325] = 25'b11111111_00101011_00101010_1;
      patterns[65326] = 25'b11111111_00101100_00101011_1;
      patterns[65327] = 25'b11111111_00101101_00101100_1;
      patterns[65328] = 25'b11111111_00101110_00101101_1;
      patterns[65329] = 25'b11111111_00101111_00101110_1;
      patterns[65330] = 25'b11111111_00110000_00101111_1;
      patterns[65331] = 25'b11111111_00110001_00110000_1;
      patterns[65332] = 25'b11111111_00110010_00110001_1;
      patterns[65333] = 25'b11111111_00110011_00110010_1;
      patterns[65334] = 25'b11111111_00110100_00110011_1;
      patterns[65335] = 25'b11111111_00110101_00110100_1;
      patterns[65336] = 25'b11111111_00110110_00110101_1;
      patterns[65337] = 25'b11111111_00110111_00110110_1;
      patterns[65338] = 25'b11111111_00111000_00110111_1;
      patterns[65339] = 25'b11111111_00111001_00111000_1;
      patterns[65340] = 25'b11111111_00111010_00111001_1;
      patterns[65341] = 25'b11111111_00111011_00111010_1;
      patterns[65342] = 25'b11111111_00111100_00111011_1;
      patterns[65343] = 25'b11111111_00111101_00111100_1;
      patterns[65344] = 25'b11111111_00111110_00111101_1;
      patterns[65345] = 25'b11111111_00111111_00111110_1;
      patterns[65346] = 25'b11111111_01000000_00111111_1;
      patterns[65347] = 25'b11111111_01000001_01000000_1;
      patterns[65348] = 25'b11111111_01000010_01000001_1;
      patterns[65349] = 25'b11111111_01000011_01000010_1;
      patterns[65350] = 25'b11111111_01000100_01000011_1;
      patterns[65351] = 25'b11111111_01000101_01000100_1;
      patterns[65352] = 25'b11111111_01000110_01000101_1;
      patterns[65353] = 25'b11111111_01000111_01000110_1;
      patterns[65354] = 25'b11111111_01001000_01000111_1;
      patterns[65355] = 25'b11111111_01001001_01001000_1;
      patterns[65356] = 25'b11111111_01001010_01001001_1;
      patterns[65357] = 25'b11111111_01001011_01001010_1;
      patterns[65358] = 25'b11111111_01001100_01001011_1;
      patterns[65359] = 25'b11111111_01001101_01001100_1;
      patterns[65360] = 25'b11111111_01001110_01001101_1;
      patterns[65361] = 25'b11111111_01001111_01001110_1;
      patterns[65362] = 25'b11111111_01010000_01001111_1;
      patterns[65363] = 25'b11111111_01010001_01010000_1;
      patterns[65364] = 25'b11111111_01010010_01010001_1;
      patterns[65365] = 25'b11111111_01010011_01010010_1;
      patterns[65366] = 25'b11111111_01010100_01010011_1;
      patterns[65367] = 25'b11111111_01010101_01010100_1;
      patterns[65368] = 25'b11111111_01010110_01010101_1;
      patterns[65369] = 25'b11111111_01010111_01010110_1;
      patterns[65370] = 25'b11111111_01011000_01010111_1;
      patterns[65371] = 25'b11111111_01011001_01011000_1;
      patterns[65372] = 25'b11111111_01011010_01011001_1;
      patterns[65373] = 25'b11111111_01011011_01011010_1;
      patterns[65374] = 25'b11111111_01011100_01011011_1;
      patterns[65375] = 25'b11111111_01011101_01011100_1;
      patterns[65376] = 25'b11111111_01011110_01011101_1;
      patterns[65377] = 25'b11111111_01011111_01011110_1;
      patterns[65378] = 25'b11111111_01100000_01011111_1;
      patterns[65379] = 25'b11111111_01100001_01100000_1;
      patterns[65380] = 25'b11111111_01100010_01100001_1;
      patterns[65381] = 25'b11111111_01100011_01100010_1;
      patterns[65382] = 25'b11111111_01100100_01100011_1;
      patterns[65383] = 25'b11111111_01100101_01100100_1;
      patterns[65384] = 25'b11111111_01100110_01100101_1;
      patterns[65385] = 25'b11111111_01100111_01100110_1;
      patterns[65386] = 25'b11111111_01101000_01100111_1;
      patterns[65387] = 25'b11111111_01101001_01101000_1;
      patterns[65388] = 25'b11111111_01101010_01101001_1;
      patterns[65389] = 25'b11111111_01101011_01101010_1;
      patterns[65390] = 25'b11111111_01101100_01101011_1;
      patterns[65391] = 25'b11111111_01101101_01101100_1;
      patterns[65392] = 25'b11111111_01101110_01101101_1;
      patterns[65393] = 25'b11111111_01101111_01101110_1;
      patterns[65394] = 25'b11111111_01110000_01101111_1;
      patterns[65395] = 25'b11111111_01110001_01110000_1;
      patterns[65396] = 25'b11111111_01110010_01110001_1;
      patterns[65397] = 25'b11111111_01110011_01110010_1;
      patterns[65398] = 25'b11111111_01110100_01110011_1;
      patterns[65399] = 25'b11111111_01110101_01110100_1;
      patterns[65400] = 25'b11111111_01110110_01110101_1;
      patterns[65401] = 25'b11111111_01110111_01110110_1;
      patterns[65402] = 25'b11111111_01111000_01110111_1;
      patterns[65403] = 25'b11111111_01111001_01111000_1;
      patterns[65404] = 25'b11111111_01111010_01111001_1;
      patterns[65405] = 25'b11111111_01111011_01111010_1;
      patterns[65406] = 25'b11111111_01111100_01111011_1;
      patterns[65407] = 25'b11111111_01111101_01111100_1;
      patterns[65408] = 25'b11111111_01111110_01111101_1;
      patterns[65409] = 25'b11111111_01111111_01111110_1;
      patterns[65410] = 25'b11111111_10000000_01111111_1;
      patterns[65411] = 25'b11111111_10000001_10000000_1;
      patterns[65412] = 25'b11111111_10000010_10000001_1;
      patterns[65413] = 25'b11111111_10000011_10000010_1;
      patterns[65414] = 25'b11111111_10000100_10000011_1;
      patterns[65415] = 25'b11111111_10000101_10000100_1;
      patterns[65416] = 25'b11111111_10000110_10000101_1;
      patterns[65417] = 25'b11111111_10000111_10000110_1;
      patterns[65418] = 25'b11111111_10001000_10000111_1;
      patterns[65419] = 25'b11111111_10001001_10001000_1;
      patterns[65420] = 25'b11111111_10001010_10001001_1;
      patterns[65421] = 25'b11111111_10001011_10001010_1;
      patterns[65422] = 25'b11111111_10001100_10001011_1;
      patterns[65423] = 25'b11111111_10001101_10001100_1;
      patterns[65424] = 25'b11111111_10001110_10001101_1;
      patterns[65425] = 25'b11111111_10001111_10001110_1;
      patterns[65426] = 25'b11111111_10010000_10001111_1;
      patterns[65427] = 25'b11111111_10010001_10010000_1;
      patterns[65428] = 25'b11111111_10010010_10010001_1;
      patterns[65429] = 25'b11111111_10010011_10010010_1;
      patterns[65430] = 25'b11111111_10010100_10010011_1;
      patterns[65431] = 25'b11111111_10010101_10010100_1;
      patterns[65432] = 25'b11111111_10010110_10010101_1;
      patterns[65433] = 25'b11111111_10010111_10010110_1;
      patterns[65434] = 25'b11111111_10011000_10010111_1;
      patterns[65435] = 25'b11111111_10011001_10011000_1;
      patterns[65436] = 25'b11111111_10011010_10011001_1;
      patterns[65437] = 25'b11111111_10011011_10011010_1;
      patterns[65438] = 25'b11111111_10011100_10011011_1;
      patterns[65439] = 25'b11111111_10011101_10011100_1;
      patterns[65440] = 25'b11111111_10011110_10011101_1;
      patterns[65441] = 25'b11111111_10011111_10011110_1;
      patterns[65442] = 25'b11111111_10100000_10011111_1;
      patterns[65443] = 25'b11111111_10100001_10100000_1;
      patterns[65444] = 25'b11111111_10100010_10100001_1;
      patterns[65445] = 25'b11111111_10100011_10100010_1;
      patterns[65446] = 25'b11111111_10100100_10100011_1;
      patterns[65447] = 25'b11111111_10100101_10100100_1;
      patterns[65448] = 25'b11111111_10100110_10100101_1;
      patterns[65449] = 25'b11111111_10100111_10100110_1;
      patterns[65450] = 25'b11111111_10101000_10100111_1;
      patterns[65451] = 25'b11111111_10101001_10101000_1;
      patterns[65452] = 25'b11111111_10101010_10101001_1;
      patterns[65453] = 25'b11111111_10101011_10101010_1;
      patterns[65454] = 25'b11111111_10101100_10101011_1;
      patterns[65455] = 25'b11111111_10101101_10101100_1;
      patterns[65456] = 25'b11111111_10101110_10101101_1;
      patterns[65457] = 25'b11111111_10101111_10101110_1;
      patterns[65458] = 25'b11111111_10110000_10101111_1;
      patterns[65459] = 25'b11111111_10110001_10110000_1;
      patterns[65460] = 25'b11111111_10110010_10110001_1;
      patterns[65461] = 25'b11111111_10110011_10110010_1;
      patterns[65462] = 25'b11111111_10110100_10110011_1;
      patterns[65463] = 25'b11111111_10110101_10110100_1;
      patterns[65464] = 25'b11111111_10110110_10110101_1;
      patterns[65465] = 25'b11111111_10110111_10110110_1;
      patterns[65466] = 25'b11111111_10111000_10110111_1;
      patterns[65467] = 25'b11111111_10111001_10111000_1;
      patterns[65468] = 25'b11111111_10111010_10111001_1;
      patterns[65469] = 25'b11111111_10111011_10111010_1;
      patterns[65470] = 25'b11111111_10111100_10111011_1;
      patterns[65471] = 25'b11111111_10111101_10111100_1;
      patterns[65472] = 25'b11111111_10111110_10111101_1;
      patterns[65473] = 25'b11111111_10111111_10111110_1;
      patterns[65474] = 25'b11111111_11000000_10111111_1;
      patterns[65475] = 25'b11111111_11000001_11000000_1;
      patterns[65476] = 25'b11111111_11000010_11000001_1;
      patterns[65477] = 25'b11111111_11000011_11000010_1;
      patterns[65478] = 25'b11111111_11000100_11000011_1;
      patterns[65479] = 25'b11111111_11000101_11000100_1;
      patterns[65480] = 25'b11111111_11000110_11000101_1;
      patterns[65481] = 25'b11111111_11000111_11000110_1;
      patterns[65482] = 25'b11111111_11001000_11000111_1;
      patterns[65483] = 25'b11111111_11001001_11001000_1;
      patterns[65484] = 25'b11111111_11001010_11001001_1;
      patterns[65485] = 25'b11111111_11001011_11001010_1;
      patterns[65486] = 25'b11111111_11001100_11001011_1;
      patterns[65487] = 25'b11111111_11001101_11001100_1;
      patterns[65488] = 25'b11111111_11001110_11001101_1;
      patterns[65489] = 25'b11111111_11001111_11001110_1;
      patterns[65490] = 25'b11111111_11010000_11001111_1;
      patterns[65491] = 25'b11111111_11010001_11010000_1;
      patterns[65492] = 25'b11111111_11010010_11010001_1;
      patterns[65493] = 25'b11111111_11010011_11010010_1;
      patterns[65494] = 25'b11111111_11010100_11010011_1;
      patterns[65495] = 25'b11111111_11010101_11010100_1;
      patterns[65496] = 25'b11111111_11010110_11010101_1;
      patterns[65497] = 25'b11111111_11010111_11010110_1;
      patterns[65498] = 25'b11111111_11011000_11010111_1;
      patterns[65499] = 25'b11111111_11011001_11011000_1;
      patterns[65500] = 25'b11111111_11011010_11011001_1;
      patterns[65501] = 25'b11111111_11011011_11011010_1;
      patterns[65502] = 25'b11111111_11011100_11011011_1;
      patterns[65503] = 25'b11111111_11011101_11011100_1;
      patterns[65504] = 25'b11111111_11011110_11011101_1;
      patterns[65505] = 25'b11111111_11011111_11011110_1;
      patterns[65506] = 25'b11111111_11100000_11011111_1;
      patterns[65507] = 25'b11111111_11100001_11100000_1;
      patterns[65508] = 25'b11111111_11100010_11100001_1;
      patterns[65509] = 25'b11111111_11100011_11100010_1;
      patterns[65510] = 25'b11111111_11100100_11100011_1;
      patterns[65511] = 25'b11111111_11100101_11100100_1;
      patterns[65512] = 25'b11111111_11100110_11100101_1;
      patterns[65513] = 25'b11111111_11100111_11100110_1;
      patterns[65514] = 25'b11111111_11101000_11100111_1;
      patterns[65515] = 25'b11111111_11101001_11101000_1;
      patterns[65516] = 25'b11111111_11101010_11101001_1;
      patterns[65517] = 25'b11111111_11101011_11101010_1;
      patterns[65518] = 25'b11111111_11101100_11101011_1;
      patterns[65519] = 25'b11111111_11101101_11101100_1;
      patterns[65520] = 25'b11111111_11101110_11101101_1;
      patterns[65521] = 25'b11111111_11101111_11101110_1;
      patterns[65522] = 25'b11111111_11110000_11101111_1;
      patterns[65523] = 25'b11111111_11110001_11110000_1;
      patterns[65524] = 25'b11111111_11110010_11110001_1;
      patterns[65525] = 25'b11111111_11110011_11110010_1;
      patterns[65526] = 25'b11111111_11110100_11110011_1;
      patterns[65527] = 25'b11111111_11110101_11110100_1;
      patterns[65528] = 25'b11111111_11110110_11110101_1;
      patterns[65529] = 25'b11111111_11110111_11110110_1;
      patterns[65530] = 25'b11111111_11111000_11110111_1;
      patterns[65531] = 25'b11111111_11111001_11111000_1;
      patterns[65532] = 25'b11111111_11111010_11111001_1;
      patterns[65533] = 25'b11111111_11111011_11111010_1;
      patterns[65534] = 25'b11111111_11111100_11111011_1;
      patterns[65535] = 25'b11111111_11111101_11111100_1;
      patterns[65536] = 25'b11111111_11111110_11111101_1;
      patterns[65537] = 25'b11111111_11111111_11111110_1;

      for (i = 0; i < 65538; i = i + 1)
      begin
        A = patterns[i][24:17];
        B = patterns[i][16:9];
        #10;
        if (patterns[i][8:1] !== 8'hx)
        begin
          if (S !== patterns[i][8:1])
          begin
            $display("%d:S: (assertion error). Expected %h, found %h", i, patterns[i][8:1], S);
            $finish;
          end
        end
        if (patterns[i][0] !== 1'hx)
        begin
          if (C !== patterns[i][0])
          begin
            $display("%d:C: (assertion error). Expected %h, found %h", i, patterns[i][0], C);
            $finish;
          end
        end
      end

      $display("All tests passed.");
    end
    endmodule
